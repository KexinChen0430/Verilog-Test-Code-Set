module ass2(a, b, out);
    input [1:0] a;
    output [3:0] out;
    assign out = a;
endmodule