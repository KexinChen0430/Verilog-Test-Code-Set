module page251;

specify
$timeskew (posedge CP &&& MODE, negedge CPN, 50,, event_based_flag,
remain_active_flag);

endspecify
endmodule