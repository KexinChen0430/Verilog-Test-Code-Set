//commit 389dc7aaae138ed820997ec66714e20a9ecb0a9e
//Author: Zihao Yu <yuzihao@ict.ac.cn>
//Date:   Tue Nov 2 09:03:54 2021 +0800
//
//    test,emu: use jumpfw for flash
//diff --git a/Makefile b/Makefile
//index 7785829..c97164e 100644
//--- a/Makefile
//+++ b/Makefile
//@@ -9,7 +9,8 @@ MEM_GEN = ./scripts/vlsi_mem_gen
// USE_READY_TO_RUN_NEMU = true
// 
// SIMTOP = top.TopMain
//-IMAGE ?= ready-to-run/linux.bin
//+#IMAGE ?= ready-to-run/linux.bin
//+IMAGE ?= /home/yzh/oscpu/NutShell/ready-to-run/busybox-ysyx3.bin
// 
// DATAWIDTH ?= 64
// BOARD ?= sim  # sim  pynq  axu3cg soctest
//@@ -52,7 +53,7 @@ $(SIM_TOP_V): $(SCALA_FILE) $(TEST_FILE)
// 	mill chiselModule.test.runMain $(SIMTOP) -td $(@D) --output-file $(@F) BOARD=$(BOARD) CORE=$(CORE)
// 	sed -i -e 's/_\(aw\|ar\|w\|r\|b\)_\(\|bits_\)/_\1/g' $@
// 
//-ysyxSoC_DIR = ../ysyxSoC-new
//+ysyxSoC_DIR = ../ysyxSoC
// SOC_DIR = $(ysyxSoC_DIR)/ysyx/peripheral
// RAM_DIR = $(ysyxSoC_DIR)/ysyx/ram
// EMU_SOC_V = $(shell find $(SOC_DIR) -name '*.v') $(shell find $(RAM_DIR) -name '*.v') $(ysyxSoC_DIR)/ysyx/soc/ysyxSoCFull.v
module ysyx_210000_SRAMTemplate(
  input         clock,
  input         reset,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [4:0]  io_rreq_bits_setIdx,
  output [31:0] io_rresp_data_0_tag,
  output [1:0]  io_rresp_data_0__type,
  output [38:0] io_rresp_data_0_target,
  output [2:0]  io_rresp_data_0_brIdx,
  output        io_rresp_data_0_valid,
  input         io_wreq_valid,
  input  [4:0]  io_wreq_bits_setIdx,
  input  [31:0] io_wreq_bits_data_tag,
  input  [1:0]  io_wreq_bits_data__type,
  input  [38:0] io_wreq_bits_data_target,
  input  [2:0]  io_wreq_bits_data_brIdx
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [95:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [4:0] array_RW0_addr; // @[SRAMTemplate.scala 128:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 128:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 128:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 128:26]
  wire [76:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 128:26]
  wire [76:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 128:26]
  reg  REG; // @[SRAMTemplate.scala 132:30]
  reg [4:0] REG_1; // @[Counter.scala 60:40]
  wire  _T = REG_1 == 5'h1f; // @[Counter.scala 72:24]
  wire [4:0] _T_2 = REG_1 + 5'h1; // @[Counter.scala 76:24]
  wire  _GEN_1 = REG & _T; // @[Counter.scala 118:17 Counter.scala 118:24]
  wire  _GEN_2 = _GEN_1 ? 1'h0 : REG; // @[SRAMTemplate.scala 134:24 SRAMTemplate.scala 134:38 SRAMTemplate.scala 132:30]
  wire  wen = io_wreq_valid | REG; // @[SRAMTemplate.scala 140:52]
  wire  _T_3 = ~wen; // @[SRAMTemplate.scala 141:41]
  wire  realRen = io_rreq_valid & ~wen; // @[SRAMTemplate.scala 141:38]
  wire [4:0] setIdx = REG ? REG_1 : io_wreq_bits_setIdx; // @[SRAMTemplate.scala 143:19]
  wire [76:0] _T_4 = {io_wreq_bits_data_tag,io_wreq_bits_data__type,io_wreq_bits_data_target,io_wreq_bits_data_brIdx
    ,1'h1}; // @[SRAMTemplate.scala 144:78]
  reg  REG_2; // @[Hold.scala 28:106]
  reg [76:0] REG_3_0; // @[Reg.scala 27:20]
  wire [76:0] _GEN_14 = REG_2 ? array_RW0_rdata_0 : REG_3_0; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  ysyx_210000_array array ( // @[SRAMTemplate.scala 128:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_rdata_0(array_RW0_rdata_0)
  );
  assign io_rreq_ready = ~REG & _T_3; // @[SRAMTemplate.scala 153:33]
  assign io_rresp_data_0_tag = _GEN_14[76:45]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_0__type = _GEN_14[44:43]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_0_target = _GEN_14[42:4]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_0_brIdx = _GEN_14[3:1]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_0_valid = _GEN_14[0]; // @[SRAMTemplate.scala 150:78]
  assign array_RW0_wdata_0 = REG ? 77'h0 : _T_4; // @[SRAMTemplate.scala 144:22]
  assign array_RW0_wmode = io_wreq_valid | REG; // @[SRAMTemplate.scala 140:52]
  assign array_RW0_clk = clock;
  assign array_RW0_en = realRen | wen;
  assign array_RW0_addr = wen ? setIdx : io_rreq_bits_setIdx;
  always @(posedge clock) begin
    REG <= reset | _GEN_2; // @[SRAMTemplate.scala 132:30 SRAMTemplate.scala 132:30]
    if (reset) begin // @[Counter.scala 60:40]
      REG_1 <= 5'h0; // @[Counter.scala 60:40]
    end else if (REG) begin // @[Counter.scala 118:17]
      REG_1 <= _T_2; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Hold.scala 28:106]
      REG_2 <= 1'h0; // @[Hold.scala 28:106]
    end else begin
      REG_2 <= realRen; // @[Hold.scala 28:106]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_0 <= 77'h0; // @[Reg.scala 27:20]
    end else if (REG_2) begin // @[Reg.scala 28:19]
      REG_3_0 <= array_RW0_rdata_0; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  REG_2 = _RAND_2[0:0];
  _RAND_3 = {3{`RANDOM}};
  REG_3_0 = _RAND_3[76:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_BPU_inorder(
  input         clock,
  input         reset,
  input         io_in_pc_valid,
  input  [38:0] io_in_pc_bits,
  output [38:0] io_out_target,
  output        io_out_valid,
  input         io_flush,
  output [2:0]  io_brIdx,
  output        io_crosslineJump,
  input         MOUFlushICache,
  input         bpuUpdateReq_valid,
  input  [38:0] bpuUpdateReq_pc,
  input         bpuUpdateReq_isMissPredict,
  input  [38:0] bpuUpdateReq_actualTarget,
  input         bpuUpdateReq_actualTaken,
  input  [6:0]  bpuUpdateReq_fuOpType,
  input  [1:0]  bpuUpdateReq_btbType,
  input         bpuUpdateReq_isRVC,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
`endif // RANDOMIZE_REG_INIT
  wire  btb_clock; // @[BPU.scala 302:19]
  wire  btb_reset; // @[BPU.scala 302:19]
  wire  btb_io_rreq_ready; // @[BPU.scala 302:19]
  wire  btb_io_rreq_valid; // @[BPU.scala 302:19]
  wire [4:0] btb_io_rreq_bits_setIdx; // @[BPU.scala 302:19]
  wire [31:0] btb_io_rresp_data_0_tag; // @[BPU.scala 302:19]
  wire [1:0] btb_io_rresp_data_0__type; // @[BPU.scala 302:19]
  wire [38:0] btb_io_rresp_data_0_target; // @[BPU.scala 302:19]
  wire [2:0] btb_io_rresp_data_0_brIdx; // @[BPU.scala 302:19]
  wire  btb_io_rresp_data_0_valid; // @[BPU.scala 302:19]
  wire  btb_io_wreq_valid; // @[BPU.scala 302:19]
  wire [4:0] btb_io_wreq_bits_setIdx; // @[BPU.scala 302:19]
  wire [31:0] btb_io_wreq_bits_data_tag; // @[BPU.scala 302:19]
  wire [1:0] btb_io_wreq_bits_data__type; // @[BPU.scala 302:19]
  wire [38:0] btb_io_wreq_bits_data_target; // @[BPU.scala 302:19]
  wire [2:0] btb_io_wreq_bits_data_brIdx; // @[BPU.scala 302:19]
  reg  flush; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_pc_valid ? 1'h0 : flush; // @[StopWatch.scala 26:19 StopWatch.scala 26:23 StopWatch.scala 24:20]
  wire  _GEN_1 = io_flush | _GEN_0; // @[StopWatch.scala 27:20 StopWatch.scala 27:24]
  reg [38:0] pcLatch; // @[Reg.scala 27:20]
  wire [31:0] btbRead_tag = btb_io_rresp_data_0_tag; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire  btbRead_valid = btb_io_rresp_data_0_valid; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire  _T_19 = btb_io_rreq_ready & btb_io_rreq_valid; // @[Decoupled.scala 40:37]
  reg  REG_1; // @[BPU.scala 320:93]
  wire [2:0] btbRead_brIdx = btb_io_rresp_data_0_brIdx; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire  btbHit = btbRead_valid & btbRead_tag == pcLatch[38:7] & ~flush & REG_1 & ~(pcLatch[1] & btbRead_brIdx[0]); // @[BPU.scala 320:131]
  wire  crosslineJump = btbRead_brIdx[2] & btbHit; // @[BPU.scala 327:40]
  wire [1:0] lo = io_out_valid ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg [1:0] pht_0; // @[BPU.scala 337:20]
  reg [1:0] pht_1; // @[BPU.scala 337:20]
  reg [1:0] pht_2; // @[BPU.scala 337:20]
  reg [1:0] pht_3; // @[BPU.scala 337:20]
  reg [1:0] pht_4; // @[BPU.scala 337:20]
  reg [1:0] pht_5; // @[BPU.scala 337:20]
  reg [1:0] pht_6; // @[BPU.scala 337:20]
  reg [1:0] pht_7; // @[BPU.scala 337:20]
  reg [1:0] pht_8; // @[BPU.scala 337:20]
  reg [1:0] pht_9; // @[BPU.scala 337:20]
  reg [1:0] pht_10; // @[BPU.scala 337:20]
  reg [1:0] pht_11; // @[BPU.scala 337:20]
  reg [1:0] pht_12; // @[BPU.scala 337:20]
  reg [1:0] pht_13; // @[BPU.scala 337:20]
  reg [1:0] pht_14; // @[BPU.scala 337:20]
  reg [1:0] pht_15; // @[BPU.scala 337:20]
  reg [1:0] pht_16; // @[BPU.scala 337:20]
  reg [1:0] pht_17; // @[BPU.scala 337:20]
  reg [1:0] pht_18; // @[BPU.scala 337:20]
  reg [1:0] pht_19; // @[BPU.scala 337:20]
  reg [1:0] pht_20; // @[BPU.scala 337:20]
  reg [1:0] pht_21; // @[BPU.scala 337:20]
  reg [1:0] pht_22; // @[BPU.scala 337:20]
  reg [1:0] pht_23; // @[BPU.scala 337:20]
  reg [1:0] pht_24; // @[BPU.scala 337:20]
  reg [1:0] pht_25; // @[BPU.scala 337:20]
  reg [1:0] pht_26; // @[BPU.scala 337:20]
  reg [1:0] pht_27; // @[BPU.scala 337:20]
  reg [1:0] pht_28; // @[BPU.scala 337:20]
  reg [1:0] pht_29; // @[BPU.scala 337:20]
  reg [1:0] pht_30; // @[BPU.scala 337:20]
  reg [1:0] pht_31; // @[BPU.scala 337:20]
  wire [1:0] _GEN_4 = 5'h1 == io_in_pc_bits[6:2] ? pht_1 : pht_0; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_5 = 5'h2 == io_in_pc_bits[6:2] ? pht_2 : _GEN_4; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_6 = 5'h3 == io_in_pc_bits[6:2] ? pht_3 : _GEN_5; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_7 = 5'h4 == io_in_pc_bits[6:2] ? pht_4 : _GEN_6; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_8 = 5'h5 == io_in_pc_bits[6:2] ? pht_5 : _GEN_7; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_9 = 5'h6 == io_in_pc_bits[6:2] ? pht_6 : _GEN_8; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_10 = 5'h7 == io_in_pc_bits[6:2] ? pht_7 : _GEN_9; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_11 = 5'h8 == io_in_pc_bits[6:2] ? pht_8 : _GEN_10; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_12 = 5'h9 == io_in_pc_bits[6:2] ? pht_9 : _GEN_11; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_13 = 5'ha == io_in_pc_bits[6:2] ? pht_10 : _GEN_12; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_14 = 5'hb == io_in_pc_bits[6:2] ? pht_11 : _GEN_13; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_15 = 5'hc == io_in_pc_bits[6:2] ? pht_12 : _GEN_14; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_16 = 5'hd == io_in_pc_bits[6:2] ? pht_13 : _GEN_15; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_17 = 5'he == io_in_pc_bits[6:2] ? pht_14 : _GEN_16; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_18 = 5'hf == io_in_pc_bits[6:2] ? pht_15 : _GEN_17; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_19 = 5'h10 == io_in_pc_bits[6:2] ? pht_16 : _GEN_18; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_20 = 5'h11 == io_in_pc_bits[6:2] ? pht_17 : _GEN_19; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_21 = 5'h12 == io_in_pc_bits[6:2] ? pht_18 : _GEN_20; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_22 = 5'h13 == io_in_pc_bits[6:2] ? pht_19 : _GEN_21; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_23 = 5'h14 == io_in_pc_bits[6:2] ? pht_20 : _GEN_22; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_24 = 5'h15 == io_in_pc_bits[6:2] ? pht_21 : _GEN_23; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_25 = 5'h16 == io_in_pc_bits[6:2] ? pht_22 : _GEN_24; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_26 = 5'h17 == io_in_pc_bits[6:2] ? pht_23 : _GEN_25; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_27 = 5'h18 == io_in_pc_bits[6:2] ? pht_24 : _GEN_26; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_28 = 5'h19 == io_in_pc_bits[6:2] ? pht_25 : _GEN_27; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_29 = 5'h1a == io_in_pc_bits[6:2] ? pht_26 : _GEN_28; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_30 = 5'h1b == io_in_pc_bits[6:2] ? pht_27 : _GEN_29; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_31 = 5'h1c == io_in_pc_bits[6:2] ? pht_28 : _GEN_30; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_32 = 5'h1d == io_in_pc_bits[6:2] ? pht_29 : _GEN_31; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_33 = 5'h1e == io_in_pc_bits[6:2] ? pht_30 : _GEN_32; // @[BPU.scala 338:62 BPU.scala 338:62]
  wire [1:0] _GEN_34 = 5'h1f == io_in_pc_bits[6:2] ? pht_31 : _GEN_33; // @[BPU.scala 338:62 BPU.scala 338:62]
  reg  phtTaken; // @[Reg.scala 27:20]
  reg [38:0] ras_0; // @[BPU.scala 344:20]
  reg [38:0] ras_1; // @[BPU.scala 344:20]
  reg [38:0] ras_2; // @[BPU.scala 344:20]
  reg [38:0] ras_3; // @[BPU.scala 344:20]
  reg [38:0] ras_4; // @[BPU.scala 344:20]
  reg [38:0] ras_5; // @[BPU.scala 344:20]
  reg [38:0] ras_6; // @[BPU.scala 344:20]
  reg [38:0] ras_7; // @[BPU.scala 344:20]
  reg [38:0] ras_8; // @[BPU.scala 344:20]
  reg [38:0] ras_9; // @[BPU.scala 344:20]
  reg [38:0] ras_10; // @[BPU.scala 344:20]
  reg [38:0] ras_11; // @[BPU.scala 344:20]
  reg [38:0] ras_12; // @[BPU.scala 344:20]
  reg [38:0] ras_13; // @[BPU.scala 344:20]
  reg [38:0] ras_14; // @[BPU.scala 344:20]
  reg [38:0] ras_15; // @[BPU.scala 344:20]
  reg [3:0] value; // @[Counter.scala 60:40]
  reg [38:0] rasTarget; // @[Reg.scala 27:20]
  wire [38:0] _GEN_37 = 4'h1 == value ? ras_1 : ras_0; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [38:0] _GEN_38 = 4'h2 == value ? ras_2 : _GEN_37; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [38:0] _GEN_39 = 4'h3 == value ? ras_3 : _GEN_38; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [38:0] _GEN_40 = 4'h4 == value ? ras_4 : _GEN_39; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [38:0] _GEN_41 = 4'h5 == value ? ras_5 : _GEN_40; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [38:0] _GEN_42 = 4'h6 == value ? ras_6 : _GEN_41; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [38:0] _GEN_43 = 4'h7 == value ? ras_7 : _GEN_42; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [38:0] _GEN_44 = 4'h8 == value ? ras_8 : _GEN_43; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [38:0] _GEN_45 = 4'h9 == value ? ras_9 : _GEN_44; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [38:0] _GEN_46 = 4'ha == value ? ras_10 : _GEN_45; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [38:0] _GEN_47 = 4'hb == value ? ras_11 : _GEN_46; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [38:0] _GEN_48 = 4'hc == value ? ras_12 : _GEN_47; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire [38:0] _GEN_49 = 4'hd == value ? ras_13 : _GEN_48; // @[Reg.scala 28:23 Reg.scala 28:23]
  wire  hi = bpuUpdateReq_pc[1]; // @[BPU.scala 355:145]
  wire  lo_1 = ~hi; // @[BPU.scala 355:150]
  wire  hi_hi = bpuUpdateReq_pc[2:0] == 3'h6 & ~bpuUpdateReq_isRVC; // @[BPU.scala 369:46]
  wire [1:0] hi_1 = {hi_hi,hi}; // @[Cat.scala 30:58]
  reg [1:0] cnt; // @[BPU.scala 391:20]
  wire [1:0] _GEN_54 = 5'h1 == bpuUpdateReq_pc[6:2] ? pht_1 : pht_0; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_55 = 5'h2 == bpuUpdateReq_pc[6:2] ? pht_2 : _GEN_54; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_56 = 5'h3 == bpuUpdateReq_pc[6:2] ? pht_3 : _GEN_55; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_57 = 5'h4 == bpuUpdateReq_pc[6:2] ? pht_4 : _GEN_56; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_58 = 5'h5 == bpuUpdateReq_pc[6:2] ? pht_5 : _GEN_57; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_59 = 5'h6 == bpuUpdateReq_pc[6:2] ? pht_6 : _GEN_58; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_60 = 5'h7 == bpuUpdateReq_pc[6:2] ? pht_7 : _GEN_59; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_61 = 5'h8 == bpuUpdateReq_pc[6:2] ? pht_8 : _GEN_60; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_62 = 5'h9 == bpuUpdateReq_pc[6:2] ? pht_9 : _GEN_61; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_63 = 5'ha == bpuUpdateReq_pc[6:2] ? pht_10 : _GEN_62; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_64 = 5'hb == bpuUpdateReq_pc[6:2] ? pht_11 : _GEN_63; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_65 = 5'hc == bpuUpdateReq_pc[6:2] ? pht_12 : _GEN_64; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_66 = 5'hd == bpuUpdateReq_pc[6:2] ? pht_13 : _GEN_65; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_67 = 5'he == bpuUpdateReq_pc[6:2] ? pht_14 : _GEN_66; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_68 = 5'hf == bpuUpdateReq_pc[6:2] ? pht_15 : _GEN_67; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_69 = 5'h10 == bpuUpdateReq_pc[6:2] ? pht_16 : _GEN_68; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_70 = 5'h11 == bpuUpdateReq_pc[6:2] ? pht_17 : _GEN_69; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_71 = 5'h12 == bpuUpdateReq_pc[6:2] ? pht_18 : _GEN_70; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_72 = 5'h13 == bpuUpdateReq_pc[6:2] ? pht_19 : _GEN_71; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_73 = 5'h14 == bpuUpdateReq_pc[6:2] ? pht_20 : _GEN_72; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_74 = 5'h15 == bpuUpdateReq_pc[6:2] ? pht_21 : _GEN_73; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_75 = 5'h16 == bpuUpdateReq_pc[6:2] ? pht_22 : _GEN_74; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_76 = 5'h17 == bpuUpdateReq_pc[6:2] ? pht_23 : _GEN_75; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_77 = 5'h18 == bpuUpdateReq_pc[6:2] ? pht_24 : _GEN_76; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_78 = 5'h19 == bpuUpdateReq_pc[6:2] ? pht_25 : _GEN_77; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_79 = 5'h1a == bpuUpdateReq_pc[6:2] ? pht_26 : _GEN_78; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_80 = 5'h1b == bpuUpdateReq_pc[6:2] ? pht_27 : _GEN_79; // @[BPU.scala 391:20 BPU.scala 391:20]
  wire [1:0] _GEN_81 = 5'h1c == bpuUpdateReq_pc[6:2] ? pht_28 : _GEN_80; // @[BPU.scala 391:20 BPU.scala 391:20]
  reg  reqLatch_valid; // @[BPU.scala 392:25]
  reg [38:0] reqLatch_pc; // @[BPU.scala 392:25]
  reg  reqLatch_actualTaken; // @[BPU.scala 392:25]
  reg [6:0] reqLatch_fuOpType; // @[BPU.scala 392:25]
  wire  _T_73 = ~reqLatch_fuOpType[3]; // @[ALU.scala 65:30]
  wire [1:0] _T_76 = cnt + 2'h1; // @[BPU.scala 395:33]
  wire [1:0] _T_78 = cnt - 2'h1; // @[BPU.scala 395:44]
  wire [1:0] _T_79 = reqLatch_actualTaken ? _T_76 : _T_78; // @[BPU.scala 395:21]
  wire  _T_85 = reqLatch_actualTaken & cnt != 2'h3 | ~reqLatch_actualTaken & cnt != 2'h0; // @[BPU.scala 396:44]
  wire [3:0] _T_91 = value + 4'h1; // @[BPU.scala 406:20]
  wire [38:0] _T_93 = bpuUpdateReq_pc + 39'h2; // @[BPU.scala 406:52]
  wire [38:0] _T_95 = bpuUpdateReq_pc + 39'h4; // @[BPU.scala 406:66]
  wire [38:0] _T_96 = bpuUpdateReq_isRVC ? _T_93 : _T_95; // @[BPU.scala 406:33]
  wire  _T_98 = value == 4'h0; // @[BPU.scala 411:21]
  wire [3:0] _value_T_4 = value - 4'h1; // @[BPU.scala 414:53]
  wire [3:0] _value_T_5 = _T_98 ? 4'h0 : _value_T_4; // @[BPU.scala 414:22]
  wire [1:0] btbRead__type = btb_io_rresp_data_0__type; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire [38:0] btbRead_target = btb_io_rresp_data_0_target; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire [3:0] _T_102 = {1'h1,crosslineJump,lo}; // @[Cat.scala 30:58]
  wire [3:0] _GEN_232 = {{1'd0}, btbRead_brIdx}; // @[BPU.scala 421:30]
  wire [3:0] _T_103 = _GEN_232 & _T_102; // @[BPU.scala 421:30]
  wire  _T_107 = btbRead__type == 2'h0 ? phtTaken : rasTarget != 39'h0; // @[BPU.scala 422:32]
  ysyx_210000_SRAMTemplate btb ( // @[BPU.scala 302:19]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_rreq_ready(btb_io_rreq_ready),
    .io_rreq_valid(btb_io_rreq_valid),
    .io_rreq_bits_setIdx(btb_io_rreq_bits_setIdx),
    .io_rresp_data_0_tag(btb_io_rresp_data_0_tag),
    .io_rresp_data_0__type(btb_io_rresp_data_0__type),
    .io_rresp_data_0_target(btb_io_rresp_data_0_target),
    .io_rresp_data_0_brIdx(btb_io_rresp_data_0_brIdx),
    .io_rresp_data_0_valid(btb_io_rresp_data_0_valid),
    .io_wreq_valid(btb_io_wreq_valid),
    .io_wreq_bits_setIdx(btb_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(btb_io_wreq_bits_data_tag),
    .io_wreq_bits_data__type(btb_io_wreq_bits_data__type),
    .io_wreq_bits_data_target(btb_io_wreq_bits_data_target),
    .io_wreq_bits_data_brIdx(btb_io_wreq_bits_data_brIdx)
  );
  assign io_out_target = btbRead__type == 2'h3 ? rasTarget : btbRead_target; // @[BPU.scala 418:23]
  assign io_out_valid = btbHit & _T_107; // @[BPU.scala 422:26]
  assign io_brIdx = _T_103[2:0]; // @[BPU.scala 421:13]
  assign io_crosslineJump = btbRead_brIdx[2] & btbHit; // @[BPU.scala 327:40]
  assign btb_clock = clock;
  assign btb_reset = reset | (MOUFlushICache | MOUFlushTLB); // @[BPU.scala 308:29]
  assign btb_io_rreq_valid = io_in_pc_valid; // @[BPU.scala 311:22]
  assign btb_io_rreq_bits_setIdx = io_in_pc_bits[6:2]; // @[BPU.scala 35:65]
  assign btb_io_wreq_valid = bpuUpdateReq_isMissPredict & bpuUpdateReq_valid; // @[BPU.scala 377:43]
  assign btb_io_wreq_bits_setIdx = bpuUpdateReq_pc[6:2]; // @[BPU.scala 35:65]
  assign btb_io_wreq_bits_data_tag = bpuUpdateReq_pc[38:7]; // @[BPU.scala 35:65]
  assign btb_io_wreq_bits_data__type = bpuUpdateReq_btbType; // @[BPU.scala 379:26]
  assign btb_io_wreq_bits_data_target = bpuUpdateReq_actualTarget; // @[BPU.scala 379:26]
  assign btb_io_wreq_bits_data_brIdx = {hi_1,lo_1}; // @[Cat.scala 30:58]
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      flush <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      flush <= _GEN_1;
    end
    if (reset) begin // @[Reg.scala 27:20]
      pcLatch <= 39'h30000000; // @[Reg.scala 27:20]
    end else if (io_in_pc_valid) begin // @[Reg.scala 28:19]
      pcLatch <= io_in_pc_bits; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[BPU.scala 320:93]
      REG_1 <= 1'h0; // @[BPU.scala 320:93]
    end else begin
      REG_1 <= _T_19; // @[BPU.scala 320:93]
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_0 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h0 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_0 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_1 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h1 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_1 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_2 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h2 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_2 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_3 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h3 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_3 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_4 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h4 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_4 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_5 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h5 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_5 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_6 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h6 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_6 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_7 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h7 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_7 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_8 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h8 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_8 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_9 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h9 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_9 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_10 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'ha == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_10 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_11 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'hb == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_11 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_12 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'hc == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_12 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_13 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'hd == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_13 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_14 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'he == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_14 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_15 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'hf == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_15 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_16 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h10 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_16 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_17 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h11 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_17 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_18 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h12 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_18 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_19 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h13 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_19 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_20 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h14 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_20 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_21 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h15 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_21 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_22 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h16 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_22 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_23 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h17 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_23 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_24 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h18 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_24 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_25 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h19 == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_25 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_26 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h1a == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_26 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_27 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h1b == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_27 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_28 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h1c == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_28 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_29 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h1d == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_29 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_30 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h1e == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_30 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[BPU.scala 337:20]
      pht_31 <= 2'h0; // @[BPU.scala 337:20]
    end else if (reqLatch_valid & _T_73) begin // @[BPU.scala 393:66]
      if (_T_85) begin // @[BPU.scala 397:16]
        if (5'h1f == reqLatch_pc[6:2]) begin // @[BPU.scala 398:40]
          pht_31 <= _T_79; // @[BPU.scala 398:40]
        end
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      phtTaken <= 1'h0; // @[Reg.scala 27:20]
    end else if (io_in_pc_valid) begin // @[Reg.scala 28:19]
      phtTaken <= _GEN_34[1]; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_0 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'h0 == _T_91) begin // @[BPU.scala 406:27]
          ras_0 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_1 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'h1 == _T_91) begin // @[BPU.scala 406:27]
          ras_1 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_2 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'h2 == _T_91) begin // @[BPU.scala 406:27]
          ras_2 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_3 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'h3 == _T_91) begin // @[BPU.scala 406:27]
          ras_3 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_4 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'h4 == _T_91) begin // @[BPU.scala 406:27]
          ras_4 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_5 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'h5 == _T_91) begin // @[BPU.scala 406:27]
          ras_5 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_6 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'h6 == _T_91) begin // @[BPU.scala 406:27]
          ras_6 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_7 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'h7 == _T_91) begin // @[BPU.scala 406:27]
          ras_7 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_8 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'h8 == _T_91) begin // @[BPU.scala 406:27]
          ras_8 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_9 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'h9 == _T_91) begin // @[BPU.scala 406:27]
          ras_9 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_10 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'ha == _T_91) begin // @[BPU.scala 406:27]
          ras_10 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_11 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'hb == _T_91) begin // @[BPU.scala 406:27]
          ras_11 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_12 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'hc == _T_91) begin // @[BPU.scala 406:27]
          ras_12 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_13 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'hd == _T_91) begin // @[BPU.scala 406:27]
          ras_13 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_14 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'he == _T_91) begin // @[BPU.scala 406:27]
          ras_14 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[BPU.scala 344:20]
      ras_15 <= 39'h0; // @[BPU.scala 344:20]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        if (4'hf == _T_91) begin // @[BPU.scala 406:27]
          ras_15 <= _T_96; // @[BPU.scala 406:27]
        end
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 4'h0; // @[Counter.scala 60:40]
    end else if (bpuUpdateReq_valid) begin // @[BPU.scala 404:20]
      if (bpuUpdateReq_fuOpType == 7'h5c) begin // @[BPU.scala 405:45]
        value <= _T_91; // @[BPU.scala 408:16]
      end else if (bpuUpdateReq_fuOpType == 7'h5e) begin // @[BPU.scala 410:48]
        value <= _value_T_5; // @[BPU.scala 414:16]
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      rasTarget <= 39'h0; // @[Reg.scala 27:20]
    end else if (io_in_pc_valid) begin // @[Reg.scala 28:19]
      if (4'hf == value) begin // @[Reg.scala 28:23]
        rasTarget <= ras_15; // @[Reg.scala 28:23]
      end else if (4'he == value) begin // @[Reg.scala 28:23]
        rasTarget <= ras_14; // @[Reg.scala 28:23]
      end else begin
        rasTarget <= _GEN_49;
      end
    end
    if (reset) begin // @[BPU.scala 391:20]
      cnt <= 2'h0; // @[BPU.scala 391:20]
    end else if (5'h1f == bpuUpdateReq_pc[6:2]) begin // @[BPU.scala 391:20]
      cnt <= pht_31; // @[BPU.scala 391:20]
    end else if (5'h1e == bpuUpdateReq_pc[6:2]) begin // @[BPU.scala 391:20]
      cnt <= pht_30; // @[BPU.scala 391:20]
    end else if (5'h1d == bpuUpdateReq_pc[6:2]) begin // @[BPU.scala 391:20]
      cnt <= pht_29; // @[BPU.scala 391:20]
    end else begin
      cnt <= _GEN_81;
    end
    if (reset) begin // @[BPU.scala 392:25]
      reqLatch_valid <= 1'h0; // @[BPU.scala 392:25]
    end else begin
      reqLatch_valid <= bpuUpdateReq_valid; // @[BPU.scala 392:25]
    end
    if (reset) begin // @[BPU.scala 392:25]
      reqLatch_pc <= 39'h0; // @[BPU.scala 392:25]
    end else begin
      reqLatch_pc <= bpuUpdateReq_pc; // @[BPU.scala 392:25]
    end
    if (reset) begin // @[BPU.scala 392:25]
      reqLatch_actualTaken <= 1'h0; // @[BPU.scala 392:25]
    end else begin
      reqLatch_actualTaken <= bpuUpdateReq_actualTaken; // @[BPU.scala 392:25]
    end
    if (reset) begin // @[BPU.scala 392:25]
      reqLatch_fuOpType <= 7'h0; // @[BPU.scala 392:25]
    end else begin
      reqLatch_fuOpType <= bpuUpdateReq_fuOpType; // @[BPU.scala 392:25]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  pcLatch = _RAND_1[38:0];
  _RAND_2 = {1{`RANDOM}};
  REG_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pht_0 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  pht_1 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  pht_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  pht_3 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  pht_4 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  pht_5 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  pht_6 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  pht_7 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  pht_8 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  pht_9 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  pht_10 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  pht_11 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  pht_12 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  pht_13 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  pht_14 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  pht_15 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  pht_16 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  pht_17 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  pht_18 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  pht_19 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  pht_20 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  pht_21 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  pht_22 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  pht_23 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  pht_24 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  pht_25 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  pht_26 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  pht_27 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  pht_28 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  pht_29 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  pht_30 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  pht_31 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  phtTaken = _RAND_35[0:0];
  _RAND_36 = {2{`RANDOM}};
  ras_0 = _RAND_36[38:0];
  _RAND_37 = {2{`RANDOM}};
  ras_1 = _RAND_37[38:0];
  _RAND_38 = {2{`RANDOM}};
  ras_2 = _RAND_38[38:0];
  _RAND_39 = {2{`RANDOM}};
  ras_3 = _RAND_39[38:0];
  _RAND_40 = {2{`RANDOM}};
  ras_4 = _RAND_40[38:0];
  _RAND_41 = {2{`RANDOM}};
  ras_5 = _RAND_41[38:0];
  _RAND_42 = {2{`RANDOM}};
  ras_6 = _RAND_42[38:0];
  _RAND_43 = {2{`RANDOM}};
  ras_7 = _RAND_43[38:0];
  _RAND_44 = {2{`RANDOM}};
  ras_8 = _RAND_44[38:0];
  _RAND_45 = {2{`RANDOM}};
  ras_9 = _RAND_45[38:0];
  _RAND_46 = {2{`RANDOM}};
  ras_10 = _RAND_46[38:0];
  _RAND_47 = {2{`RANDOM}};
  ras_11 = _RAND_47[38:0];
  _RAND_48 = {2{`RANDOM}};
  ras_12 = _RAND_48[38:0];
  _RAND_49 = {2{`RANDOM}};
  ras_13 = _RAND_49[38:0];
  _RAND_50 = {2{`RANDOM}};
  ras_14 = _RAND_50[38:0];
  _RAND_51 = {2{`RANDOM}};
  ras_15 = _RAND_51[38:0];
  _RAND_52 = {1{`RANDOM}};
  value = _RAND_52[3:0];
  _RAND_53 = {2{`RANDOM}};
  rasTarget = _RAND_53[38:0];
  _RAND_54 = {1{`RANDOM}};
  cnt = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  reqLatch_valid = _RAND_55[0:0];
  _RAND_56 = {2{`RANDOM}};
  reqLatch_pc = _RAND_56[38:0];
  _RAND_57 = {1{`RANDOM}};
  reqLatch_actualTaken = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  reqLatch_fuOpType = _RAND_58[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_IFU_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [38:0] io_imem_req_bits_addr,
  output [81:0] io_imem_req_bits_user,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input  [81:0] io_imem_resp_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_instr,
  output [38:0] io_out_bits_pc,
  output [38:0] io_out_bits_pnpc,
  output        io_out_bits_exceptionVec_12,
  output [3:0]  io_out_bits_brIdx,
  input  [38:0] io_redirect_target,
  input         io_redirect_valid,
  output [3:0]  io_flushVec,
  input         io_ipf,
  input         flushICache,
  input         REG_6_valid,
  input  [38:0] REG_6_pc,
  input         REG_6_isMissPredict,
  input  [38:0] REG_6_actualTarget,
  input         REG_6_actualTaken,
  input  [6:0]  REG_6_fuOpType,
  input  [1:0]  REG_6_btbType,
  input         REG_6_isRVC,
  input         flushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  bp1_clock; // @[IFU.scala 325:19]
  wire  bp1_reset; // @[IFU.scala 325:19]
  wire  bp1_io_in_pc_valid; // @[IFU.scala 325:19]
  wire [38:0] bp1_io_in_pc_bits; // @[IFU.scala 325:19]
  wire [38:0] bp1_io_out_target; // @[IFU.scala 325:19]
  wire  bp1_io_out_valid; // @[IFU.scala 325:19]
  wire  bp1_io_flush; // @[IFU.scala 325:19]
  wire [2:0] bp1_io_brIdx; // @[IFU.scala 325:19]
  wire  bp1_io_crosslineJump; // @[IFU.scala 325:19]
  wire  bp1_MOUFlushICache; // @[IFU.scala 325:19]
  wire  bp1_bpuUpdateReq_valid; // @[IFU.scala 325:19]
  wire [38:0] bp1_bpuUpdateReq_pc; // @[IFU.scala 325:19]
  wire  bp1_bpuUpdateReq_isMissPredict; // @[IFU.scala 325:19]
  wire [38:0] bp1_bpuUpdateReq_actualTarget; // @[IFU.scala 325:19]
  wire  bp1_bpuUpdateReq_actualTaken; // @[IFU.scala 325:19]
  wire [6:0] bp1_bpuUpdateReq_fuOpType; // @[IFU.scala 325:19]
  wire [1:0] bp1_bpuUpdateReq_btbType; // @[IFU.scala 325:19]
  wire  bp1_bpuUpdateReq_isRVC; // @[IFU.scala 325:19]
  wire  bp1_MOUFlushTLB; // @[IFU.scala 325:19]
  reg [38:0] pc; // @[IFU.scala 321:19]
  wire  _T = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 40:37]
  wire  pcUpdate = io_redirect_valid | _T; // @[IFU.scala 322:36]
  wire [38:0] _T_3 = pc + 39'h2; // @[IFU.scala 323:28]
  wire [38:0] _T_5 = pc + 39'h4; // @[IFU.scala 323:38]
  wire [38:0] snpc = pc[1] ? _T_3 : _T_5; // @[IFU.scala 323:17]
  reg  crosslineJumpLatch; // @[IFU.scala 328:35]
  reg [38:0] crosslineJumpTarget; // @[Reg.scala 27:20]
  wire [38:0] pnpc = bp1_io_crosslineJump ? snpc : bp1_io_out_target; // @[IFU.scala 337:17]
  wire [38:0] _T_11 = bp1_io_out_valid ? pnpc : snpc; // @[IFU.scala 339:104]
  wire [38:0] _T_12 = crosslineJumpLatch ? crosslineJumpTarget : _T_11; // @[IFU.scala 339:59]
  wire [38:0] npc = io_redirect_valid ? io_redirect_target : _T_12; // @[IFU.scala 339:16]
  wire  _T_13 = bp1_io_out_valid ? 1'h0 : 1'h1; // @[IFU.scala 340:114]
  wire  _T_15 = crosslineJumpLatch ? 1'h0 : bp1_io_crosslineJump | _T_13; // @[IFU.scala 340:54]
  wire  npcIsSeq = io_redirect_valid ? 1'h0 : _T_15; // @[IFU.scala 340:21]
  wire [2:0] lo = io_redirect_valid ? 3'h0 : bp1_io_brIdx; // @[IFU.scala 348:29]
  wire [37:0] hi = pc[38:1]; // @[IFU.scala 369:39]
  wire [42:0] hi_1 = {npcIsSeq,lo,npc}; // @[Cat.scala 30:58]
  wire  _T_40 = io_imem_resp_ready & io_imem_resp_valid; // @[Decoupled.scala 40:37]
  reg  REG_3; // @[StopWatch.scala 24:20]
  wire  _GEN_3 = io_imem_req_valid | REG_3; // @[StopWatch.scala 30:20 StopWatch.scala 30:24 StopWatch.scala 24:20]
  wire  _T_41 = |io_flushVec; // @[IFU.scala 393:37]
  ysyx_210000_BPU_inorder bp1 ( // @[IFU.scala 325:19]
    .clock(bp1_clock),
    .reset(bp1_reset),
    .io_in_pc_valid(bp1_io_in_pc_valid),
    .io_in_pc_bits(bp1_io_in_pc_bits),
    .io_out_target(bp1_io_out_target),
    .io_out_valid(bp1_io_out_valid),
    .io_flush(bp1_io_flush),
    .io_brIdx(bp1_io_brIdx),
    .io_crosslineJump(bp1_io_crosslineJump),
    .MOUFlushICache(bp1_MOUFlushICache),
    .bpuUpdateReq_valid(bp1_bpuUpdateReq_valid),
    .bpuUpdateReq_pc(bp1_bpuUpdateReq_pc),
    .bpuUpdateReq_isMissPredict(bp1_bpuUpdateReq_isMissPredict),
    .bpuUpdateReq_actualTarget(bp1_bpuUpdateReq_actualTarget),
    .bpuUpdateReq_actualTaken(bp1_bpuUpdateReq_actualTaken),
    .bpuUpdateReq_fuOpType(bp1_bpuUpdateReq_fuOpType),
    .bpuUpdateReq_btbType(bp1_bpuUpdateReq_btbType),
    .bpuUpdateReq_isRVC(bp1_bpuUpdateReq_isRVC),
    .MOUFlushTLB(bp1_MOUFlushTLB)
  );
  assign io_imem_req_valid = io_out_ready; // @[IFU.scala 371:21]
  assign io_imem_req_bits_addr = {hi,1'h0}; // @[Cat.scala 30:58]
  assign io_imem_req_bits_user = {hi_1,pc}; // @[Cat.scala 30:58]
  assign io_imem_resp_ready = io_out_ready | io_flushVec[0]; // @[IFU.scala 373:38]
  assign io_out_valid = io_imem_resp_valid & ~io_flushVec[0]; // @[IFU.scala 390:38]
  assign io_out_bits_instr = io_imem_resp_bits_rdata; // @[IFU.scala 383:21]
  assign io_out_bits_pc = io_imem_resp_bits_user[38:0]; // @[IFU.scala 385:24]
  assign io_out_bits_pnpc = io_imem_resp_bits_user[77:39]; // @[IFU.scala 386:26]
  assign io_out_bits_exceptionVec_12 = io_ipf; // @[IFU.scala 389:44]
  assign io_out_bits_brIdx = io_imem_resp_bits_user[81:78]; // @[IFU.scala 387:27]
  assign io_flushVec = io_redirect_valid ? 4'hf : 4'h0; // @[IFU.scala 366:21]
  assign bp1_clock = clock;
  assign bp1_reset = reset;
  assign bp1_io_in_pc_valid = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 40:37]
  assign bp1_io_in_pc_bits = io_redirect_valid ? io_redirect_target : _T_12; // @[IFU.scala 339:16]
  assign bp1_io_flush = io_redirect_valid; // @[IFU.scala 357:16]
  assign bp1_MOUFlushICache = flushICache;
  assign bp1_bpuUpdateReq_valid = REG_6_valid;
  assign bp1_bpuUpdateReq_pc = REG_6_pc;
  assign bp1_bpuUpdateReq_isMissPredict = REG_6_isMissPredict;
  assign bp1_bpuUpdateReq_actualTarget = REG_6_actualTarget;
  assign bp1_bpuUpdateReq_actualTaken = REG_6_actualTaken;
  assign bp1_bpuUpdateReq_fuOpType = REG_6_fuOpType;
  assign bp1_bpuUpdateReq_btbType = REG_6_btbType;
  assign bp1_bpuUpdateReq_isRVC = REG_6_isRVC;
  assign bp1_MOUFlushTLB = flushTLB;
  always @(posedge clock) begin
    if (reset) begin // @[IFU.scala 321:19]
      pc <= 39'h30000000; // @[IFU.scala 321:19]
    end else if (pcUpdate) begin // @[IFU.scala 359:19]
      if (io_redirect_valid) begin // @[IFU.scala 339:16]
        pc <= io_redirect_target;
      end else if (crosslineJumpLatch) begin // @[IFU.scala 339:59]
        pc <= crosslineJumpTarget;
      end else begin
        pc <= _T_11;
      end
    end
    if (reset) begin // @[IFU.scala 328:35]
      crosslineJumpLatch <= 1'h0; // @[IFU.scala 328:35]
    end else if (pcUpdate | bp1_io_flush) begin // @[IFU.scala 329:34]
      if (bp1_io_flush) begin // @[IFU.scala 330:30]
        crosslineJumpLatch <= 1'h0;
      end else begin
        crosslineJumpLatch <= bp1_io_crosslineJump & ~crosslineJumpLatch;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      crosslineJumpTarget <= 39'h0; // @[Reg.scala 27:20]
    end else if (bp1_io_crosslineJump) begin // @[Reg.scala 28:19]
      crosslineJumpTarget <= bp1_io_out_target; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_3 <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (_T_40) begin // @[StopWatch.scala 31:19]
      REG_3 <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      REG_3 <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[38:0];
  _RAND_1 = {1{`RANDOM}};
  crosslineJumpLatch = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  crosslineJumpTarget = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  REG_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_NaiveRVCAlignBuffer(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_instr,
  input  [38:0] io_in_bits_pc,
  input  [38:0] io_in_bits_pnpc,
  input         io_in_bits_exceptionVec_12,
  input  [3:0]  io_in_bits_brIdx,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_instr,
  output [38:0] io_out_bits_pc,
  output [38:0] io_out_bits_pnpc,
  output        io_out_bits_exceptionVec_12,
  output [3:0]  io_out_bits_brIdx,
  output        io_out_bits_crossPageIPFFix,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[NaiveIBF.scala 39:22]
  wire  _T_76 = state == 2'h2; // @[NaiveIBF.scala 90:23]
  wire  _T_77 = state == 2'h3; // @[NaiveIBF.scala 90:47]
  wire [79:0] instIn = {16'h0,io_in_bits_instr}; // @[Cat.scala 30:58]
  wire [15:0] hi_1 = instIn[15:0]; // @[NaiveIBF.scala 90:80]
  reg [15:0] specialInstR; // @[NaiveIBF.scala 66:29]
  wire [31:0] _T_79 = {hi_1,specialInstR}; // @[Cat.scala 30:58]
  wire  _T_1 = state == 2'h0; // @[NaiveIBF.scala 41:28]
  reg [2:0] pcOffsetR; // @[NaiveIBF.scala 40:26]
  wire [2:0] pcOffset = state == 2'h0 ? io_in_bits_pc[2:0] : pcOffsetR; // @[NaiveIBF.scala 41:21]
  wire  _T_84 = 3'h0 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_88 = _T_84 ? instIn[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire  _T_85 = 3'h2 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_89 = _T_85 ? instIn[47:16] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_92 = _T_88 | _T_89; // @[Mux.scala 27:72]
  wire  _T_86 = 3'h4 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_90 = _T_86 ? instIn[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_93 = _T_92 | _T_90; // @[Mux.scala 27:72]
  wire  _T_87 = 3'h6 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_91 = _T_87 ? instIn[79:48] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_94 = _T_93 | _T_91; // @[Mux.scala 27:72]
  wire [31:0] instr = state == 2'h2 | state == 2'h3 ? _T_79 : _T_94; // @[NaiveIBF.scala 90:15]
  wire  isRVC = instr[1:0] != 2'h3; // @[NaiveIBF.scala 34:26]
  wire  _T_3 = pcOffset == 3'h0; // @[NaiveIBF.scala 48:28]
  wire  _T_4 = ~isRVC; // @[NaiveIBF.scala 48:40]
  wire  _T_8 = pcOffset == 3'h4; // @[NaiveIBF.scala 48:72]
  wire  _T_14 = pcOffset == 3'h2; // @[NaiveIBF.scala 48:116]
  wire  _T_19 = pcOffset == 3'h6; // @[NaiveIBF.scala 48:159]
  wire  rvcFinish = pcOffset == 3'h0 & (~isRVC | io_in_bits_brIdx[0]) | pcOffset == 3'h4 & (~isRVC | io_in_bits_brIdx[0]
    ) | pcOffset == 3'h2 & (isRVC | io_in_bits_brIdx[1]) | pcOffset == 3'h6 & isRVC; // @[NaiveIBF.scala 48:147]
  wire  _T_34 = _T_14 & _T_4; // @[NaiveIBF.scala 51:122]
  wire  _T_36 = ~io_in_bits_brIdx[1]; // @[NaiveIBF.scala 51:135]
  wire  rvcNext = _T_3 & (isRVC & ~io_in_bits_brIdx[0]) | _T_8 & (isRVC & ~io_in_bits_brIdx[0]) | _T_14 & _T_4 & ~
    io_in_bits_brIdx[1]; // @[NaiveIBF.scala 51:102]
  wire  _T_40 = _T_19 & _T_4; // @[NaiveIBF.scala 52:37]
  wire  rvcSpecial = _T_19 & _T_4 & ~io_in_bits_brIdx[2]; // @[NaiveIBF.scala 52:47]
  wire  rvcSpecialJump = _T_40 & io_in_bits_brIdx[2]; // @[NaiveIBF.scala 53:51]
  wire  pnpcIsSeq = io_in_bits_brIdx[3]; // @[NaiveIBF.scala 54:24]
  wire  _T_49 = _T_1 | state == 2'h1; // @[NaiveIBF.scala 57:36]
  wire  flushIFU = (_T_1 | state == 2'h1) & rvcSpecial & io_in_valid & ~pnpcIsSeq; // @[NaiveIBF.scala 57:87]
  wire  loadNextInstline = _T_49 & (rvcSpecial | rvcSpecialJump) & io_in_valid & pnpcIsSeq; // @[NaiveIBF.scala 60:115]
  reg [38:0] specialPCR; // @[NaiveIBF.scala 64:27]
  reg [38:0] specialNPCR; // @[NaiveIBF.scala 65:28]
  reg  specialIPFR; // @[NaiveIBF.scala 67:28]
  wire [35:0] hi = io_in_bits_pc[38:3]; // @[NaiveIBF.scala 68:37]
  wire  rvcForceLoadNext = _T_34 & io_in_bits_pnpc[2:0] == 3'h4 & _T_36; // @[NaiveIBF.scala 69:86]
  wire  _T_97 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_98 = rvcFinish | rvcNext; // @[NaiveIBF.scala 100:28]
  wire  _T_99 = rvcFinish | rvcForceLoadNext; // @[NaiveIBF.scala 101:28]
  wire [38:0] _T_101 = io_in_bits_pc + 39'h2; // @[NaiveIBF.scala 103:76]
  wire [38:0] _T_103 = io_in_bits_pc + 39'h4; // @[NaiveIBF.scala 103:95]
  wire [38:0] _T_104 = isRVC ? _T_101 : _T_103; // @[NaiveIBF.scala 103:55]
  wire [38:0] _T_105 = rvcFinish ? io_in_bits_pnpc : _T_104; // @[NaiveIBF.scala 103:23]
  wire  _T_106 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_0 = _T_106 & rvcFinish ? 2'h0 : state; // @[NaiveIBF.scala 104:41 NaiveIBF.scala 104:48 NaiveIBF.scala 39:22]
  wire [2:0] _T_110 = isRVC ? 3'h2 : 3'h4; // @[NaiveIBF.scala 107:38]
  wire [2:0] _T_112 = pcOffset + _T_110; // @[NaiveIBF.scala 107:33]
  wire [1:0] _GEN_1 = _T_106 & rvcNext ? 2'h1 : _GEN_0; // @[NaiveIBF.scala 105:39 NaiveIBF.scala 106:17]
  wire [2:0] _GEN_2 = _T_106 & rvcNext ? _T_112 : pcOffsetR; // @[NaiveIBF.scala 105:39 NaiveIBF.scala 107:21 NaiveIBF.scala 40:26]
  wire [1:0] _GEN_3 = rvcSpecial & io_in_valid ? 2'h2 : _GEN_1; // @[NaiveIBF.scala 109:40 NaiveIBF.scala 110:17]
  wire  _T_115 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [38:0] _T_118 = {hi,pcOffsetR}; // @[Cat.scala 30:58]
  wire  _T_134 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_138 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [38:0] _GEN_27 = _T_138 ? specialPCR : 39'h0; // @[Conditional.scala 39:67 NaiveIBF.scala 161:15]
  wire [38:0] _GEN_32 = _T_134 ? specialPCR : _GEN_27; // @[Conditional.scala 39:67 NaiveIBF.scala 149:15]
  wire [38:0] _GEN_40 = _T_115 ? _T_118 : _GEN_32; // @[Conditional.scala 39:67 NaiveIBF.scala 126:15]
  wire [38:0] pcOut = _T_97 ? io_in_bits_pc : _GEN_40; // @[Conditional.scala 40:58 NaiveIBF.scala 102:15]
  wire [38:0] _GEN_4 = rvcSpecial & io_in_valid ? pcOut : specialPCR; // @[NaiveIBF.scala 109:40 NaiveIBF.scala 111:22 NaiveIBF.scala 64:27]
  wire [15:0] _GEN_5 = rvcSpecial & io_in_valid ? io_in_bits_instr[63:48] : specialInstR; // @[NaiveIBF.scala 109:40 NaiveIBF.scala 112:24 NaiveIBF.scala 66:29]
  wire  _GEN_6 = rvcSpecial & io_in_valid ? io_in_bits_exceptionVec_12 : specialIPFR; // @[NaiveIBF.scala 109:40 NaiveIBF.scala 113:23 NaiveIBF.scala 67:28]
  wire [1:0] _GEN_7 = rvcSpecialJump & io_in_valid ? 2'h3 : _GEN_3; // @[NaiveIBF.scala 115:44 NaiveIBF.scala 116:17]
  wire [38:0] _GEN_8 = rvcSpecialJump & io_in_valid ? pcOut : _GEN_4; // @[NaiveIBF.scala 115:44 NaiveIBF.scala 117:22]
  wire [38:0] _GEN_9 = rvcSpecialJump & io_in_valid ? io_in_bits_pnpc : specialNPCR; // @[NaiveIBF.scala 115:44 NaiveIBF.scala 118:23 NaiveIBF.scala 65:28]
  wire [15:0] _GEN_10 = rvcSpecialJump & io_in_valid ? io_in_bits_instr[63:48] : _GEN_5; // @[NaiveIBF.scala 115:44 NaiveIBF.scala 119:24]
  wire  _GEN_11 = rvcSpecialJump & io_in_valid ? io_in_bits_exceptionVec_12 : _GEN_6; // @[NaiveIBF.scala 115:44 NaiveIBF.scala 120:23]
  wire [38:0] _T_120 = pcOut + 39'h2; // @[NaiveIBF.scala 127:68]
  wire [38:0] _T_122 = pcOut + 39'h4; // @[NaiveIBF.scala 127:79]
  wire [38:0] _T_123 = isRVC ? _T_120 : _T_122; // @[NaiveIBF.scala 127:55]
  wire [38:0] _T_124 = rvcFinish ? io_in_bits_pnpc : _T_123; // @[NaiveIBF.scala 127:23]
  wire [38:0] _T_136 = specialPCR + 39'h4; // @[NaiveIBF.scala 150:31]
  wire [1:0] _GEN_24 = _T_106 ? 2'h1 : state; // @[NaiveIBF.scala 154:28 NaiveIBF.scala 155:17 NaiveIBF.scala 39:22]
  wire [2:0] _GEN_25 = _T_106 ? 3'h2 : pcOffsetR; // @[NaiveIBF.scala 154:28 NaiveIBF.scala 156:21 NaiveIBF.scala 40:26]
  wire [1:0] _GEN_26 = _T_106 ? 2'h0 : state; // @[NaiveIBF.scala 166:28 NaiveIBF.scala 167:17 NaiveIBF.scala 39:22]
  wire [38:0] _GEN_28 = _T_138 ? specialNPCR : 39'h0; // @[Conditional.scala 39:67 NaiveIBF.scala 162:17]
  wire  _GEN_29 = _T_138 & io_in_valid; // @[Conditional.scala 39:67 NaiveIBF.scala 164:15]
  wire [1:0] _GEN_31 = _T_138 ? _GEN_26 : state; // @[Conditional.scala 39:67 NaiveIBF.scala 39:22]
  wire [38:0] _GEN_33 = _T_134 ? _T_136 : _GEN_28; // @[Conditional.scala 39:67 NaiveIBF.scala 150:17]
  wire  _GEN_34 = _T_134 ? io_in_valid : _GEN_29; // @[Conditional.scala 39:67 NaiveIBF.scala 152:15]
  wire  _GEN_35 = _T_134 ? 1'h0 : _T_138; // @[Conditional.scala 39:67 NaiveIBF.scala 153:15]
  wire [1:0] _GEN_36 = _T_134 ? _GEN_24 : _GEN_31; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_37 = _T_134 ? _GEN_25 : pcOffsetR; // @[Conditional.scala 39:67 NaiveIBF.scala 40:26]
  wire  _GEN_38 = _T_115 ? _T_98 : _GEN_34; // @[Conditional.scala 39:67 NaiveIBF.scala 124:15]
  wire  _GEN_39 = _T_115 ? _T_99 : _GEN_35; // @[Conditional.scala 39:67 NaiveIBF.scala 125:15]
  wire [38:0] _GEN_41 = _T_115 ? _T_124 : _GEN_33; // @[Conditional.scala 39:67 NaiveIBF.scala 127:17]
  wire  canGo = _T_97 ? rvcFinish | rvcNext : _GEN_38; // @[Conditional.scala 40:58 NaiveIBF.scala 100:15]
  wire  canIn = _T_97 ? rvcFinish | rvcForceLoadNext : _GEN_39; // @[Conditional.scala 40:58 NaiveIBF.scala 101:15]
  wire [38:0] pnpcOut = _T_97 ? _T_105 : _GEN_41; // @[Conditional.scala 40:58 NaiveIBF.scala 103:17]
  wire  _T_150 = pnpcOut == _T_122 & _T_4 | pnpcOut == _T_120 & isRVC ? 1'h0 : 1'h1; // @[NaiveIBF.scala 185:27]
  wire  _T_159 = _T_77 | _T_76; // @[NaiveIBF.scala 191:133]
  assign io_in_ready = ~io_in_valid | _T_106 & canIn | loadNextInstline; // @[NaiveIBF.scala 188:60]
  assign io_out_valid = io_in_valid & canGo; // @[NaiveIBF.scala 187:31]
  assign io_out_bits_instr = {{32'd0}, instr}; // @[NaiveIBF.scala 90:15]
  assign io_out_bits_pc = _T_97 ? io_in_bits_pc : _GEN_40; // @[Conditional.scala 40:58 NaiveIBF.scala 102:15]
  assign io_out_bits_pnpc = _T_97 ? _T_105 : _GEN_41; // @[Conditional.scala 40:58 NaiveIBF.scala 103:17]
  assign io_out_bits_exceptionVec_12 = io_in_bits_exceptionVec_12 | specialIPFR & (_T_77 | _T_76); // @[NaiveIBF.scala 191:87]
  assign io_out_bits_brIdx = {{3'd0}, _T_150}; // @[NaiveIBF.scala 185:27]
  assign io_out_bits_crossPageIPFFix = io_in_bits_exceptionVec_12 & _T_159 & ~specialIPFR; // @[NaiveIBF.scala 192:130]
  always @(posedge clock) begin
    if (reset) begin // @[NaiveIBF.scala 39:22]
      state <= 2'h0; // @[NaiveIBF.scala 39:22]
    end else if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (_T_97) begin // @[Conditional.scala 40:58]
        state <= _GEN_7;
      end else if (_T_115) begin // @[Conditional.scala 39:67]
        state <= _GEN_7;
      end else begin
        state <= _GEN_36;
      end
    end else begin
      state <= 2'h0; // @[NaiveIBF.scala 172:11]
    end
    if (reset) begin // @[NaiveIBF.scala 66:29]
      specialInstR <= 16'h0; // @[NaiveIBF.scala 66:29]
    end else if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (_T_97) begin // @[Conditional.scala 40:58]
        specialInstR <= _GEN_10;
      end else if (_T_115) begin // @[Conditional.scala 39:67]
        specialInstR <= _GEN_10;
      end
    end
    if (reset) begin // @[NaiveIBF.scala 40:26]
      pcOffsetR <= 3'h0; // @[NaiveIBF.scala 40:26]
    end else if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (_T_97) begin // @[Conditional.scala 40:58]
        pcOffsetR <= _GEN_2;
      end else if (_T_115) begin // @[Conditional.scala 39:67]
        pcOffsetR <= _GEN_2;
      end else begin
        pcOffsetR <= _GEN_37;
      end
    end
    if (reset) begin // @[NaiveIBF.scala 64:27]
      specialPCR <= 39'h0; // @[NaiveIBF.scala 64:27]
    end else if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (_T_97) begin // @[Conditional.scala 40:58]
        specialPCR <= _GEN_8;
      end else if (_T_115) begin // @[Conditional.scala 39:67]
        specialPCR <= _GEN_8;
      end
    end
    if (reset) begin // @[NaiveIBF.scala 65:28]
      specialNPCR <= 39'h0; // @[NaiveIBF.scala 65:28]
    end else if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (_T_97) begin // @[Conditional.scala 40:58]
        specialNPCR <= _GEN_9;
      end else if (_T_115) begin // @[Conditional.scala 39:67]
        specialNPCR <= _GEN_9;
      end
    end
    if (reset) begin // @[NaiveIBF.scala 67:28]
      specialIPFR <= 1'h0; // @[NaiveIBF.scala 67:28]
    end else if (~io_flush) begin // @[NaiveIBF.scala 97:18]
      if (_T_97) begin // @[Conditional.scala 40:58]
        specialIPFR <= _GEN_11;
      end else if (_T_115) begin // @[Conditional.scala 39:67]
        specialIPFR <= _GEN_11;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~flushIFU | reset)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NaiveIBF.scala:59 assert(!flushIFU)\n"); // @[NaiveIBF.scala 59:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~flushIFU | reset)) begin
          $fatal; // @[NaiveIBF.scala 59:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  specialInstR = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  pcOffsetR = _RAND_2[2:0];
  _RAND_3 = {2{`RANDOM}};
  specialPCR = _RAND_3[38:0];
  _RAND_4 = {2{`RANDOM}};
  specialNPCR = _RAND_4[38:0];
  _RAND_5 = {1{`RANDOM}};
  specialIPFR = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_Decoder(
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_instr,
  input  [38:0] io_in_bits_pc,
  input  [38:0] io_in_bits_pnpc,
  input         io_in_bits_exceptionVec_12,
  input  [3:0]  io_in_bits_brIdx,
  input         io_in_bits_crossPageIPFFix,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_cf_instr,
  output [38:0] io_out_bits_cf_pc,
  output [38:0] io_out_bits_cf_pnpc,
  output        io_out_bits_cf_exceptionVec_1,
  output        io_out_bits_cf_exceptionVec_2,
  output        io_out_bits_cf_exceptionVec_12,
  output        io_out_bits_cf_intrVec_0,
  output        io_out_bits_cf_intrVec_1,
  output        io_out_bits_cf_intrVec_2,
  output        io_out_bits_cf_intrVec_3,
  output        io_out_bits_cf_intrVec_4,
  output        io_out_bits_cf_intrVec_5,
  output        io_out_bits_cf_intrVec_6,
  output        io_out_bits_cf_intrVec_7,
  output        io_out_bits_cf_intrVec_8,
  output        io_out_bits_cf_intrVec_9,
  output        io_out_bits_cf_intrVec_10,
  output        io_out_bits_cf_intrVec_11,
  output [3:0]  io_out_bits_cf_brIdx,
  output        io_out_bits_cf_crossPageIPFFix,
  output        io_out_bits_ctrl_src1Type,
  output        io_out_bits_ctrl_src2Type,
  output [2:0]  io_out_bits_ctrl_fuType,
  output [6:0]  io_out_bits_ctrl_fuOpType,
  output [4:0]  io_out_bits_ctrl_rfSrc1,
  output [4:0]  io_out_bits_ctrl_rfSrc2,
  output        io_out_bits_ctrl_rfWen,
  output [4:0]  io_out_bits_ctrl_rfDest,
  output [63:0] io_out_bits_data_imm,
  input         DTLBENABLE,
  input  [11:0] intrVecIDU
);
  wire [63:0] _T = io_in_bits_instr & 64'h707f; // @[Lookup.scala 31:38]
  wire  _T_1 = 64'h13 == _T; // @[Lookup.scala 31:38]
  wire [63:0] _T_2 = io_in_bits_instr & 64'hfc00707f; // @[Lookup.scala 31:38]
  wire  _T_3 = 64'h1013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_5 = 64'h2013 == _T; // @[Lookup.scala 31:38]
  wire  _T_7 = 64'h3013 == _T; // @[Lookup.scala 31:38]
  wire  _T_9 = 64'h4013 == _T; // @[Lookup.scala 31:38]
  wire  _T_11 = 64'h5013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_13 = 64'h6013 == _T; // @[Lookup.scala 31:38]
  wire  _T_15 = 64'h7013 == _T; // @[Lookup.scala 31:38]
  wire  _T_17 = 64'h40005013 == _T_2; // @[Lookup.scala 31:38]
  wire [63:0] _T_18 = io_in_bits_instr & 64'hfe00707f; // @[Lookup.scala 31:38]
  wire  _T_19 = 64'h33 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_21 = 64'h1033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_23 = 64'h2033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_25 = 64'h3033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_27 = 64'h4033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_29 = 64'h5033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_31 = 64'h6033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_33 = 64'h7033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_35 = 64'h40000033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_37 = 64'h40005033 == _T_18; // @[Lookup.scala 31:38]
  wire [63:0] _T_38 = io_in_bits_instr & 64'h7f; // @[Lookup.scala 31:38]
  wire  _T_39 = 64'h17 == _T_38; // @[Lookup.scala 31:38]
  wire  _T_41 = 64'h37 == _T_38; // @[Lookup.scala 31:38]
  wire  _T_43 = 64'h6f == _T_38; // @[Lookup.scala 31:38]
  wire  _T_45 = 64'h67 == _T; // @[Lookup.scala 31:38]
  wire  _T_47 = 64'h63 == _T; // @[Lookup.scala 31:38]
  wire  _T_49 = 64'h1063 == _T; // @[Lookup.scala 31:38]
  wire  _T_51 = 64'h4063 == _T; // @[Lookup.scala 31:38]
  wire  _T_53 = 64'h5063 == _T; // @[Lookup.scala 31:38]
  wire  _T_55 = 64'h6063 == _T; // @[Lookup.scala 31:38]
  wire  _T_57 = 64'h7063 == _T; // @[Lookup.scala 31:38]
  wire  _T_59 = 64'h3 == _T; // @[Lookup.scala 31:38]
  wire  _T_61 = 64'h1003 == _T; // @[Lookup.scala 31:38]
  wire  _T_63 = 64'h2003 == _T; // @[Lookup.scala 31:38]
  wire  _T_65 = 64'h4003 == _T; // @[Lookup.scala 31:38]
  wire  _T_67 = 64'h5003 == _T; // @[Lookup.scala 31:38]
  wire  _T_69 = 64'h23 == _T; // @[Lookup.scala 31:38]
  wire  _T_71 = 64'h1023 == _T; // @[Lookup.scala 31:38]
  wire  _T_73 = 64'h2023 == _T; // @[Lookup.scala 31:38]
  wire  _T_75 = 64'h1b == _T; // @[Lookup.scala 31:38]
  wire  _T_77 = 64'h101b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_79 = 64'h501b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_81 = 64'h4000501b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_83 = 64'h103b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_85 = 64'h503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_87 = 64'h4000503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_89 = 64'h3b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_91 = 64'h4000003b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_93 = 64'h6003 == _T; // @[Lookup.scala 31:38]
  wire  _T_95 = 64'h3003 == _T; // @[Lookup.scala 31:38]
  wire  _T_97 = 64'h3023 == _T; // @[Lookup.scala 31:38]
  wire  _T_99 = 64'h6b == _T; // @[Lookup.scala 31:38]
  wire  _T_101 = 64'h2000033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_103 = 64'h2001033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_105 = 64'h2002033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_107 = 64'h2003033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_109 = 64'h2004033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_111 = 64'h2005033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_113 = 64'h2006033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_115 = 64'h2007033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_117 = 64'h200003b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_119 = 64'h200403b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_121 = 64'h200503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_123 = 64'h200603b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_125 = 64'h200703b == _T_18; // @[Lookup.scala 31:38]
  wire [63:0] _T_126 = io_in_bits_instr & 64'hffffffff; // @[Lookup.scala 31:38]
  wire  _T_127 = 64'h0 == _T_126; // @[Lookup.scala 31:38]
  wire [63:0] _T_128 = io_in_bits_instr & 64'he003; // @[Lookup.scala 31:38]
  wire  _T_129 = 64'h0 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_131 = 64'h4000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_133 = 64'h6000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_135 = 64'hc000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_137 = 64'he000 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_138 = io_in_bits_instr & 64'hef83; // @[Lookup.scala 31:38]
  wire  _T_139 = 64'h1 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_141 = 64'h1 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_143 = 64'h2001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_145 = 64'h4001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_147 = 64'h6101 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_149 = 64'h6001 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_150 = io_in_bits_instr & 64'hec03; // @[Lookup.scala 31:38]
  wire  _T_151 = 64'h8001 == _T_150; // @[Lookup.scala 31:38]
  wire  _T_153 = 64'h8401 == _T_150; // @[Lookup.scala 31:38]
  wire  _T_155 = 64'h8801 == _T_150; // @[Lookup.scala 31:38]
  wire [63:0] _T_156 = io_in_bits_instr & 64'hfc63; // @[Lookup.scala 31:38]
  wire  _T_157 = 64'h8c01 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_159 = 64'h8c21 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_161 = 64'h8c41 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_163 = 64'h8c61 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_165 = 64'h9c01 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_167 = 64'h9c21 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_169 = 64'ha001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_171 = 64'hc001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_173 = 64'he001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_175 = 64'h2 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_177 = 64'h4002 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_179 = 64'h6002 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_180 = io_in_bits_instr & 64'hf07f; // @[Lookup.scala 31:38]
  wire  _T_181 = 64'h8002 == _T_180; // @[Lookup.scala 31:38]
  wire [63:0] _T_182 = io_in_bits_instr & 64'hf003; // @[Lookup.scala 31:38]
  wire  _T_183 = 64'h8002 == _T_182; // @[Lookup.scala 31:38]
  wire [63:0] _T_184 = io_in_bits_instr & 64'hffff; // @[Lookup.scala 31:38]
  wire  _T_185 = 64'h9002 == _T_184; // @[Lookup.scala 31:38]
  wire  _T_187 = 64'h9002 == _T_180; // @[Lookup.scala 31:38]
  wire  _T_189 = 64'h9002 == _T_182; // @[Lookup.scala 31:38]
  wire  _T_191 = 64'hc002 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_193 = 64'he002 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_195 = 64'h73 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_197 = 64'h100073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_199 = 64'h30200073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_201 = 64'hf == _T; // @[Lookup.scala 31:38]
  wire  _T_203 = 64'h10500073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_205 = 64'h10200073 == _T_126; // @[Lookup.scala 31:38]
  wire [63:0] _T_206 = io_in_bits_instr & 64'hfe007fff; // @[Lookup.scala 31:38]
  wire  _T_207 = 64'h12000073 == _T_206; // @[Lookup.scala 31:38]
  wire  _T_209 = 64'h200073 == _T_126; // @[Lookup.scala 31:38]
  wire [63:0] _T_210 = io_in_bits_instr & 64'hf9f0707f; // @[Lookup.scala 31:38]
  wire  _T_211 = 64'h1000302f == _T_210; // @[Lookup.scala 31:38]
  wire  _T_213 = 64'h1000202f == _T_210; // @[Lookup.scala 31:38]
  wire [63:0] _T_214 = io_in_bits_instr & 64'hf800707f; // @[Lookup.scala 31:38]
  wire  _T_215 = 64'h1800302f == _T_214; // @[Lookup.scala 31:38]
  wire  _T_217 = 64'h1800202f == _T_214; // @[Lookup.scala 31:38]
  wire [63:0] _T_218 = io_in_bits_instr & 64'hf800607f; // @[Lookup.scala 31:38]
  wire  _T_219 = 64'h800202f == _T_218; // @[Lookup.scala 31:38]
  wire  _T_221 = 64'h202f == _T_218; // @[Lookup.scala 31:38]
  wire  _T_223 = 64'h2000202f == _T_218; // @[Lookup.scala 31:38]
  wire  _T_225 = 64'h6000202f == _T_218; // @[Lookup.scala 31:38]
  wire  _T_227 = 64'h4000202f == _T_218; // @[Lookup.scala 31:38]
  wire  _T_229 = 64'h8000202f == _T_218; // @[Lookup.scala 31:38]
  wire  _T_231 = 64'ha000202f == _T_218; // @[Lookup.scala 31:38]
  wire  _T_233 = 64'hc000202f == _T_218; // @[Lookup.scala 31:38]
  wire  _T_235 = 64'he000202f == _T_218; // @[Lookup.scala 31:38]
  wire  _T_237 = 64'h1073 == _T; // @[Lookup.scala 31:38]
  wire  _T_239 = 64'h2073 == _T; // @[Lookup.scala 31:38]
  wire  _T_241 = 64'h3073 == _T; // @[Lookup.scala 31:38]
  wire  _T_243 = 64'h5073 == _T; // @[Lookup.scala 31:38]
  wire  _T_245 = 64'h6073 == _T; // @[Lookup.scala 31:38]
  wire  _T_247 = 64'h7073 == _T; // @[Lookup.scala 31:38]
  wire  _T_249 = 64'h100f == _T_126; // @[Lookup.scala 31:38]
  wire  _T_251 = 64'h700b == _T; // @[Lookup.scala 31:38]
  wire [2:0] _T_252 = _T_251 ? 3'h4 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_253 = _T_249 ? 3'h1 : _T_252; // @[Lookup.scala 33:37]
  wire [2:0] _T_254 = _T_247 ? 3'h4 : _T_253; // @[Lookup.scala 33:37]
  wire [2:0] _T_255 = _T_245 ? 3'h4 : _T_254; // @[Lookup.scala 33:37]
  wire [2:0] _T_256 = _T_243 ? 3'h4 : _T_255; // @[Lookup.scala 33:37]
  wire [2:0] _T_257 = _T_241 ? 3'h4 : _T_256; // @[Lookup.scala 33:37]
  wire [2:0] _T_258 = _T_239 ? 3'h4 : _T_257; // @[Lookup.scala 33:37]
  wire [2:0] _T_259 = _T_237 ? 3'h4 : _T_258; // @[Lookup.scala 33:37]
  wire [2:0] _T_260 = _T_235 ? 3'h5 : _T_259; // @[Lookup.scala 33:37]
  wire [2:0] _T_261 = _T_233 ? 3'h5 : _T_260; // @[Lookup.scala 33:37]
  wire [2:0] _T_262 = _T_231 ? 3'h5 : _T_261; // @[Lookup.scala 33:37]
  wire [2:0] _T_263 = _T_229 ? 3'h5 : _T_262; // @[Lookup.scala 33:37]
  wire [2:0] _T_264 = _T_227 ? 3'h5 : _T_263; // @[Lookup.scala 33:37]
  wire [2:0] _T_265 = _T_225 ? 3'h5 : _T_264; // @[Lookup.scala 33:37]
  wire [2:0] _T_266 = _T_223 ? 3'h5 : _T_265; // @[Lookup.scala 33:37]
  wire [2:0] _T_267 = _T_221 ? 3'h5 : _T_266; // @[Lookup.scala 33:37]
  wire [2:0] _T_268 = _T_219 ? 3'h5 : _T_267; // @[Lookup.scala 33:37]
  wire [3:0] _T_269 = _T_217 ? 4'hf : {{1'd0}, _T_268}; // @[Lookup.scala 33:37]
  wire [3:0] _T_270 = _T_215 ? 4'hf : _T_269; // @[Lookup.scala 33:37]
  wire [3:0] _T_271 = _T_213 ? 4'h4 : _T_270; // @[Lookup.scala 33:37]
  wire [3:0] _T_272 = _T_211 ? 4'h4 : _T_271; // @[Lookup.scala 33:37]
  wire [3:0] _T_273 = _T_209 ? 4'h4 : _T_272; // @[Lookup.scala 33:37]
  wire [3:0] _T_274 = _T_207 ? 4'h5 : _T_273; // @[Lookup.scala 33:37]
  wire [3:0] _T_275 = _T_205 ? 4'h4 : _T_274; // @[Lookup.scala 33:37]
  wire [3:0] _T_276 = _T_203 ? 4'h4 : _T_275; // @[Lookup.scala 33:37]
  wire [3:0] _T_277 = _T_201 ? 4'h2 : _T_276; // @[Lookup.scala 33:37]
  wire [3:0] _T_278 = _T_199 ? 4'h4 : _T_277; // @[Lookup.scala 33:37]
  wire [3:0] _T_279 = _T_197 ? 4'h4 : _T_278; // @[Lookup.scala 33:37]
  wire [3:0] _T_280 = _T_195 ? 4'h4 : _T_279; // @[Lookup.scala 33:37]
  wire [3:0] _T_281 = _T_193 ? 4'h2 : _T_280; // @[Lookup.scala 33:37]
  wire [3:0] _T_282 = _T_191 ? 4'h2 : _T_281; // @[Lookup.scala 33:37]
  wire [3:0] _T_283 = _T_189 ? 4'h5 : _T_282; // @[Lookup.scala 33:37]
  wire [3:0] _T_284 = _T_187 ? 4'h4 : _T_283; // @[Lookup.scala 33:37]
  wire [3:0] _T_285 = _T_185 ? 4'h4 : _T_284; // @[Lookup.scala 33:37]
  wire [3:0] _T_286 = _T_183 ? 4'h5 : _T_285; // @[Lookup.scala 33:37]
  wire [3:0] _T_287 = _T_181 ? 4'h4 : _T_286; // @[Lookup.scala 33:37]
  wire [3:0] _T_288 = _T_179 ? 4'h4 : _T_287; // @[Lookup.scala 33:37]
  wire [3:0] _T_289 = _T_177 ? 4'h4 : _T_288; // @[Lookup.scala 33:37]
  wire [3:0] _T_290 = _T_175 ? 4'h4 : _T_289; // @[Lookup.scala 33:37]
  wire [3:0] _T_291 = _T_173 ? 4'h1 : _T_290; // @[Lookup.scala 33:37]
  wire [3:0] _T_292 = _T_171 ? 4'h1 : _T_291; // @[Lookup.scala 33:37]
  wire [3:0] _T_293 = _T_169 ? 4'h7 : _T_292; // @[Lookup.scala 33:37]
  wire [3:0] _T_294 = _T_167 ? 4'h5 : _T_293; // @[Lookup.scala 33:37]
  wire [3:0] _T_295 = _T_165 ? 4'h5 : _T_294; // @[Lookup.scala 33:37]
  wire [3:0] _T_296 = _T_163 ? 4'h5 : _T_295; // @[Lookup.scala 33:37]
  wire [3:0] _T_297 = _T_161 ? 4'h5 : _T_296; // @[Lookup.scala 33:37]
  wire [3:0] _T_298 = _T_159 ? 4'h5 : _T_297; // @[Lookup.scala 33:37]
  wire [3:0] _T_299 = _T_157 ? 4'h5 : _T_298; // @[Lookup.scala 33:37]
  wire [3:0] _T_300 = _T_155 ? 4'h4 : _T_299; // @[Lookup.scala 33:37]
  wire [3:0] _T_301 = _T_153 ? 4'h4 : _T_300; // @[Lookup.scala 33:37]
  wire [3:0] _T_302 = _T_151 ? 4'h4 : _T_301; // @[Lookup.scala 33:37]
  wire [3:0] _T_303 = _T_149 ? 4'h4 : _T_302; // @[Lookup.scala 33:37]
  wire [3:0] _T_304 = _T_147 ? 4'h4 : _T_303; // @[Lookup.scala 33:37]
  wire [3:0] _T_305 = _T_145 ? 4'h4 : _T_304; // @[Lookup.scala 33:37]
  wire [3:0] _T_306 = _T_143 ? 4'h4 : _T_305; // @[Lookup.scala 33:37]
  wire [3:0] _T_307 = _T_141 ? 4'h4 : _T_306; // @[Lookup.scala 33:37]
  wire [3:0] _T_308 = _T_139 ? 4'h4 : _T_307; // @[Lookup.scala 33:37]
  wire [3:0] _T_309 = _T_137 ? 4'h2 : _T_308; // @[Lookup.scala 33:37]
  wire [3:0] _T_310 = _T_135 ? 4'h2 : _T_309; // @[Lookup.scala 33:37]
  wire [3:0] _T_311 = _T_133 ? 4'h4 : _T_310; // @[Lookup.scala 33:37]
  wire [3:0] _T_312 = _T_131 ? 4'h4 : _T_311; // @[Lookup.scala 33:37]
  wire [3:0] _T_313 = _T_129 ? 4'h4 : _T_312; // @[Lookup.scala 33:37]
  wire [3:0] _T_314 = _T_127 ? 4'h0 : _T_313; // @[Lookup.scala 33:37]
  wire [3:0] _T_315 = _T_125 ? 4'h5 : _T_314; // @[Lookup.scala 33:37]
  wire [3:0] _T_316 = _T_123 ? 4'h5 : _T_315; // @[Lookup.scala 33:37]
  wire [3:0] _T_317 = _T_121 ? 4'h5 : _T_316; // @[Lookup.scala 33:37]
  wire [3:0] _T_318 = _T_119 ? 4'h5 : _T_317; // @[Lookup.scala 33:37]
  wire [3:0] _T_319 = _T_117 ? 4'h5 : _T_318; // @[Lookup.scala 33:37]
  wire [3:0] _T_320 = _T_115 ? 4'h5 : _T_319; // @[Lookup.scala 33:37]
  wire [3:0] _T_321 = _T_113 ? 4'h5 : _T_320; // @[Lookup.scala 33:37]
  wire [3:0] _T_322 = _T_111 ? 4'h5 : _T_321; // @[Lookup.scala 33:37]
  wire [3:0] _T_323 = _T_109 ? 4'h5 : _T_322; // @[Lookup.scala 33:37]
  wire [3:0] _T_324 = _T_107 ? 4'h5 : _T_323; // @[Lookup.scala 33:37]
  wire [3:0] _T_325 = _T_105 ? 4'h5 : _T_324; // @[Lookup.scala 33:37]
  wire [3:0] _T_326 = _T_103 ? 4'h5 : _T_325; // @[Lookup.scala 33:37]
  wire [3:0] _T_327 = _T_101 ? 4'h5 : _T_326; // @[Lookup.scala 33:37]
  wire [3:0] _T_328 = _T_99 ? 4'h4 : _T_327; // @[Lookup.scala 33:37]
  wire [3:0] _T_329 = _T_97 ? 4'h2 : _T_328; // @[Lookup.scala 33:37]
  wire [3:0] _T_330 = _T_95 ? 4'h4 : _T_329; // @[Lookup.scala 33:37]
  wire [3:0] _T_331 = _T_93 ? 4'h4 : _T_330; // @[Lookup.scala 33:37]
  wire [3:0] _T_332 = _T_91 ? 4'h5 : _T_331; // @[Lookup.scala 33:37]
  wire [3:0] _T_333 = _T_89 ? 4'h5 : _T_332; // @[Lookup.scala 33:37]
  wire [3:0] _T_334 = _T_87 ? 4'h5 : _T_333; // @[Lookup.scala 33:37]
  wire [3:0] _T_335 = _T_85 ? 4'h5 : _T_334; // @[Lookup.scala 33:37]
  wire [3:0] _T_336 = _T_83 ? 4'h5 : _T_335; // @[Lookup.scala 33:37]
  wire [3:0] _T_337 = _T_81 ? 4'h4 : _T_336; // @[Lookup.scala 33:37]
  wire [3:0] _T_338 = _T_79 ? 4'h4 : _T_337; // @[Lookup.scala 33:37]
  wire [3:0] _T_339 = _T_77 ? 4'h4 : _T_338; // @[Lookup.scala 33:37]
  wire [3:0] _T_340 = _T_75 ? 4'h4 : _T_339; // @[Lookup.scala 33:37]
  wire [3:0] _T_341 = _T_73 ? 4'h2 : _T_340; // @[Lookup.scala 33:37]
  wire [3:0] _T_342 = _T_71 ? 4'h2 : _T_341; // @[Lookup.scala 33:37]
  wire [3:0] _T_343 = _T_69 ? 4'h2 : _T_342; // @[Lookup.scala 33:37]
  wire [3:0] _T_344 = _T_67 ? 4'h4 : _T_343; // @[Lookup.scala 33:37]
  wire [3:0] _T_345 = _T_65 ? 4'h4 : _T_344; // @[Lookup.scala 33:37]
  wire [3:0] _T_346 = _T_63 ? 4'h4 : _T_345; // @[Lookup.scala 33:37]
  wire [3:0] _T_347 = _T_61 ? 4'h4 : _T_346; // @[Lookup.scala 33:37]
  wire [3:0] _T_348 = _T_59 ? 4'h4 : _T_347; // @[Lookup.scala 33:37]
  wire [3:0] _T_349 = _T_57 ? 4'h1 : _T_348; // @[Lookup.scala 33:37]
  wire [3:0] _T_350 = _T_55 ? 4'h1 : _T_349; // @[Lookup.scala 33:37]
  wire [3:0] _T_351 = _T_53 ? 4'h1 : _T_350; // @[Lookup.scala 33:37]
  wire [3:0] _T_352 = _T_51 ? 4'h1 : _T_351; // @[Lookup.scala 33:37]
  wire [3:0] _T_353 = _T_49 ? 4'h1 : _T_352; // @[Lookup.scala 33:37]
  wire [3:0] _T_354 = _T_47 ? 4'h1 : _T_353; // @[Lookup.scala 33:37]
  wire [3:0] _T_355 = _T_45 ? 4'h4 : _T_354; // @[Lookup.scala 33:37]
  wire [3:0] _T_356 = _T_43 ? 4'h7 : _T_355; // @[Lookup.scala 33:37]
  wire [3:0] _T_357 = _T_41 ? 4'h6 : _T_356; // @[Lookup.scala 33:37]
  wire [3:0] _T_358 = _T_39 ? 4'h6 : _T_357; // @[Lookup.scala 33:37]
  wire [3:0] _T_359 = _T_37 ? 4'h5 : _T_358; // @[Lookup.scala 33:37]
  wire [3:0] _T_360 = _T_35 ? 4'h5 : _T_359; // @[Lookup.scala 33:37]
  wire [3:0] _T_361 = _T_33 ? 4'h5 : _T_360; // @[Lookup.scala 33:37]
  wire [3:0] _T_362 = _T_31 ? 4'h5 : _T_361; // @[Lookup.scala 33:37]
  wire [3:0] _T_363 = _T_29 ? 4'h5 : _T_362; // @[Lookup.scala 33:37]
  wire [3:0] _T_364 = _T_27 ? 4'h5 : _T_363; // @[Lookup.scala 33:37]
  wire [3:0] _T_365 = _T_25 ? 4'h5 : _T_364; // @[Lookup.scala 33:37]
  wire [3:0] _T_366 = _T_23 ? 4'h5 : _T_365; // @[Lookup.scala 33:37]
  wire [3:0] _T_367 = _T_21 ? 4'h5 : _T_366; // @[Lookup.scala 33:37]
  wire [3:0] _T_368 = _T_19 ? 4'h5 : _T_367; // @[Lookup.scala 33:37]
  wire [3:0] _T_369 = _T_17 ? 4'h4 : _T_368; // @[Lookup.scala 33:37]
  wire [3:0] _T_370 = _T_15 ? 4'h4 : _T_369; // @[Lookup.scala 33:37]
  wire [3:0] _T_371 = _T_13 ? 4'h4 : _T_370; // @[Lookup.scala 33:37]
  wire [3:0] _T_372 = _T_11 ? 4'h4 : _T_371; // @[Lookup.scala 33:37]
  wire [3:0] _T_373 = _T_9 ? 4'h4 : _T_372; // @[Lookup.scala 33:37]
  wire [3:0] _T_374 = _T_7 ? 4'h4 : _T_373; // @[Lookup.scala 33:37]
  wire [3:0] _T_375 = _T_5 ? 4'h4 : _T_374; // @[Lookup.scala 33:37]
  wire [3:0] _T_376 = _T_3 ? 4'h4 : _T_375; // @[Lookup.scala 33:37]
  wire [3:0] decodeList_0 = _T_1 ? 4'h4 : _T_376; // @[Lookup.scala 33:37]
  wire [1:0] _T_377 = _T_251 ? 2'h0 : 2'h3; // @[Lookup.scala 33:37]
  wire [2:0] _T_378 = _T_249 ? 3'h4 : {{1'd0}, _T_377}; // @[Lookup.scala 33:37]
  wire [2:0] _T_379 = _T_247 ? 3'h3 : _T_378; // @[Lookup.scala 33:37]
  wire [2:0] _T_380 = _T_245 ? 3'h3 : _T_379; // @[Lookup.scala 33:37]
  wire [2:0] _T_381 = _T_243 ? 3'h3 : _T_380; // @[Lookup.scala 33:37]
  wire [2:0] _T_382 = _T_241 ? 3'h3 : _T_381; // @[Lookup.scala 33:37]
  wire [2:0] _T_383 = _T_239 ? 3'h3 : _T_382; // @[Lookup.scala 33:37]
  wire [2:0] _T_384 = _T_237 ? 3'h3 : _T_383; // @[Lookup.scala 33:37]
  wire [2:0] _T_385 = _T_235 ? 3'h1 : _T_384; // @[Lookup.scala 33:37]
  wire [2:0] _T_386 = _T_233 ? 3'h1 : _T_385; // @[Lookup.scala 33:37]
  wire [2:0] _T_387 = _T_231 ? 3'h1 : _T_386; // @[Lookup.scala 33:37]
  wire [2:0] _T_388 = _T_229 ? 3'h1 : _T_387; // @[Lookup.scala 33:37]
  wire [2:0] _T_389 = _T_227 ? 3'h1 : _T_388; // @[Lookup.scala 33:37]
  wire [2:0] _T_390 = _T_225 ? 3'h1 : _T_389; // @[Lookup.scala 33:37]
  wire [2:0] _T_391 = _T_223 ? 3'h1 : _T_390; // @[Lookup.scala 33:37]
  wire [2:0] _T_392 = _T_221 ? 3'h1 : _T_391; // @[Lookup.scala 33:37]
  wire [2:0] _T_393 = _T_219 ? 3'h1 : _T_392; // @[Lookup.scala 33:37]
  wire [2:0] _T_394 = _T_217 ? 3'h1 : _T_393; // @[Lookup.scala 33:37]
  wire [2:0] _T_395 = _T_215 ? 3'h1 : _T_394; // @[Lookup.scala 33:37]
  wire [2:0] _T_396 = _T_213 ? 3'h1 : _T_395; // @[Lookup.scala 33:37]
  wire [2:0] _T_397 = _T_211 ? 3'h1 : _T_396; // @[Lookup.scala 33:37]
  wire [2:0] _T_398 = _T_209 ? 3'h3 : _T_397; // @[Lookup.scala 33:37]
  wire [2:0] _T_399 = _T_207 ? 3'h4 : _T_398; // @[Lookup.scala 33:37]
  wire [2:0] _T_400 = _T_205 ? 3'h3 : _T_399; // @[Lookup.scala 33:37]
  wire [2:0] _T_401 = _T_203 ? 3'h0 : _T_400; // @[Lookup.scala 33:37]
  wire [2:0] _T_402 = _T_201 ? 3'h4 : _T_401; // @[Lookup.scala 33:37]
  wire [2:0] _T_403 = _T_199 ? 3'h3 : _T_402; // @[Lookup.scala 33:37]
  wire [2:0] _T_404 = _T_197 ? 3'h3 : _T_403; // @[Lookup.scala 33:37]
  wire [2:0] _T_405 = _T_195 ? 3'h3 : _T_404; // @[Lookup.scala 33:37]
  wire [2:0] _T_406 = _T_193 ? 3'h1 : _T_405; // @[Lookup.scala 33:37]
  wire [2:0] _T_407 = _T_191 ? 3'h1 : _T_406; // @[Lookup.scala 33:37]
  wire [2:0] _T_408 = _T_189 ? 3'h0 : _T_407; // @[Lookup.scala 33:37]
  wire [2:0] _T_409 = _T_187 ? 3'h0 : _T_408; // @[Lookup.scala 33:37]
  wire [2:0] _T_410 = _T_185 ? 3'h3 : _T_409; // @[Lookup.scala 33:37]
  wire [2:0] _T_411 = _T_183 ? 3'h0 : _T_410; // @[Lookup.scala 33:37]
  wire [2:0] _T_412 = _T_181 ? 3'h0 : _T_411; // @[Lookup.scala 33:37]
  wire [2:0] _T_413 = _T_179 ? 3'h1 : _T_412; // @[Lookup.scala 33:37]
  wire [2:0] _T_414 = _T_177 ? 3'h1 : _T_413; // @[Lookup.scala 33:37]
  wire [2:0] _T_415 = _T_175 ? 3'h0 : _T_414; // @[Lookup.scala 33:37]
  wire [2:0] _T_416 = _T_173 ? 3'h0 : _T_415; // @[Lookup.scala 33:37]
  wire [2:0] _T_417 = _T_171 ? 3'h0 : _T_416; // @[Lookup.scala 33:37]
  wire [2:0] _T_418 = _T_169 ? 3'h0 : _T_417; // @[Lookup.scala 33:37]
  wire [2:0] _T_419 = _T_167 ? 3'h0 : _T_418; // @[Lookup.scala 33:37]
  wire [2:0] _T_420 = _T_165 ? 3'h0 : _T_419; // @[Lookup.scala 33:37]
  wire [2:0] _T_421 = _T_163 ? 3'h0 : _T_420; // @[Lookup.scala 33:37]
  wire [2:0] _T_422 = _T_161 ? 3'h0 : _T_421; // @[Lookup.scala 33:37]
  wire [2:0] _T_423 = _T_159 ? 3'h0 : _T_422; // @[Lookup.scala 33:37]
  wire [2:0] _T_424 = _T_157 ? 3'h0 : _T_423; // @[Lookup.scala 33:37]
  wire [2:0] _T_425 = _T_155 ? 3'h0 : _T_424; // @[Lookup.scala 33:37]
  wire [2:0] _T_426 = _T_153 ? 3'h0 : _T_425; // @[Lookup.scala 33:37]
  wire [2:0] _T_427 = _T_151 ? 3'h0 : _T_426; // @[Lookup.scala 33:37]
  wire [2:0] _T_428 = _T_149 ? 3'h0 : _T_427; // @[Lookup.scala 33:37]
  wire [2:0] _T_429 = _T_147 ? 3'h0 : _T_428; // @[Lookup.scala 33:37]
  wire [2:0] _T_430 = _T_145 ? 3'h0 : _T_429; // @[Lookup.scala 33:37]
  wire [2:0] _T_431 = _T_143 ? 3'h0 : _T_430; // @[Lookup.scala 33:37]
  wire [2:0] _T_432 = _T_141 ? 3'h0 : _T_431; // @[Lookup.scala 33:37]
  wire [2:0] _T_433 = _T_139 ? 3'h0 : _T_432; // @[Lookup.scala 33:37]
  wire [2:0] _T_434 = _T_137 ? 3'h1 : _T_433; // @[Lookup.scala 33:37]
  wire [2:0] _T_435 = _T_135 ? 3'h1 : _T_434; // @[Lookup.scala 33:37]
  wire [2:0] _T_436 = _T_133 ? 3'h1 : _T_435; // @[Lookup.scala 33:37]
  wire [2:0] _T_437 = _T_131 ? 3'h1 : _T_436; // @[Lookup.scala 33:37]
  wire [2:0] _T_438 = _T_129 ? 3'h0 : _T_437; // @[Lookup.scala 33:37]
  wire [2:0] _T_439 = _T_127 ? 3'h3 : _T_438; // @[Lookup.scala 33:37]
  wire [2:0] _T_440 = _T_125 ? 3'h2 : _T_439; // @[Lookup.scala 33:37]
  wire [2:0] _T_441 = _T_123 ? 3'h2 : _T_440; // @[Lookup.scala 33:37]
  wire [2:0] _T_442 = _T_121 ? 3'h2 : _T_441; // @[Lookup.scala 33:37]
  wire [2:0] _T_443 = _T_119 ? 3'h2 : _T_442; // @[Lookup.scala 33:37]
  wire [2:0] _T_444 = _T_117 ? 3'h2 : _T_443; // @[Lookup.scala 33:37]
  wire [2:0] _T_445 = _T_115 ? 3'h2 : _T_444; // @[Lookup.scala 33:37]
  wire [2:0] _T_446 = _T_113 ? 3'h2 : _T_445; // @[Lookup.scala 33:37]
  wire [2:0] _T_447 = _T_111 ? 3'h2 : _T_446; // @[Lookup.scala 33:37]
  wire [2:0] _T_448 = _T_109 ? 3'h2 : _T_447; // @[Lookup.scala 33:37]
  wire [2:0] _T_449 = _T_107 ? 3'h2 : _T_448; // @[Lookup.scala 33:37]
  wire [2:0] _T_450 = _T_105 ? 3'h2 : _T_449; // @[Lookup.scala 33:37]
  wire [2:0] _T_451 = _T_103 ? 3'h2 : _T_450; // @[Lookup.scala 33:37]
  wire [2:0] _T_452 = _T_101 ? 3'h2 : _T_451; // @[Lookup.scala 33:37]
  wire [2:0] _T_453 = _T_99 ? 3'h3 : _T_452; // @[Lookup.scala 33:37]
  wire [2:0] _T_454 = _T_97 ? 3'h1 : _T_453; // @[Lookup.scala 33:37]
  wire [2:0] _T_455 = _T_95 ? 3'h1 : _T_454; // @[Lookup.scala 33:37]
  wire [2:0] _T_456 = _T_93 ? 3'h1 : _T_455; // @[Lookup.scala 33:37]
  wire [2:0] _T_457 = _T_91 ? 3'h0 : _T_456; // @[Lookup.scala 33:37]
  wire [2:0] _T_458 = _T_89 ? 3'h0 : _T_457; // @[Lookup.scala 33:37]
  wire [2:0] _T_459 = _T_87 ? 3'h0 : _T_458; // @[Lookup.scala 33:37]
  wire [2:0] _T_460 = _T_85 ? 3'h0 : _T_459; // @[Lookup.scala 33:37]
  wire [2:0] _T_461 = _T_83 ? 3'h0 : _T_460; // @[Lookup.scala 33:37]
  wire [2:0] _T_462 = _T_81 ? 3'h0 : _T_461; // @[Lookup.scala 33:37]
  wire [2:0] _T_463 = _T_79 ? 3'h0 : _T_462; // @[Lookup.scala 33:37]
  wire [2:0] _T_464 = _T_77 ? 3'h0 : _T_463; // @[Lookup.scala 33:37]
  wire [2:0] _T_465 = _T_75 ? 3'h0 : _T_464; // @[Lookup.scala 33:37]
  wire [2:0] _T_466 = _T_73 ? 3'h1 : _T_465; // @[Lookup.scala 33:37]
  wire [2:0] _T_467 = _T_71 ? 3'h1 : _T_466; // @[Lookup.scala 33:37]
  wire [2:0] _T_468 = _T_69 ? 3'h1 : _T_467; // @[Lookup.scala 33:37]
  wire [2:0] _T_469 = _T_67 ? 3'h1 : _T_468; // @[Lookup.scala 33:37]
  wire [2:0] _T_470 = _T_65 ? 3'h1 : _T_469; // @[Lookup.scala 33:37]
  wire [2:0] _T_471 = _T_63 ? 3'h1 : _T_470; // @[Lookup.scala 33:37]
  wire [2:0] _T_472 = _T_61 ? 3'h1 : _T_471; // @[Lookup.scala 33:37]
  wire [2:0] _T_473 = _T_59 ? 3'h1 : _T_472; // @[Lookup.scala 33:37]
  wire [2:0] _T_474 = _T_57 ? 3'h0 : _T_473; // @[Lookup.scala 33:37]
  wire [2:0] _T_475 = _T_55 ? 3'h0 : _T_474; // @[Lookup.scala 33:37]
  wire [2:0] _T_476 = _T_53 ? 3'h0 : _T_475; // @[Lookup.scala 33:37]
  wire [2:0] _T_477 = _T_51 ? 3'h0 : _T_476; // @[Lookup.scala 33:37]
  wire [2:0] _T_478 = _T_49 ? 3'h0 : _T_477; // @[Lookup.scala 33:37]
  wire [2:0] _T_479 = _T_47 ? 3'h0 : _T_478; // @[Lookup.scala 33:37]
  wire [2:0] _T_480 = _T_45 ? 3'h0 : _T_479; // @[Lookup.scala 33:37]
  wire [2:0] _T_481 = _T_43 ? 3'h0 : _T_480; // @[Lookup.scala 33:37]
  wire [2:0] _T_482 = _T_41 ? 3'h0 : _T_481; // @[Lookup.scala 33:37]
  wire [2:0] _T_483 = _T_39 ? 3'h0 : _T_482; // @[Lookup.scala 33:37]
  wire [2:0] _T_484 = _T_37 ? 3'h0 : _T_483; // @[Lookup.scala 33:37]
  wire [2:0] _T_485 = _T_35 ? 3'h0 : _T_484; // @[Lookup.scala 33:37]
  wire [2:0] _T_486 = _T_33 ? 3'h0 : _T_485; // @[Lookup.scala 33:37]
  wire [2:0] _T_487 = _T_31 ? 3'h0 : _T_486; // @[Lookup.scala 33:37]
  wire [2:0] _T_488 = _T_29 ? 3'h0 : _T_487; // @[Lookup.scala 33:37]
  wire [2:0] _T_489 = _T_27 ? 3'h0 : _T_488; // @[Lookup.scala 33:37]
  wire [2:0] _T_490 = _T_25 ? 3'h0 : _T_489; // @[Lookup.scala 33:37]
  wire [2:0] _T_491 = _T_23 ? 3'h0 : _T_490; // @[Lookup.scala 33:37]
  wire [2:0] _T_492 = _T_21 ? 3'h0 : _T_491; // @[Lookup.scala 33:37]
  wire [2:0] _T_493 = _T_19 ? 3'h0 : _T_492; // @[Lookup.scala 33:37]
  wire [2:0] _T_494 = _T_17 ? 3'h0 : _T_493; // @[Lookup.scala 33:37]
  wire [2:0] _T_495 = _T_15 ? 3'h0 : _T_494; // @[Lookup.scala 33:37]
  wire [2:0] _T_496 = _T_13 ? 3'h0 : _T_495; // @[Lookup.scala 33:37]
  wire [2:0] _T_497 = _T_11 ? 3'h0 : _T_496; // @[Lookup.scala 33:37]
  wire [2:0] _T_498 = _T_9 ? 3'h0 : _T_497; // @[Lookup.scala 33:37]
  wire [2:0] _T_499 = _T_7 ? 3'h0 : _T_498; // @[Lookup.scala 33:37]
  wire [2:0] _T_500 = _T_5 ? 3'h0 : _T_499; // @[Lookup.scala 33:37]
  wire [2:0] _T_501 = _T_3 ? 3'h0 : _T_500; // @[Lookup.scala 33:37]
  wire [2:0] decodeList_1 = _T_1 ? 3'h0 : _T_501; // @[Lookup.scala 33:37]
  wire [6:0] _T_502 = _T_251 ? 7'h7e : 7'h0; // @[Lookup.scala 33:37]
  wire [6:0] _T_503 = _T_249 ? 7'h1 : _T_502; // @[Lookup.scala 33:37]
  wire [6:0] _T_504 = _T_247 ? 7'h7 : _T_503; // @[Lookup.scala 33:37]
  wire [6:0] _T_505 = _T_245 ? 7'h6 : _T_504; // @[Lookup.scala 33:37]
  wire [6:0] _T_506 = _T_243 ? 7'h5 : _T_505; // @[Lookup.scala 33:37]
  wire [6:0] _T_507 = _T_241 ? 7'h3 : _T_506; // @[Lookup.scala 33:37]
  wire [6:0] _T_508 = _T_239 ? 7'h2 : _T_507; // @[Lookup.scala 33:37]
  wire [6:0] _T_509 = _T_237 ? 7'h1 : _T_508; // @[Lookup.scala 33:37]
  wire [6:0] _T_510 = _T_235 ? 7'h32 : _T_509; // @[Lookup.scala 33:37]
  wire [6:0] _T_511 = _T_233 ? 7'h31 : _T_510; // @[Lookup.scala 33:37]
  wire [6:0] _T_512 = _T_231 ? 7'h30 : _T_511; // @[Lookup.scala 33:37]
  wire [6:0] _T_513 = _T_229 ? 7'h37 : _T_512; // @[Lookup.scala 33:37]
  wire [6:0] _T_514 = _T_227 ? 7'h26 : _T_513; // @[Lookup.scala 33:37]
  wire [6:0] _T_515 = _T_225 ? 7'h25 : _T_514; // @[Lookup.scala 33:37]
  wire [6:0] _T_516 = _T_223 ? 7'h24 : _T_515; // @[Lookup.scala 33:37]
  wire [6:0] _T_517 = _T_221 ? 7'h63 : _T_516; // @[Lookup.scala 33:37]
  wire [6:0] _T_518 = _T_219 ? 7'h22 : _T_517; // @[Lookup.scala 33:37]
  wire [6:0] _T_519 = _T_217 ? 7'h21 : _T_518; // @[Lookup.scala 33:37]
  wire [6:0] _T_520 = _T_215 ? 7'h21 : _T_519; // @[Lookup.scala 33:37]
  wire [6:0] _T_521 = _T_213 ? 7'h20 : _T_520; // @[Lookup.scala 33:37]
  wire [6:0] _T_522 = _T_211 ? 7'h20 : _T_521; // @[Lookup.scala 33:37]
  wire [6:0] _T_523 = _T_209 ? 7'h0 : _T_522; // @[Lookup.scala 33:37]
  wire [6:0] _T_524 = _T_207 ? 7'h2 : _T_523; // @[Lookup.scala 33:37]
  wire [6:0] _T_525 = _T_205 ? 7'h0 : _T_524; // @[Lookup.scala 33:37]
  wire [6:0] _T_526 = _T_203 ? 7'h40 : _T_525; // @[Lookup.scala 33:37]
  wire [6:0] _T_527 = _T_201 ? 7'h0 : _T_526; // @[Lookup.scala 33:37]
  wire [6:0] _T_528 = _T_199 ? 7'h0 : _T_527; // @[Lookup.scala 33:37]
  wire [6:0] _T_529 = _T_197 ? 7'h0 : _T_528; // @[Lookup.scala 33:37]
  wire [6:0] _T_530 = _T_195 ? 7'h0 : _T_529; // @[Lookup.scala 33:37]
  wire [6:0] _T_531 = _T_193 ? 7'hb : _T_530; // @[Lookup.scala 33:37]
  wire [6:0] _T_532 = _T_191 ? 7'ha : _T_531; // @[Lookup.scala 33:37]
  wire [6:0] _T_533 = _T_189 ? 7'h40 : _T_532; // @[Lookup.scala 33:37]
  wire [6:0] _T_534 = _T_187 ? 7'h5a : _T_533; // @[Lookup.scala 33:37]
  wire [6:0] _T_535 = _T_185 ? 7'h0 : _T_534; // @[Lookup.scala 33:37]
  wire [6:0] _T_536 = _T_183 ? 7'h40 : _T_535; // @[Lookup.scala 33:37]
  wire [6:0] _T_537 = _T_181 ? 7'h5a : _T_536; // @[Lookup.scala 33:37]
  wire [6:0] _T_538 = _T_179 ? 7'h3 : _T_537; // @[Lookup.scala 33:37]
  wire [6:0] _T_539 = _T_177 ? 7'h2 : _T_538; // @[Lookup.scala 33:37]
  wire [6:0] _T_540 = _T_175 ? 7'h1 : _T_539; // @[Lookup.scala 33:37]
  wire [6:0] _T_541 = _T_173 ? 7'h11 : _T_540; // @[Lookup.scala 33:37]
  wire [6:0] _T_542 = _T_171 ? 7'h10 : _T_541; // @[Lookup.scala 33:37]
  wire [6:0] _T_543 = _T_169 ? 7'h58 : _T_542; // @[Lookup.scala 33:37]
  wire [6:0] _T_544 = _T_167 ? 7'h60 : _T_543; // @[Lookup.scala 33:37]
  wire [6:0] _T_545 = _T_165 ? 7'h28 : _T_544; // @[Lookup.scala 33:37]
  wire [6:0] _T_546 = _T_163 ? 7'h7 : _T_545; // @[Lookup.scala 33:37]
  wire [6:0] _T_547 = _T_161 ? 7'h6 : _T_546; // @[Lookup.scala 33:37]
  wire [6:0] _T_548 = _T_159 ? 7'h4 : _T_547; // @[Lookup.scala 33:37]
  wire [6:0] _T_549 = _T_157 ? 7'h8 : _T_548; // @[Lookup.scala 33:37]
  wire [6:0] _T_550 = _T_155 ? 7'h7 : _T_549; // @[Lookup.scala 33:37]
  wire [6:0] _T_551 = _T_153 ? 7'hd : _T_550; // @[Lookup.scala 33:37]
  wire [6:0] _T_552 = _T_151 ? 7'h5 : _T_551; // @[Lookup.scala 33:37]
  wire [6:0] _T_553 = _T_149 ? 7'h40 : _T_552; // @[Lookup.scala 33:37]
  wire [6:0] _T_554 = _T_147 ? 7'h40 : _T_553; // @[Lookup.scala 33:37]
  wire [6:0] _T_555 = _T_145 ? 7'h40 : _T_554; // @[Lookup.scala 33:37]
  wire [6:0] _T_556 = _T_143 ? 7'h60 : _T_555; // @[Lookup.scala 33:37]
  wire [6:0] _T_557 = _T_141 ? 7'h40 : _T_556; // @[Lookup.scala 33:37]
  wire [6:0] _T_558 = _T_139 ? 7'h40 : _T_557; // @[Lookup.scala 33:37]
  wire [6:0] _T_559 = _T_137 ? 7'hb : _T_558; // @[Lookup.scala 33:37]
  wire [6:0] _T_560 = _T_135 ? 7'ha : _T_559; // @[Lookup.scala 33:37]
  wire [6:0] _T_561 = _T_133 ? 7'h3 : _T_560; // @[Lookup.scala 33:37]
  wire [6:0] _T_562 = _T_131 ? 7'h2 : _T_561; // @[Lookup.scala 33:37]
  wire [6:0] _T_563 = _T_129 ? 7'h40 : _T_562; // @[Lookup.scala 33:37]
  wire [6:0] _T_564 = _T_127 ? 7'h0 : _T_563; // @[Lookup.scala 33:37]
  wire [6:0] _T_565 = _T_125 ? 7'hf : _T_564; // @[Lookup.scala 33:37]
  wire [6:0] _T_566 = _T_123 ? 7'he : _T_565; // @[Lookup.scala 33:37]
  wire [6:0] _T_567 = _T_121 ? 7'hd : _T_566; // @[Lookup.scala 33:37]
  wire [6:0] _T_568 = _T_119 ? 7'hc : _T_567; // @[Lookup.scala 33:37]
  wire [6:0] _T_569 = _T_117 ? 7'h8 : _T_568; // @[Lookup.scala 33:37]
  wire [6:0] _T_570 = _T_115 ? 7'h7 : _T_569; // @[Lookup.scala 33:37]
  wire [6:0] _T_571 = _T_113 ? 7'h6 : _T_570; // @[Lookup.scala 33:37]
  wire [6:0] _T_572 = _T_111 ? 7'h5 : _T_571; // @[Lookup.scala 33:37]
  wire [6:0] _T_573 = _T_109 ? 7'h4 : _T_572; // @[Lookup.scala 33:37]
  wire [6:0] _T_574 = _T_107 ? 7'h3 : _T_573; // @[Lookup.scala 33:37]
  wire [6:0] _T_575 = _T_105 ? 7'h2 : _T_574; // @[Lookup.scala 33:37]
  wire [6:0] _T_576 = _T_103 ? 7'h1 : _T_575; // @[Lookup.scala 33:37]
  wire [6:0] _T_577 = _T_101 ? 7'h0 : _T_576; // @[Lookup.scala 33:37]
  wire [6:0] _T_578 = _T_99 ? 7'h2 : _T_577; // @[Lookup.scala 33:37]
  wire [6:0] _T_579 = _T_97 ? 7'hb : _T_578; // @[Lookup.scala 33:37]
  wire [6:0] _T_580 = _T_95 ? 7'h3 : _T_579; // @[Lookup.scala 33:37]
  wire [6:0] _T_581 = _T_93 ? 7'h6 : _T_580; // @[Lookup.scala 33:37]
  wire [6:0] _T_582 = _T_91 ? 7'h28 : _T_581; // @[Lookup.scala 33:37]
  wire [6:0] _T_583 = _T_89 ? 7'h60 : _T_582; // @[Lookup.scala 33:37]
  wire [6:0] _T_584 = _T_87 ? 7'h2d : _T_583; // @[Lookup.scala 33:37]
  wire [6:0] _T_585 = _T_85 ? 7'h25 : _T_584; // @[Lookup.scala 33:37]
  wire [6:0] _T_586 = _T_83 ? 7'h21 : _T_585; // @[Lookup.scala 33:37]
  wire [6:0] _T_587 = _T_81 ? 7'h2d : _T_586; // @[Lookup.scala 33:37]
  wire [6:0] _T_588 = _T_79 ? 7'h25 : _T_587; // @[Lookup.scala 33:37]
  wire [6:0] _T_589 = _T_77 ? 7'h21 : _T_588; // @[Lookup.scala 33:37]
  wire [6:0] _T_590 = _T_75 ? 7'h60 : _T_589; // @[Lookup.scala 33:37]
  wire [6:0] _T_591 = _T_73 ? 7'ha : _T_590; // @[Lookup.scala 33:37]
  wire [6:0] _T_592 = _T_71 ? 7'h9 : _T_591; // @[Lookup.scala 33:37]
  wire [6:0] _T_593 = _T_69 ? 7'h8 : _T_592; // @[Lookup.scala 33:37]
  wire [6:0] _T_594 = _T_67 ? 7'h5 : _T_593; // @[Lookup.scala 33:37]
  wire [6:0] _T_595 = _T_65 ? 7'h4 : _T_594; // @[Lookup.scala 33:37]
  wire [6:0] _T_596 = _T_63 ? 7'h2 : _T_595; // @[Lookup.scala 33:37]
  wire [6:0] _T_597 = _T_61 ? 7'h1 : _T_596; // @[Lookup.scala 33:37]
  wire [6:0] _T_598 = _T_59 ? 7'h0 : _T_597; // @[Lookup.scala 33:37]
  wire [6:0] _T_599 = _T_57 ? 7'h17 : _T_598; // @[Lookup.scala 33:37]
  wire [6:0] _T_600 = _T_55 ? 7'h16 : _T_599; // @[Lookup.scala 33:37]
  wire [6:0] _T_601 = _T_53 ? 7'h15 : _T_600; // @[Lookup.scala 33:37]
  wire [6:0] _T_602 = _T_51 ? 7'h14 : _T_601; // @[Lookup.scala 33:37]
  wire [6:0] _T_603 = _T_49 ? 7'h11 : _T_602; // @[Lookup.scala 33:37]
  wire [6:0] _T_604 = _T_47 ? 7'h10 : _T_603; // @[Lookup.scala 33:37]
  wire [6:0] _T_605 = _T_45 ? 7'h5a : _T_604; // @[Lookup.scala 33:37]
  wire [6:0] _T_606 = _T_43 ? 7'h58 : _T_605; // @[Lookup.scala 33:37]
  wire [6:0] _T_607 = _T_41 ? 7'h40 : _T_606; // @[Lookup.scala 33:37]
  wire [6:0] _T_608 = _T_39 ? 7'h40 : _T_607; // @[Lookup.scala 33:37]
  wire [6:0] _T_609 = _T_37 ? 7'hd : _T_608; // @[Lookup.scala 33:37]
  wire [6:0] _T_610 = _T_35 ? 7'h8 : _T_609; // @[Lookup.scala 33:37]
  wire [6:0] _T_611 = _T_33 ? 7'h7 : _T_610; // @[Lookup.scala 33:37]
  wire [6:0] _T_612 = _T_31 ? 7'h6 : _T_611; // @[Lookup.scala 33:37]
  wire [6:0] _T_613 = _T_29 ? 7'h5 : _T_612; // @[Lookup.scala 33:37]
  wire [6:0] _T_614 = _T_27 ? 7'h4 : _T_613; // @[Lookup.scala 33:37]
  wire [6:0] _T_615 = _T_25 ? 7'h3 : _T_614; // @[Lookup.scala 33:37]
  wire [6:0] _T_616 = _T_23 ? 7'h2 : _T_615; // @[Lookup.scala 33:37]
  wire [6:0] _T_617 = _T_21 ? 7'h1 : _T_616; // @[Lookup.scala 33:37]
  wire [6:0] _T_618 = _T_19 ? 7'h40 : _T_617; // @[Lookup.scala 33:37]
  wire [6:0] _T_619 = _T_17 ? 7'hd : _T_618; // @[Lookup.scala 33:37]
  wire [6:0] _T_620 = _T_15 ? 7'h7 : _T_619; // @[Lookup.scala 33:37]
  wire [6:0] _T_621 = _T_13 ? 7'h6 : _T_620; // @[Lookup.scala 33:37]
  wire [6:0] _T_622 = _T_11 ? 7'h5 : _T_621; // @[Lookup.scala 33:37]
  wire [6:0] _T_623 = _T_9 ? 7'h4 : _T_622; // @[Lookup.scala 33:37]
  wire [6:0] _T_624 = _T_7 ? 7'h3 : _T_623; // @[Lookup.scala 33:37]
  wire [6:0] _T_625 = _T_5 ? 7'h2 : _T_624; // @[Lookup.scala 33:37]
  wire [6:0] _T_626 = _T_3 ? 7'h1 : _T_625; // @[Lookup.scala 33:37]
  wire [6:0] decodeList_2 = _T_1 ? 7'h40 : _T_626; // @[Lookup.scala 33:37]
  wire  hasIntr = |intrVecIDU; // @[IDU.scala 170:22]
  wire [3:0] instrType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 4'h0 : decodeList_0; // @[IDU.scala 36:75]
  wire [2:0] fuType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 3'h3 : decodeList_1; // @[IDU.scala 36:75]
  wire [6:0] fuOpType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 7'h0 : decodeList_2; // @[IDU.scala 36:75]
  wire  isRVC = io_in_bits_instr[1:0] != 2'h3; // @[IDU.scala 38:45]
  wire [4:0] _T_700 = _T_193 ? 5'h3 : 5'h10; // @[Lookup.scala 33:37]
  wire [4:0] _T_701 = _T_191 ? 5'h2 : _T_700; // @[Lookup.scala 33:37]
  wire [4:0] _T_702 = _T_189 ? 5'h10 : _T_701; // @[Lookup.scala 33:37]
  wire [4:0] _T_703 = _T_187 ? 5'h10 : _T_702; // @[Lookup.scala 33:37]
  wire [4:0] _T_704 = _T_185 ? 5'hf : _T_703; // @[Lookup.scala 33:37]
  wire [4:0] _T_705 = _T_183 ? 5'h10 : _T_704; // @[Lookup.scala 33:37]
  wire [4:0] _T_706 = _T_181 ? 5'h10 : _T_705; // @[Lookup.scala 33:37]
  wire [4:0] _T_707 = _T_179 ? 5'h1 : _T_706; // @[Lookup.scala 33:37]
  wire [4:0] _T_708 = _T_177 ? 5'h0 : _T_707; // @[Lookup.scala 33:37]
  wire [4:0] _T_709 = _T_175 ? 5'ha : _T_708; // @[Lookup.scala 33:37]
  wire [4:0] _T_710 = _T_173 ? 5'h9 : _T_709; // @[Lookup.scala 33:37]
  wire [4:0] _T_711 = _T_171 ? 5'h9 : _T_710; // @[Lookup.scala 33:37]
  wire [4:0] _T_712 = _T_169 ? 5'h8 : _T_711; // @[Lookup.scala 33:37]
  wire [4:0] _T_713 = _T_167 ? 5'h10 : _T_712; // @[Lookup.scala 33:37]
  wire [4:0] _T_714 = _T_165 ? 5'h10 : _T_713; // @[Lookup.scala 33:37]
  wire [4:0] _T_715 = _T_163 ? 5'h10 : _T_714; // @[Lookup.scala 33:37]
  wire [4:0] _T_716 = _T_161 ? 5'h10 : _T_715; // @[Lookup.scala 33:37]
  wire [4:0] _T_717 = _T_159 ? 5'h10 : _T_716; // @[Lookup.scala 33:37]
  wire [4:0] _T_718 = _T_157 ? 5'h10 : _T_717; // @[Lookup.scala 33:37]
  wire [4:0] _T_719 = _T_155 ? 5'ha : _T_718; // @[Lookup.scala 33:37]
  wire [4:0] _T_720 = _T_153 ? 5'ha : _T_719; // @[Lookup.scala 33:37]
  wire [4:0] _T_721 = _T_151 ? 5'ha : _T_720; // @[Lookup.scala 33:37]
  wire [4:0] _T_722 = _T_149 ? 5'hb : _T_721; // @[Lookup.scala 33:37]
  wire [4:0] _T_723 = _T_147 ? 5'hd : _T_722; // @[Lookup.scala 33:37]
  wire [4:0] _T_724 = _T_145 ? 5'ha : _T_723; // @[Lookup.scala 33:37]
  wire [4:0] _T_725 = _T_143 ? 5'hc : _T_724; // @[Lookup.scala 33:37]
  wire [4:0] _T_726 = _T_141 ? 5'hc : _T_725; // @[Lookup.scala 33:37]
  wire [4:0] _T_727 = _T_139 ? 5'h10 : _T_726; // @[Lookup.scala 33:37]
  wire [4:0] _T_728 = _T_137 ? 5'h5 : _T_727; // @[Lookup.scala 33:37]
  wire [4:0] _T_729 = _T_135 ? 5'h4 : _T_728; // @[Lookup.scala 33:37]
  wire [4:0] _T_730 = _T_133 ? 5'h7 : _T_729; // @[Lookup.scala 33:37]
  wire [4:0] _T_731 = _T_131 ? 5'h6 : _T_730; // @[Lookup.scala 33:37]
  wire [4:0] rvcImmType = _T_129 ? 5'he : _T_731; // @[Lookup.scala 33:37]
  wire [3:0] _T_732 = _T_193 ? 4'h9 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_733 = _T_191 ? 4'h9 : _T_732; // @[Lookup.scala 33:37]
  wire [3:0] _T_734 = _T_189 ? 4'h2 : _T_733; // @[Lookup.scala 33:37]
  wire [3:0] _T_735 = _T_187 ? 4'h4 : _T_734; // @[Lookup.scala 33:37]
  wire [3:0] _T_736 = _T_185 ? 4'h0 : _T_735; // @[Lookup.scala 33:37]
  wire [3:0] _T_737 = _T_183 ? 4'h5 : _T_736; // @[Lookup.scala 33:37]
  wire [3:0] _T_738 = _T_181 ? 4'h4 : _T_737; // @[Lookup.scala 33:37]
  wire [3:0] _T_739 = _T_179 ? 4'h9 : _T_738; // @[Lookup.scala 33:37]
  wire [3:0] _T_740 = _T_177 ? 4'h9 : _T_739; // @[Lookup.scala 33:37]
  wire [3:0] _T_741 = _T_175 ? 4'h2 : _T_740; // @[Lookup.scala 33:37]
  wire [3:0] _T_742 = _T_173 ? 4'h6 : _T_741; // @[Lookup.scala 33:37]
  wire [3:0] _T_743 = _T_171 ? 4'h6 : _T_742; // @[Lookup.scala 33:37]
  wire [3:0] _T_744 = _T_169 ? 4'h0 : _T_743; // @[Lookup.scala 33:37]
  wire [3:0] _T_745 = _T_167 ? 4'h6 : _T_744; // @[Lookup.scala 33:37]
  wire [3:0] _T_746 = _T_165 ? 4'h6 : _T_745; // @[Lookup.scala 33:37]
  wire [3:0] _T_747 = _T_163 ? 4'h6 : _T_746; // @[Lookup.scala 33:37]
  wire [3:0] _T_748 = _T_161 ? 4'h6 : _T_747; // @[Lookup.scala 33:37]
  wire [3:0] _T_749 = _T_159 ? 4'h6 : _T_748; // @[Lookup.scala 33:37]
  wire [3:0] _T_750 = _T_157 ? 4'h6 : _T_749; // @[Lookup.scala 33:37]
  wire [3:0] _T_751 = _T_155 ? 4'h6 : _T_750; // @[Lookup.scala 33:37]
  wire [3:0] _T_752 = _T_153 ? 4'h6 : _T_751; // @[Lookup.scala 33:37]
  wire [3:0] _T_753 = _T_151 ? 4'h6 : _T_752; // @[Lookup.scala 33:37]
  wire [3:0] _T_754 = _T_149 ? 4'h0 : _T_753; // @[Lookup.scala 33:37]
  wire [3:0] _T_755 = _T_147 ? 4'h9 : _T_754; // @[Lookup.scala 33:37]
  wire [3:0] _T_756 = _T_145 ? 4'h0 : _T_755; // @[Lookup.scala 33:37]
  wire [3:0] _T_757 = _T_143 ? 4'h2 : _T_756; // @[Lookup.scala 33:37]
  wire [3:0] _T_758 = _T_141 ? 4'h2 : _T_757; // @[Lookup.scala 33:37]
  wire [3:0] _T_759 = _T_139 ? 4'h0 : _T_758; // @[Lookup.scala 33:37]
  wire [3:0] _T_760 = _T_137 ? 4'h6 : _T_759; // @[Lookup.scala 33:37]
  wire [3:0] _T_761 = _T_135 ? 4'h6 : _T_760; // @[Lookup.scala 33:37]
  wire [3:0] _T_762 = _T_133 ? 4'h6 : _T_761; // @[Lookup.scala 33:37]
  wire [3:0] _T_763 = _T_131 ? 4'h6 : _T_762; // @[Lookup.scala 33:37]
  wire [3:0] rvcSrc1Type = _T_129 ? 4'h9 : _T_763; // @[Lookup.scala 33:37]
  wire [2:0] _T_764 = _T_193 ? 3'h5 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_765 = _T_191 ? 3'h5 : _T_764; // @[Lookup.scala 33:37]
  wire [2:0] _T_766 = _T_189 ? 3'h5 : _T_765; // @[Lookup.scala 33:37]
  wire [2:0] _T_767 = _T_187 ? 3'h0 : _T_766; // @[Lookup.scala 33:37]
  wire [2:0] _T_768 = _T_185 ? 3'h0 : _T_767; // @[Lookup.scala 33:37]
  wire [2:0] _T_769 = _T_183 ? 3'h0 : _T_768; // @[Lookup.scala 33:37]
  wire [2:0] _T_770 = _T_181 ? 3'h0 : _T_769; // @[Lookup.scala 33:37]
  wire [2:0] _T_771 = _T_179 ? 3'h0 : _T_770; // @[Lookup.scala 33:37]
  wire [2:0] _T_772 = _T_177 ? 3'h0 : _T_771; // @[Lookup.scala 33:37]
  wire [2:0] _T_773 = _T_175 ? 3'h0 : _T_772; // @[Lookup.scala 33:37]
  wire [2:0] _T_774 = _T_173 ? 3'h0 : _T_773; // @[Lookup.scala 33:37]
  wire [2:0] _T_775 = _T_171 ? 3'h0 : _T_774; // @[Lookup.scala 33:37]
  wire [2:0] _T_776 = _T_169 ? 3'h0 : _T_775; // @[Lookup.scala 33:37]
  wire [2:0] _T_777 = _T_167 ? 3'h7 : _T_776; // @[Lookup.scala 33:37]
  wire [2:0] _T_778 = _T_165 ? 3'h7 : _T_777; // @[Lookup.scala 33:37]
  wire [2:0] _T_779 = _T_163 ? 3'h7 : _T_778; // @[Lookup.scala 33:37]
  wire [2:0] _T_780 = _T_161 ? 3'h7 : _T_779; // @[Lookup.scala 33:37]
  wire [2:0] _T_781 = _T_159 ? 3'h7 : _T_780; // @[Lookup.scala 33:37]
  wire [2:0] _T_782 = _T_157 ? 3'h7 : _T_781; // @[Lookup.scala 33:37]
  wire [2:0] _T_783 = _T_155 ? 3'h0 : _T_782; // @[Lookup.scala 33:37]
  wire [2:0] _T_784 = _T_153 ? 3'h0 : _T_783; // @[Lookup.scala 33:37]
  wire [2:0] _T_785 = _T_151 ? 3'h0 : _T_784; // @[Lookup.scala 33:37]
  wire [2:0] _T_786 = _T_149 ? 3'h0 : _T_785; // @[Lookup.scala 33:37]
  wire [2:0] _T_787 = _T_147 ? 3'h0 : _T_786; // @[Lookup.scala 33:37]
  wire [2:0] _T_788 = _T_145 ? 3'h0 : _T_787; // @[Lookup.scala 33:37]
  wire [2:0] _T_789 = _T_143 ? 3'h0 : _T_788; // @[Lookup.scala 33:37]
  wire [2:0] _T_790 = _T_141 ? 3'h0 : _T_789; // @[Lookup.scala 33:37]
  wire [2:0] _T_791 = _T_139 ? 3'h0 : _T_790; // @[Lookup.scala 33:37]
  wire [2:0] _T_792 = _T_137 ? 3'h7 : _T_791; // @[Lookup.scala 33:37]
  wire [2:0] _T_793 = _T_135 ? 3'h7 : _T_792; // @[Lookup.scala 33:37]
  wire [2:0] _T_794 = _T_133 ? 3'h0 : _T_793; // @[Lookup.scala 33:37]
  wire [2:0] _T_795 = _T_131 ? 3'h0 : _T_794; // @[Lookup.scala 33:37]
  wire [2:0] rvcSrc2Type = _T_129 ? 3'h0 : _T_795; // @[Lookup.scala 33:37]
  wire [1:0] _T_798 = _T_189 ? 2'h2 : 2'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_799 = _T_187 ? 4'h8 : {{2'd0}, _T_798}; // @[Lookup.scala 33:37]
  wire [3:0] _T_800 = _T_185 ? 4'h0 : _T_799; // @[Lookup.scala 33:37]
  wire [3:0] _T_801 = _T_183 ? 4'h2 : _T_800; // @[Lookup.scala 33:37]
  wire [3:0] _T_802 = _T_181 ? 4'h0 : _T_801; // @[Lookup.scala 33:37]
  wire [3:0] _T_803 = _T_179 ? 4'h2 : _T_802; // @[Lookup.scala 33:37]
  wire [3:0] _T_804 = _T_177 ? 4'h2 : _T_803; // @[Lookup.scala 33:37]
  wire [3:0] _T_805 = _T_175 ? 4'h2 : _T_804; // @[Lookup.scala 33:37]
  wire [3:0] _T_806 = _T_173 ? 4'h0 : _T_805; // @[Lookup.scala 33:37]
  wire [3:0] _T_807 = _T_171 ? 4'h0 : _T_806; // @[Lookup.scala 33:37]
  wire [3:0] _T_808 = _T_169 ? 4'h0 : _T_807; // @[Lookup.scala 33:37]
  wire [3:0] _T_809 = _T_167 ? 4'h6 : _T_808; // @[Lookup.scala 33:37]
  wire [3:0] _T_810 = _T_165 ? 4'h6 : _T_809; // @[Lookup.scala 33:37]
  wire [3:0] _T_811 = _T_163 ? 4'h6 : _T_810; // @[Lookup.scala 33:37]
  wire [3:0] _T_812 = _T_161 ? 4'h6 : _T_811; // @[Lookup.scala 33:37]
  wire [3:0] _T_813 = _T_159 ? 4'h6 : _T_812; // @[Lookup.scala 33:37]
  wire [3:0] _T_814 = _T_157 ? 4'h6 : _T_813; // @[Lookup.scala 33:37]
  wire [3:0] _T_815 = _T_155 ? 4'h6 : _T_814; // @[Lookup.scala 33:37]
  wire [3:0] _T_816 = _T_153 ? 4'h6 : _T_815; // @[Lookup.scala 33:37]
  wire [3:0] _T_817 = _T_151 ? 4'h6 : _T_816; // @[Lookup.scala 33:37]
  wire [3:0] _T_818 = _T_149 ? 4'h2 : _T_817; // @[Lookup.scala 33:37]
  wire [3:0] _T_819 = _T_147 ? 4'h9 : _T_818; // @[Lookup.scala 33:37]
  wire [3:0] _T_820 = _T_145 ? 4'h2 : _T_819; // @[Lookup.scala 33:37]
  wire [3:0] _T_821 = _T_143 ? 4'h2 : _T_820; // @[Lookup.scala 33:37]
  wire [3:0] _T_822 = _T_141 ? 4'h2 : _T_821; // @[Lookup.scala 33:37]
  wire [3:0] _T_823 = _T_139 ? 4'h0 : _T_822; // @[Lookup.scala 33:37]
  wire [3:0] _T_824 = _T_137 ? 4'h0 : _T_823; // @[Lookup.scala 33:37]
  wire [3:0] _T_825 = _T_135 ? 4'h0 : _T_824; // @[Lookup.scala 33:37]
  wire [3:0] _T_826 = _T_133 ? 4'h7 : _T_825; // @[Lookup.scala 33:37]
  wire [3:0] _T_827 = _T_131 ? 4'h7 : _T_826; // @[Lookup.scala 33:37]
  wire [3:0] rvcDestType = _T_129 ? 4'h7 : _T_827; // @[Lookup.scala 33:37]
  wire  _T_828 = 4'h4 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_830 = 4'h2 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_831 = 4'hf == instrType; // @[LookupTree.scala 24:34]
  wire  _T_832 = 4'h1 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_833 = 4'h6 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_834 = 4'h7 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_835 = 4'h0 == instrType; // @[LookupTree.scala 24:34]
  wire  src1Type = _T_833 | _T_834 | _T_835; // @[Mux.scala 27:72]
  wire  src2Type = _T_828 | _T_833 | _T_834 | _T_835; // @[Mux.scala 27:72]
  wire [4:0] rs = io_in_bits_instr[19:15]; // @[IDU.scala 60:28]
  wire [4:0] rt = io_in_bits_instr[24:20]; // @[IDU.scala 60:43]
  wire [4:0] rd = io_in_bits_instr[11:7]; // @[IDU.scala 60:58]
  wire [4:0] rs2 = io_in_bits_instr[6:2]; // @[IDU.scala 63:24]
  wire  _T_875 = 3'h0 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_876 = 3'h1 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_877 = 3'h2 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_878 = 3'h3 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_879 = 3'h4 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_880 = 3'h5 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_881 = 3'h6 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_882 = 3'h7 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire [3:0] _T_883 = _T_875 ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_884 = _T_876 ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_885 = _T_877 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_886 = _T_878 ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_887 = _T_879 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_888 = _T_880 ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_889 = _T_881 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_890 = _T_882 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_891 = _T_883 | _T_884; // @[Mux.scala 27:72]
  wire [3:0] _T_892 = _T_891 | _T_885; // @[Mux.scala 27:72]
  wire [3:0] _T_893 = _T_892 | _T_886; // @[Mux.scala 27:72]
  wire [3:0] _T_894 = _T_893 | _T_887; // @[Mux.scala 27:72]
  wire [3:0] _T_895 = _T_894 | _T_888; // @[Mux.scala 27:72]
  wire [3:0] _T_896 = _T_895 | _T_889; // @[Mux.scala 27:72]
  wire [3:0] rs1p = _T_896 | _T_890; // @[Mux.scala 27:72]
  wire  _T_899 = 3'h0 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_900 = 3'h1 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_901 = 3'h2 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_902 = 3'h3 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_903 = 3'h4 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_904 = 3'h5 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_905 = 3'h6 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_906 = 3'h7 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire [3:0] _T_907 = _T_899 ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_908 = _T_900 ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_909 = _T_901 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_910 = _T_902 ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_911 = _T_903 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_912 = _T_904 ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_913 = _T_905 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_914 = _T_906 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_915 = _T_907 | _T_908; // @[Mux.scala 27:72]
  wire [3:0] _T_916 = _T_915 | _T_909; // @[Mux.scala 27:72]
  wire [3:0] _T_917 = _T_916 | _T_910; // @[Mux.scala 27:72]
  wire [3:0] _T_918 = _T_917 | _T_911; // @[Mux.scala 27:72]
  wire [3:0] _T_919 = _T_918 | _T_912; // @[Mux.scala 27:72]
  wire [3:0] _T_920 = _T_919 | _T_913; // @[Mux.scala 27:72]
  wire [3:0] rs2p = _T_920 | _T_914; // @[Mux.scala 27:72]
  wire  hi = io_in_bits_instr[12]; // @[IDU.scala 66:28]
  wire [5:0] rvc_shamt = {hi,rs2}; // @[Cat.scala 30:58]
  wire  _T_923 = 4'h3 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_924 = 4'h1 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_925 = 4'h2 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_926 = 4'h4 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_927 = 4'h5 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_928 = 4'h6 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_929 = 4'h7 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_930 = 4'h8 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_931 = 4'h9 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire [4:0] _T_933 = _T_923 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_934 = _T_924 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_935 = _T_925 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_936 = _T_926 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_937 = _T_927 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_938 = _T_928 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_939 = _T_929 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_941 = _T_931 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_943 = _T_933 | _T_934; // @[Mux.scala 27:72]
  wire [4:0] _T_944 = _T_943 | _T_935; // @[Mux.scala 27:72]
  wire [4:0] _T_945 = _T_944 | _T_936; // @[Mux.scala 27:72]
  wire [4:0] _T_946 = _T_945 | _T_937; // @[Mux.scala 27:72]
  wire [4:0] _GEN_5 = {{1'd0}, _T_938}; // @[Mux.scala 27:72]
  wire [4:0] _T_947 = _T_946 | _GEN_5; // @[Mux.scala 27:72]
  wire [4:0] _GEN_6 = {{1'd0}, _T_939}; // @[Mux.scala 27:72]
  wire [4:0] _T_948 = _T_947 | _GEN_6; // @[Mux.scala 27:72]
  wire [4:0] _GEN_7 = {{4'd0}, _T_930}; // @[Mux.scala 27:72]
  wire [4:0] _T_949 = _T_948 | _GEN_7; // @[Mux.scala 27:72]
  wire [4:0] _GEN_8 = {{3'd0}, _T_941}; // @[Mux.scala 27:72]
  wire [4:0] rvc_src1 = _T_949 | _GEN_8; // @[Mux.scala 27:72]
  wire  _T_952 = 3'h3 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_953 = 3'h1 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_954 = 3'h2 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_955 = 3'h4 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_956 = 3'h5 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_957 = 3'h6 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_958 = 3'h7 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire [3:0] _GEN_9 = {{1'd0}, rvcSrc2Type}; // @[LookupTree.scala 24:34]
  wire  _T_959 = 4'h8 == _GEN_9; // @[LookupTree.scala 24:34]
  wire  _T_960 = 4'h9 == _GEN_9; // @[LookupTree.scala 24:34]
  wire [4:0] _T_962 = _T_952 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_963 = _T_953 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_964 = _T_954 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_965 = _T_955 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_966 = _T_956 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_967 = _T_957 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_968 = _T_958 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_970 = _T_960 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_972 = _T_962 | _T_963; // @[Mux.scala 27:72]
  wire [4:0] _T_973 = _T_972 | _T_964; // @[Mux.scala 27:72]
  wire [4:0] _T_974 = _T_973 | _T_965; // @[Mux.scala 27:72]
  wire [4:0] _T_975 = _T_974 | _T_966; // @[Mux.scala 27:72]
  wire [4:0] _GEN_11 = {{1'd0}, _T_967}; // @[Mux.scala 27:72]
  wire [4:0] _T_976 = _T_975 | _GEN_11; // @[Mux.scala 27:72]
  wire [4:0] _GEN_12 = {{1'd0}, _T_968}; // @[Mux.scala 27:72]
  wire [4:0] _T_977 = _T_976 | _GEN_12; // @[Mux.scala 27:72]
  wire [4:0] _GEN_13 = {{4'd0}, _T_959}; // @[Mux.scala 27:72]
  wire [4:0] _T_978 = _T_977 | _GEN_13; // @[Mux.scala 27:72]
  wire [4:0] _GEN_14 = {{3'd0}, _T_970}; // @[Mux.scala 27:72]
  wire [4:0] rvc_src2 = _T_978 | _GEN_14; // @[Mux.scala 27:72]
  wire  _T_981 = 4'h3 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_982 = 4'h1 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_983 = 4'h2 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_984 = 4'h4 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_985 = 4'h5 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_986 = 4'h6 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_987 = 4'h7 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_988 = 4'h8 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_989 = 4'h9 == rvcDestType; // @[LookupTree.scala 24:34]
  wire [4:0] _T_991 = _T_981 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_992 = _T_982 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_993 = _T_983 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_994 = _T_984 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_995 = _T_985 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_996 = _T_986 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_997 = _T_987 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_999 = _T_989 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1001 = _T_991 | _T_992; // @[Mux.scala 27:72]
  wire [4:0] _T_1002 = _T_1001 | _T_993; // @[Mux.scala 27:72]
  wire [4:0] _T_1003 = _T_1002 | _T_994; // @[Mux.scala 27:72]
  wire [4:0] _T_1004 = _T_1003 | _T_995; // @[Mux.scala 27:72]
  wire [4:0] _GEN_15 = {{1'd0}, _T_996}; // @[Mux.scala 27:72]
  wire [4:0] _T_1005 = _T_1004 | _GEN_15; // @[Mux.scala 27:72]
  wire [4:0] _GEN_16 = {{1'd0}, _T_997}; // @[Mux.scala 27:72]
  wire [4:0] _T_1006 = _T_1005 | _GEN_16; // @[Mux.scala 27:72]
  wire [4:0] _GEN_17 = {{4'd0}, _T_988}; // @[Mux.scala 27:72]
  wire [4:0] _T_1007 = _T_1006 | _GEN_17; // @[Mux.scala 27:72]
  wire [4:0] _GEN_18 = {{3'd0}, _T_999}; // @[Mux.scala 27:72]
  wire [4:0] rvc_dest = _T_1007 | _GEN_18; // @[Mux.scala 27:72]
  wire [4:0] rfSrc1 = isRVC ? rvc_src1 : rs; // @[IDU.scala 87:19]
  wire [4:0] rfSrc2 = isRVC ? rvc_src2 : rt; // @[IDU.scala 88:19]
  wire [4:0] rfDest = isRVC ? rvc_dest : rd; // @[IDU.scala 89:19]
  wire [11:0] lo_1 = io_in_bits_instr[31:20]; // @[IDU.scala 99:29]
  wire [51:0] hi_1 = lo_1[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1018 = {hi_1,lo_1}; // @[Cat.scala 30:58]
  wire [6:0] hi_2 = io_in_bits_instr[31:25]; // @[IDU.scala 100:33]
  wire [11:0] lo_3 = {hi_2,rd}; // @[Cat.scala 30:58]
  wire [51:0] hi_3 = lo_3[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1021 = {hi_3,hi_2,rd}; // @[Cat.scala 30:58]
  wire  hi_hi_hi = io_in_bits_instr[31]; // @[IDU.scala 102:33]
  wire  hi_hi_lo = io_in_bits_instr[7]; // @[IDU.scala 102:44]
  wire [5:0] hi_lo = io_in_bits_instr[30:25]; // @[IDU.scala 102:54]
  wire [3:0] lo_hi = io_in_bits_instr[11:8]; // @[IDU.scala 102:69]
  wire [12:0] lo_7 = {hi_hi_hi,hi_hi_lo,hi_lo,lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire [50:0] hi_7 = lo_7[12] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1027 = {hi_7,hi_hi_hi,hi_hi_lo,hi_lo,lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire [19:0] hi_8 = io_in_bits_instr[31:12]; // @[IDU.scala 103:33]
  wire [31:0] lo_8 = {hi_8,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] hi_9 = lo_8[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1030 = {hi_9,hi_8,12'h0}; // @[Cat.scala 30:58]
  wire [7:0] hi_hi_lo_1 = io_in_bits_instr[19:12]; // @[IDU.scala 104:44]
  wire  hi_lo_1 = io_in_bits_instr[20]; // @[IDU.scala 104:59]
  wire [9:0] lo_hi_1 = io_in_bits_instr[30:21]; // @[IDU.scala 104:70]
  wire [20:0] lo_10 = {hi_hi_hi,hi_hi_lo_1,hi_lo_1,lo_hi_1,1'h0}; // @[Cat.scala 30:58]
  wire [42:0] hi_11 = lo_10[20] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1033 = {hi_11,hi_hi_hi,hi_hi_lo_1,hi_lo_1,lo_hi_1,1'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_1040 = _T_828 ? _T_1018 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1041 = _T_830 ? _T_1021 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1042 = _T_831 ? _T_1021 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1043 = _T_832 ? _T_1027 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1044 = _T_833 ? _T_1030 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1045 = _T_834 ? _T_1033 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1046 = _T_1040 | _T_1041; // @[Mux.scala 27:72]
  wire [63:0] _T_1047 = _T_1046 | _T_1042; // @[Mux.scala 27:72]
  wire [63:0] _T_1048 = _T_1047 | _T_1043; // @[Mux.scala 27:72]
  wire [63:0] _T_1049 = _T_1048 | _T_1044; // @[Mux.scala 27:72]
  wire [63:0] imm = _T_1049 | _T_1045; // @[Mux.scala 27:72]
  wire [1:0] hi_hi_2 = io_in_bits_instr[3:2]; // @[IDU.scala 109:43]
  wire [2:0] lo_hi_2 = io_in_bits_instr[6:4]; // @[IDU.scala 109:66]
  wire [63:0] _T_1051 = {56'h0,hi_hi_2,hi,lo_hi_2,2'h0}; // @[Cat.scala 30:58]
  wire [1:0] lo_hi_3 = io_in_bits_instr[6:5]; // @[IDU.scala 110:66]
  wire [63:0] _T_1052 = {55'h0,io_in_bits_instr[4:2],hi,lo_hi_3,3'h0}; // @[Cat.scala 30:58]
  wire [1:0] hi_hi_4 = io_in_bits_instr[8:7]; // @[IDU.scala 111:43]
  wire [3:0] hi_lo_4 = io_in_bits_instr[12:9]; // @[IDU.scala 111:55]
  wire [63:0] _T_1053 = {56'h0,hi_hi_4,hi_lo_4,2'h0}; // @[Cat.scala 30:58]
  wire [2:0] hi_lo_5 = io_in_bits_instr[12:10]; // @[IDU.scala 112:55]
  wire [63:0] _T_1054 = {55'h0,io_in_bits_instr[9:7],hi_lo_5,3'h0}; // @[Cat.scala 30:58]
  wire  hi_hi_6 = io_in_bits_instr[5]; // @[IDU.scala 113:43]
  wire  lo_hi_4 = io_in_bits_instr[6]; // @[IDU.scala 113:67]
  wire [63:0] _T_1055 = {57'h0,hi_hi_6,hi_lo_5,lo_hi_4,2'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_1056 = {56'h0,lo_hi_3,hi_lo_5,3'h0}; // @[Cat.scala 30:58]
  wire  hi_hi_hi_lo = io_in_bits_instr[8]; // @[IDU.scala 117:54]
  wire [1:0] hi_hi_lo_2 = io_in_bits_instr[10:9]; // @[IDU.scala 117:64]
  wire  lo_hi_hi = io_in_bits_instr[2]; // @[IDU.scala 117:97]
  wire  lo_hi_lo = io_in_bits_instr[11]; // @[IDU.scala 117:107]
  wire [2:0] lo_lo_hi = io_in_bits_instr[5:3]; // @[IDU.scala 117:118]
  wire [11:0] lo_24 = {hi,hi_hi_hi_lo,hi_hi_lo_2,lo_hi_4,hi_hi_lo,lo_hi_hi,lo_hi_lo,lo_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire [51:0] hi_21 = lo_24[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1061 = {hi_21,hi,hi_hi_hi_lo,hi_hi_lo_2,lo_hi_4,hi_hi_lo,lo_hi_hi,lo_hi_lo,lo_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire [1:0] lo_hi_hi_1 = io_in_bits_instr[11:10]; // @[IDU.scala 118:76]
  wire [1:0] lo_hi_lo_1 = io_in_bits_instr[4:3]; // @[IDU.scala 118:90]
  wire [8:0] lo_26 = {hi,lo_hi_3,lo_hi_hi,lo_hi_hi_1,lo_hi_lo_1,1'h0}; // @[Cat.scala 30:58]
  wire [54:0] hi_23 = lo_26[8] ? 55'h7fffffffffffff : 55'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1064 = {hi_23,hi,lo_hi_3,lo_hi_hi,lo_hi_hi_1,lo_hi_lo_1,1'h0}; // @[Cat.scala 30:58]
  wire [57:0] hi_25 = rvc_shamt[5] ? 58'h3ffffffffffffff : 58'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1067 = {hi_25,hi,rs2}; // @[Cat.scala 30:58]
  wire [17:0] lo_29 = {hi,rs2,12'h0}; // @[Cat.scala 30:58]
  wire [45:0] hi_27 = lo_29[17] ? 46'h3fffffffffff : 46'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1070 = {hi_27,hi,rs2,12'h0}; // @[Cat.scala 30:58]
  wire [9:0] lo_33 = {hi,lo_hi_lo_1,hi_hi_6,lo_hi_hi,lo_hi_4,4'h0}; // @[Cat.scala 30:58]
  wire [53:0] hi_31 = lo_33[9] ? 54'h3fffffffffffff : 54'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1076 = {hi_31,hi,lo_hi_lo_1,hi_hi_6,lo_hi_hi,lo_hi_4,4'h0}; // @[Cat.scala 30:58]
  wire [3:0] hi_hi_hi_5 = io_in_bits_instr[10:7]; // @[IDU.scala 123:44]
  wire [1:0] hi_hi_lo_5 = io_in_bits_instr[12:11]; // @[IDU.scala 123:57]
  wire [63:0] _T_1077 = {54'h0,hi_hi_hi_5,hi_hi_lo_5,hi_hi_6,lo_hi_4,2'h0}; // @[Cat.scala 30:58]
  wire  _T_1079 = 5'h0 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1080 = 5'h1 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1081 = 5'h2 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1082 = 5'h3 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1083 = 5'h4 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1084 = 5'h5 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1085 = 5'h6 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1086 = 5'h7 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1087 = 5'h8 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1088 = 5'h9 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1089 = 5'ha == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1090 = 5'hb == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1091 = 5'hc == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1092 = 5'hd == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1093 = 5'he == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1094 = 5'hf == rvcImmType; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1096 = _T_1079 ? _T_1051 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1097 = _T_1080 ? _T_1052 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1098 = _T_1081 ? _T_1053 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1099 = _T_1082 ? _T_1054 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1100 = _T_1083 ? _T_1055 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1101 = _T_1084 ? _T_1056 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1102 = _T_1085 ? _T_1055 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1103 = _T_1086 ? _T_1056 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1104 = _T_1087 ? _T_1061 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1105 = _T_1088 ? _T_1064 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1106 = _T_1089 ? _T_1067 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1107 = _T_1090 ? _T_1070 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1108 = _T_1091 ? _T_1067 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1109 = _T_1092 ? _T_1076 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1110 = _T_1093 ? _T_1077 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1111 = _T_1094 ? 64'h1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1113 = _T_1096 | _T_1097; // @[Mux.scala 27:72]
  wire [63:0] _T_1114 = _T_1113 | _T_1098; // @[Mux.scala 27:72]
  wire [63:0] _T_1115 = _T_1114 | _T_1099; // @[Mux.scala 27:72]
  wire [63:0] _T_1116 = _T_1115 | _T_1100; // @[Mux.scala 27:72]
  wire [63:0] _T_1117 = _T_1116 | _T_1101; // @[Mux.scala 27:72]
  wire [63:0] _T_1118 = _T_1117 | _T_1102; // @[Mux.scala 27:72]
  wire [63:0] _T_1119 = _T_1118 | _T_1103; // @[Mux.scala 27:72]
  wire [63:0] _T_1120 = _T_1119 | _T_1104; // @[Mux.scala 27:72]
  wire [63:0] _T_1121 = _T_1120 | _T_1105; // @[Mux.scala 27:72]
  wire [63:0] _T_1122 = _T_1121 | _T_1106; // @[Mux.scala 27:72]
  wire [63:0] _T_1123 = _T_1122 | _T_1107; // @[Mux.scala 27:72]
  wire [63:0] _T_1124 = _T_1123 | _T_1108; // @[Mux.scala 27:72]
  wire [63:0] _T_1125 = _T_1124 | _T_1109; // @[Mux.scala 27:72]
  wire [63:0] _T_1126 = _T_1125 | _T_1110; // @[Mux.scala 27:72]
  wire [63:0] immrvc = _T_1126 | _T_1111; // @[Mux.scala 27:72]
  wire  _T_1132 = rfDest == 5'h1 | rfDest == 5'h5; // @[IDU.scala 131:42]
  wire [6:0] _GEN_0 = _T_1132 & fuOpType == 7'h58 ? 7'h5c : fuOpType; // @[IDU.scala 132:57 IDU.scala 132:85 IDU.scala 45:29]
  wire  _T_1138 = rfSrc1 == 5'h1 | rfSrc1 == 5'h5; // @[IDU.scala 131:42]
  wire [6:0] _GEN_1 = _T_1138 ? 7'h5e : _GEN_0; // @[IDU.scala 134:29 IDU.scala 134:57]
  wire [6:0] _GEN_2 = _T_1132 ? 7'h5c : _GEN_1; // @[IDU.scala 135:29 IDU.scala 135:57]
  wire [6:0] _GEN_3 = fuOpType == 7'h5a ? _GEN_2 : _GEN_0; // @[IDU.scala 133:40]
  wire  _T_1156 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_1157 = ~hasIntr; // @[IDU.scala 160:51]
  assign io_in_ready = ~io_in_valid | _T_1156 & ~hasIntr; // @[IDU.scala 160:31]
  assign io_out_valid = io_in_valid; // @[IDU.scala 159:16]
  assign io_out_bits_cf_instr = io_in_bits_instr; // @[IDU.scala 161:18]
  assign io_out_bits_cf_pc = io_in_bits_pc; // @[IDU.scala 161:18]
  assign io_out_bits_cf_pnpc = io_in_bits_pnpc; // @[IDU.scala 161:18]
  assign io_out_bits_cf_exceptionVec_1 = |io_in_bits_pc[38:32] & ~DTLBENABLE; // @[IDU.scala 179:98]
  assign io_out_bits_cf_exceptionVec_2 = instrType == 4'h0 & _T_1157 & io_in_valid; // @[IDU.scala 176:83]
  assign io_out_bits_cf_exceptionVec_12 = io_in_bits_exceptionVec_12; // @[IDU.scala 177:47]
  assign io_out_bits_cf_intrVec_0 = intrVecIDU[0]; // @[IDU.scala 169:38]
  assign io_out_bits_cf_intrVec_1 = intrVecIDU[1]; // @[IDU.scala 169:38]
  assign io_out_bits_cf_intrVec_2 = intrVecIDU[2]; // @[IDU.scala 169:38]
  assign io_out_bits_cf_intrVec_3 = intrVecIDU[3]; // @[IDU.scala 169:38]
  assign io_out_bits_cf_intrVec_4 = intrVecIDU[4]; // @[IDU.scala 169:38]
  assign io_out_bits_cf_intrVec_5 = intrVecIDU[5]; // @[IDU.scala 169:38]
  assign io_out_bits_cf_intrVec_6 = intrVecIDU[6]; // @[IDU.scala 169:38]
  assign io_out_bits_cf_intrVec_7 = intrVecIDU[7]; // @[IDU.scala 169:38]
  assign io_out_bits_cf_intrVec_8 = intrVecIDU[8]; // @[IDU.scala 169:38]
  assign io_out_bits_cf_intrVec_9 = intrVecIDU[9]; // @[IDU.scala 169:38]
  assign io_out_bits_cf_intrVec_10 = intrVecIDU[10]; // @[IDU.scala 169:38]
  assign io_out_bits_cf_intrVec_11 = intrVecIDU[11]; // @[IDU.scala 169:38]
  assign io_out_bits_cf_brIdx = io_in_bits_brIdx; // @[IDU.scala 161:18]
  assign io_out_bits_cf_crossPageIPFFix = io_in_bits_crossPageIPFFix; // @[IDU.scala 161:18]
  assign io_out_bits_ctrl_src1Type = io_in_bits_instr[6:0] == 7'h37 ? 1'h0 : src1Type; // @[IDU.scala 139:35]
  assign io_out_bits_ctrl_src2Type = _T_828 | _T_833 | _T_834 | _T_835; // @[Mux.scala 27:72]
  assign io_out_bits_ctrl_fuType = hasIntr | io_in_bits_exceptionVec_12 | io_out_bits_cf_exceptionVec_1 ? 3'h3 :
    decodeList_1; // @[IDU.scala 36:75]
  assign io_out_bits_ctrl_fuOpType = fuType == 3'h0 ? _GEN_3 : fuOpType; // @[IDU.scala 130:32 IDU.scala 45:29]
  assign io_out_bits_ctrl_rfSrc1 = src1Type ? 5'h0 : rfSrc1; // @[IDU.scala 92:33]
  assign io_out_bits_ctrl_rfSrc2 = ~src2Type ? rfSrc2 : 5'h0; // @[IDU.scala 93:33]
  assign io_out_bits_ctrl_rfWen = instrType[2]; // @[Decode.scala 33:50]
  assign io_out_bits_ctrl_rfDest = instrType[2] ? rfDest : 5'h0; // @[IDU.scala 95:33]
  assign io_out_bits_data_imm = isRVC ? immrvc : imm; // @[IDU.scala 128:31]
endmodule
module ysyx_210000_IDU(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_instr,
  input  [38:0] io_in_0_bits_pc,
  input  [38:0] io_in_0_bits_pnpc,
  input         io_in_0_bits_exceptionVec_12,
  input  [3:0]  io_in_0_bits_brIdx,
  input         io_in_0_bits_crossPageIPFFix,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [63:0] io_out_0_bits_cf_instr,
  output [38:0] io_out_0_bits_cf_pc,
  output [38:0] io_out_0_bits_cf_pnpc,
  output        io_out_0_bits_cf_exceptionVec_1,
  output        io_out_0_bits_cf_exceptionVec_2,
  output        io_out_0_bits_cf_exceptionVec_12,
  output        io_out_0_bits_cf_intrVec_0,
  output        io_out_0_bits_cf_intrVec_1,
  output        io_out_0_bits_cf_intrVec_2,
  output        io_out_0_bits_cf_intrVec_3,
  output        io_out_0_bits_cf_intrVec_4,
  output        io_out_0_bits_cf_intrVec_5,
  output        io_out_0_bits_cf_intrVec_6,
  output        io_out_0_bits_cf_intrVec_7,
  output        io_out_0_bits_cf_intrVec_8,
  output        io_out_0_bits_cf_intrVec_9,
  output        io_out_0_bits_cf_intrVec_10,
  output        io_out_0_bits_cf_intrVec_11,
  output [3:0]  io_out_0_bits_cf_brIdx,
  output        io_out_0_bits_cf_crossPageIPFFix,
  output        io_out_0_bits_ctrl_src1Type,
  output        io_out_0_bits_ctrl_src2Type,
  output [2:0]  io_out_0_bits_ctrl_fuType,
  output [6:0]  io_out_0_bits_ctrl_fuOpType,
  output [4:0]  io_out_0_bits_ctrl_rfSrc1,
  output [4:0]  io_out_0_bits_ctrl_rfSrc2,
  output        io_out_0_bits_ctrl_rfWen,
  output [4:0]  io_out_0_bits_ctrl_rfDest,
  output [63:0] io_out_0_bits_data_imm,
  input         io_out_1_ready,
  output        io_out_1_valid,
  output [63:0] io_out_1_bits_cf_instr,
  output [38:0] io_out_1_bits_cf_pc,
  output [38:0] io_out_1_bits_cf_pnpc,
  output        io_out_1_bits_cf_exceptionVec_1,
  output        io_out_1_bits_cf_exceptionVec_2,
  output        io_out_1_bits_cf_exceptionVec_12,
  output        io_out_1_bits_cf_intrVec_0,
  output        io_out_1_bits_cf_intrVec_1,
  output        io_out_1_bits_cf_intrVec_2,
  output        io_out_1_bits_cf_intrVec_3,
  output        io_out_1_bits_cf_intrVec_4,
  output        io_out_1_bits_cf_intrVec_5,
  output        io_out_1_bits_cf_intrVec_6,
  output        io_out_1_bits_cf_intrVec_7,
  output        io_out_1_bits_cf_intrVec_8,
  output        io_out_1_bits_cf_intrVec_9,
  output        io_out_1_bits_cf_intrVec_10,
  output        io_out_1_bits_cf_intrVec_11,
  output [3:0]  io_out_1_bits_cf_brIdx,
  output        io_out_1_bits_cf_crossPageIPFFix,
  output        io_out_1_bits_ctrl_src1Type,
  output        io_out_1_bits_ctrl_src2Type,
  output [2:0]  io_out_1_bits_ctrl_fuType,
  output [6:0]  io_out_1_bits_ctrl_fuOpType,
  output [4:0]  io_out_1_bits_ctrl_rfSrc1,
  output [4:0]  io_out_1_bits_ctrl_rfSrc2,
  output        io_out_1_bits_ctrl_rfWen,
  output [4:0]  io_out_1_bits_ctrl_rfDest,
  output [63:0] io_out_1_bits_data_imm,
  input         vmEnable,
  input  [11:0] intrVec
);
  wire  decoder1_io_in_ready; // @[IDU.scala 194:25]
  wire  decoder1_io_in_valid; // @[IDU.scala 194:25]
  wire [63:0] decoder1_io_in_bits_instr; // @[IDU.scala 194:25]
  wire [38:0] decoder1_io_in_bits_pc; // @[IDU.scala 194:25]
  wire [38:0] decoder1_io_in_bits_pnpc; // @[IDU.scala 194:25]
  wire  decoder1_io_in_bits_exceptionVec_12; // @[IDU.scala 194:25]
  wire [3:0] decoder1_io_in_bits_brIdx; // @[IDU.scala 194:25]
  wire  decoder1_io_in_bits_crossPageIPFFix; // @[IDU.scala 194:25]
  wire  decoder1_io_out_ready; // @[IDU.scala 194:25]
  wire  decoder1_io_out_valid; // @[IDU.scala 194:25]
  wire [63:0] decoder1_io_out_bits_cf_instr; // @[IDU.scala 194:25]
  wire [38:0] decoder1_io_out_bits_cf_pc; // @[IDU.scala 194:25]
  wire [38:0] decoder1_io_out_bits_cf_pnpc; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_1; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_2; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_12; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_0; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_1; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_2; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_3; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_4; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_5; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_6; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_7; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_8; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_9; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_10; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_11; // @[IDU.scala 194:25]
  wire [3:0] decoder1_io_out_bits_cf_brIdx; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_crossPageIPFFix; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_ctrl_src1Type; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_ctrl_src2Type; // @[IDU.scala 194:25]
  wire [2:0] decoder1_io_out_bits_ctrl_fuType; // @[IDU.scala 194:25]
  wire [6:0] decoder1_io_out_bits_ctrl_fuOpType; // @[IDU.scala 194:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc1; // @[IDU.scala 194:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc2; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_ctrl_rfWen; // @[IDU.scala 194:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfDest; // @[IDU.scala 194:25]
  wire [63:0] decoder1_io_out_bits_data_imm; // @[IDU.scala 194:25]
  wire  decoder1_DTLBENABLE; // @[IDU.scala 194:25]
  wire [11:0] decoder1_intrVecIDU; // @[IDU.scala 194:25]
  wire  decoder2_io_in_ready; // @[IDU.scala 195:25]
  wire  decoder2_io_in_valid; // @[IDU.scala 195:25]
  wire [63:0] decoder2_io_in_bits_instr; // @[IDU.scala 195:25]
  wire [38:0] decoder2_io_in_bits_pc; // @[IDU.scala 195:25]
  wire [38:0] decoder2_io_in_bits_pnpc; // @[IDU.scala 195:25]
  wire  decoder2_io_in_bits_exceptionVec_12; // @[IDU.scala 195:25]
  wire [3:0] decoder2_io_in_bits_brIdx; // @[IDU.scala 195:25]
  wire  decoder2_io_in_bits_crossPageIPFFix; // @[IDU.scala 195:25]
  wire  decoder2_io_out_ready; // @[IDU.scala 195:25]
  wire  decoder2_io_out_valid; // @[IDU.scala 195:25]
  wire [63:0] decoder2_io_out_bits_cf_instr; // @[IDU.scala 195:25]
  wire [38:0] decoder2_io_out_bits_cf_pc; // @[IDU.scala 195:25]
  wire [38:0] decoder2_io_out_bits_cf_pnpc; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_exceptionVec_1; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_exceptionVec_2; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_exceptionVec_12; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_0; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_1; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_2; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_3; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_4; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_5; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_6; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_7; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_8; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_9; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_10; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_11; // @[IDU.scala 195:25]
  wire [3:0] decoder2_io_out_bits_cf_brIdx; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_crossPageIPFFix; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_ctrl_src1Type; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_ctrl_src2Type; // @[IDU.scala 195:25]
  wire [2:0] decoder2_io_out_bits_ctrl_fuType; // @[IDU.scala 195:25]
  wire [6:0] decoder2_io_out_bits_ctrl_fuOpType; // @[IDU.scala 195:25]
  wire [4:0] decoder2_io_out_bits_ctrl_rfSrc1; // @[IDU.scala 195:25]
  wire [4:0] decoder2_io_out_bits_ctrl_rfSrc2; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_ctrl_rfWen; // @[IDU.scala 195:25]
  wire [4:0] decoder2_io_out_bits_ctrl_rfDest; // @[IDU.scala 195:25]
  wire [63:0] decoder2_io_out_bits_data_imm; // @[IDU.scala 195:25]
  wire  decoder2_DTLBENABLE; // @[IDU.scala 195:25]
  wire [11:0] decoder2_intrVecIDU; // @[IDU.scala 195:25]
  ysyx_210000_Decoder decoder1 ( // @[IDU.scala 194:25]
    .io_in_ready(decoder1_io_in_ready),
    .io_in_valid(decoder1_io_in_valid),
    .io_in_bits_instr(decoder1_io_in_bits_instr),
    .io_in_bits_pc(decoder1_io_in_bits_pc),
    .io_in_bits_pnpc(decoder1_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_12(decoder1_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(decoder1_io_in_bits_brIdx),
    .io_in_bits_crossPageIPFFix(decoder1_io_in_bits_crossPageIPFFix),
    .io_out_ready(decoder1_io_out_ready),
    .io_out_valid(decoder1_io_out_valid),
    .io_out_bits_cf_instr(decoder1_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(decoder1_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(decoder1_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(decoder1_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(decoder1_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(decoder1_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_0(decoder1_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(decoder1_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(decoder1_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(decoder1_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(decoder1_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(decoder1_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(decoder1_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(decoder1_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(decoder1_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(decoder1_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(decoder1_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(decoder1_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(decoder1_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossPageIPFFix(decoder1_io_out_bits_cf_crossPageIPFFix),
    .io_out_bits_ctrl_src1Type(decoder1_io_out_bits_ctrl_src1Type),
    .io_out_bits_ctrl_src2Type(decoder1_io_out_bits_ctrl_src2Type),
    .io_out_bits_ctrl_fuType(decoder1_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(decoder1_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfSrc1(decoder1_io_out_bits_ctrl_rfSrc1),
    .io_out_bits_ctrl_rfSrc2(decoder1_io_out_bits_ctrl_rfSrc2),
    .io_out_bits_ctrl_rfWen(decoder1_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(decoder1_io_out_bits_ctrl_rfDest),
    .io_out_bits_data_imm(decoder1_io_out_bits_data_imm),
    .DTLBENABLE(decoder1_DTLBENABLE),
    .intrVecIDU(decoder1_intrVecIDU)
  );
  ysyx_210000_Decoder decoder2 ( // @[IDU.scala 195:25]
    .io_in_ready(decoder2_io_in_ready),
    .io_in_valid(decoder2_io_in_valid),
    .io_in_bits_instr(decoder2_io_in_bits_instr),
    .io_in_bits_pc(decoder2_io_in_bits_pc),
    .io_in_bits_pnpc(decoder2_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_12(decoder2_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(decoder2_io_in_bits_brIdx),
    .io_in_bits_crossPageIPFFix(decoder2_io_in_bits_crossPageIPFFix),
    .io_out_ready(decoder2_io_out_ready),
    .io_out_valid(decoder2_io_out_valid),
    .io_out_bits_cf_instr(decoder2_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(decoder2_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(decoder2_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(decoder2_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(decoder2_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(decoder2_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_0(decoder2_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(decoder2_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(decoder2_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(decoder2_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(decoder2_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(decoder2_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(decoder2_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(decoder2_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(decoder2_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(decoder2_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(decoder2_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(decoder2_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(decoder2_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossPageIPFFix(decoder2_io_out_bits_cf_crossPageIPFFix),
    .io_out_bits_ctrl_src1Type(decoder2_io_out_bits_ctrl_src1Type),
    .io_out_bits_ctrl_src2Type(decoder2_io_out_bits_ctrl_src2Type),
    .io_out_bits_ctrl_fuType(decoder2_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(decoder2_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfSrc1(decoder2_io_out_bits_ctrl_rfSrc1),
    .io_out_bits_ctrl_rfSrc2(decoder2_io_out_bits_ctrl_rfSrc2),
    .io_out_bits_ctrl_rfWen(decoder2_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(decoder2_io_out_bits_ctrl_rfDest),
    .io_out_bits_data_imm(decoder2_io_out_bits_data_imm),
    .DTLBENABLE(decoder2_DTLBENABLE),
    .intrVecIDU(decoder2_intrVecIDU)
  );
  assign io_in_0_ready = decoder1_io_in_ready; // @[IDU.scala 196:12]
  assign io_out_0_valid = decoder1_io_out_valid; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_instr = decoder1_io_out_bits_cf_instr; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_pc = decoder1_io_out_bits_cf_pc; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_pnpc = decoder1_io_out_bits_cf_pnpc; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_exceptionVec_1 = decoder1_io_out_bits_cf_exceptionVec_1; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_exceptionVec_2 = decoder1_io_out_bits_cf_exceptionVec_2; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_exceptionVec_12 = decoder1_io_out_bits_cf_exceptionVec_12; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_0 = decoder1_io_out_bits_cf_intrVec_0; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_1 = decoder1_io_out_bits_cf_intrVec_1; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_2 = decoder1_io_out_bits_cf_intrVec_2; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_3 = decoder1_io_out_bits_cf_intrVec_3; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_4 = decoder1_io_out_bits_cf_intrVec_4; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_5 = decoder1_io_out_bits_cf_intrVec_5; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_6 = decoder1_io_out_bits_cf_intrVec_6; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_7 = decoder1_io_out_bits_cf_intrVec_7; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_8 = decoder1_io_out_bits_cf_intrVec_8; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_9 = decoder1_io_out_bits_cf_intrVec_9; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_10 = decoder1_io_out_bits_cf_intrVec_10; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_11 = decoder1_io_out_bits_cf_intrVec_11; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_brIdx = decoder1_io_out_bits_cf_brIdx; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_crossPageIPFFix = decoder1_io_out_bits_cf_crossPageIPFFix; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_src1Type = decoder1_io_out_bits_ctrl_src1Type; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_src2Type = decoder1_io_out_bits_ctrl_src2Type; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_fuType = decoder1_io_out_bits_ctrl_fuType; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_fuOpType = decoder1_io_out_bits_ctrl_fuOpType; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_rfSrc1 = decoder1_io_out_bits_ctrl_rfSrc1; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_rfSrc2 = decoder1_io_out_bits_ctrl_rfSrc2; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_rfWen = decoder1_io_out_bits_ctrl_rfWen; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_rfDest = decoder1_io_out_bits_ctrl_rfDest; // @[IDU.scala 198:13]
  assign io_out_0_bits_data_imm = decoder1_io_out_bits_data_imm; // @[IDU.scala 198:13]
  assign io_out_1_valid = decoder2_io_out_valid; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_instr = decoder2_io_out_bits_cf_instr; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_pc = decoder2_io_out_bits_cf_pc; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_pnpc = decoder2_io_out_bits_cf_pnpc; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_exceptionVec_1 = decoder2_io_out_bits_cf_exceptionVec_1; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_exceptionVec_2 = decoder2_io_out_bits_cf_exceptionVec_2; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_exceptionVec_12 = decoder2_io_out_bits_cf_exceptionVec_12; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_0 = decoder2_io_out_bits_cf_intrVec_0; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_1 = decoder2_io_out_bits_cf_intrVec_1; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_2 = decoder2_io_out_bits_cf_intrVec_2; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_3 = decoder2_io_out_bits_cf_intrVec_3; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_4 = decoder2_io_out_bits_cf_intrVec_4; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_5 = decoder2_io_out_bits_cf_intrVec_5; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_6 = decoder2_io_out_bits_cf_intrVec_6; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_7 = decoder2_io_out_bits_cf_intrVec_7; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_8 = decoder2_io_out_bits_cf_intrVec_8; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_9 = decoder2_io_out_bits_cf_intrVec_9; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_10 = decoder2_io_out_bits_cf_intrVec_10; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_11 = decoder2_io_out_bits_cf_intrVec_11; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_brIdx = decoder2_io_out_bits_cf_brIdx; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_crossPageIPFFix = decoder2_io_out_bits_cf_crossPageIPFFix; // @[IDU.scala 199:13]
  assign io_out_1_bits_ctrl_src1Type = decoder2_io_out_bits_ctrl_src1Type; // @[IDU.scala 199:13]
  assign io_out_1_bits_ctrl_src2Type = decoder2_io_out_bits_ctrl_src2Type; // @[IDU.scala 199:13]
  assign io_out_1_bits_ctrl_fuType = decoder2_io_out_bits_ctrl_fuType; // @[IDU.scala 199:13]
  assign io_out_1_bits_ctrl_fuOpType = decoder2_io_out_bits_ctrl_fuOpType; // @[IDU.scala 199:13]
  assign io_out_1_bits_ctrl_rfSrc1 = decoder2_io_out_bits_ctrl_rfSrc1; // @[IDU.scala 199:13]
  assign io_out_1_bits_ctrl_rfSrc2 = decoder2_io_out_bits_ctrl_rfSrc2; // @[IDU.scala 199:13]
  assign io_out_1_bits_ctrl_rfWen = decoder2_io_out_bits_ctrl_rfWen; // @[IDU.scala 199:13]
  assign io_out_1_bits_ctrl_rfDest = decoder2_io_out_bits_ctrl_rfDest; // @[IDU.scala 199:13]
  assign io_out_1_bits_data_imm = decoder2_io_out_bits_data_imm; // @[IDU.scala 199:13]
  assign decoder1_io_in_valid = io_in_0_valid; // @[IDU.scala 196:12]
  assign decoder1_io_in_bits_instr = io_in_0_bits_instr; // @[IDU.scala 196:12]
  assign decoder1_io_in_bits_pc = io_in_0_bits_pc; // @[IDU.scala 196:12]
  assign decoder1_io_in_bits_pnpc = io_in_0_bits_pnpc; // @[IDU.scala 196:12]
  assign decoder1_io_in_bits_exceptionVec_12 = io_in_0_bits_exceptionVec_12; // @[IDU.scala 196:12]
  assign decoder1_io_in_bits_brIdx = io_in_0_bits_brIdx; // @[IDU.scala 196:12]
  assign decoder1_io_in_bits_crossPageIPFFix = io_in_0_bits_crossPageIPFFix; // @[IDU.scala 196:12]
  assign decoder1_io_out_ready = io_out_0_ready; // @[IDU.scala 198:13]
  assign decoder1_DTLBENABLE = vmEnable;
  assign decoder1_intrVecIDU = intrVec;
  assign decoder2_io_in_valid = 1'h0; // @[IDU.scala 202:26]
  assign decoder2_io_in_bits_instr = 64'h0; // @[IDU.scala 197:12]
  assign decoder2_io_in_bits_pc = 39'h0; // @[IDU.scala 197:12]
  assign decoder2_io_in_bits_pnpc = 39'h0; // @[IDU.scala 197:12]
  assign decoder2_io_in_bits_exceptionVec_12 = 1'h0; // @[IDU.scala 197:12]
  assign decoder2_io_in_bits_brIdx = 4'h0; // @[IDU.scala 197:12]
  assign decoder2_io_in_bits_crossPageIPFFix = 1'h0; // @[IDU.scala 197:12]
  assign decoder2_io_out_ready = io_out_1_ready; // @[IDU.scala 199:13]
  assign decoder2_DTLBENABLE = vmEnable;
  assign decoder2_intrVecIDU = intrVec;
endmodule
module ysyx_210000_FlushableQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_instr,
  input  [38:0] io_enq_bits_pc,
  input  [38:0] io_enq_bits_pnpc,
  input         io_enq_bits_exceptionVec_12,
  input  [3:0]  io_enq_bits_brIdx,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_instr,
  output [38:0] io_deq_bits_pc,
  output [38:0] io_deq_bits_pnpc,
  output        io_deq_bits_exceptionVec_12,
  output [3:0]  io_deq_bits_brIdx,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] REG__0_instr; // @[FlushableQueue.scala 34:28]
  reg [38:0] REG__0_pc; // @[FlushableQueue.scala 34:28]
  reg [38:0] REG__0_pnpc; // @[FlushableQueue.scala 34:28]
  reg  REG__0_exceptionVec_12; // @[FlushableQueue.scala 34:28]
  reg [3:0] REG__0_brIdx; // @[FlushableQueue.scala 34:28]
  reg [63:0] REG__1_instr; // @[FlushableQueue.scala 34:28]
  reg [38:0] REG__1_pc; // @[FlushableQueue.scala 34:28]
  reg [38:0] REG__1_pnpc; // @[FlushableQueue.scala 34:28]
  reg  REG__1_exceptionVec_12; // @[FlushableQueue.scala 34:28]
  reg [3:0] REG__1_brIdx; // @[FlushableQueue.scala 34:28]
  reg [63:0] REG__2_instr; // @[FlushableQueue.scala 34:28]
  reg [38:0] REG__2_pc; // @[FlushableQueue.scala 34:28]
  reg [38:0] REG__2_pnpc; // @[FlushableQueue.scala 34:28]
  reg  REG__2_exceptionVec_12; // @[FlushableQueue.scala 34:28]
  reg [3:0] REG__2_brIdx; // @[FlushableQueue.scala 34:28]
  reg [63:0] REG__3_instr; // @[FlushableQueue.scala 34:28]
  reg [38:0] REG__3_pc; // @[FlushableQueue.scala 34:28]
  reg [38:0] REG__3_pnpc; // @[FlushableQueue.scala 34:28]
  reg  REG__3_exceptionVec_12; // @[FlushableQueue.scala 34:28]
  reg [3:0] REG__3_brIdx; // @[FlushableQueue.scala 34:28]
  reg [1:0] value; // @[Counter.scala 60:40]
  reg [1:0] value_1; // @[Counter.scala 60:40]
  reg  REG_1; // @[FlushableQueue.scala 37:35]
  wire  _T = value == value_1; // @[FlushableQueue.scala 39:41]
  wire  _T_2 = _T & ~REG_1; // @[FlushableQueue.scala 40:33]
  wire  _T_3 = _T & REG_1; // @[FlushableQueue.scala 41:32]
  wire  _T_4 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_5 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _value_T_1 = value + 2'h1; // @[Counter.scala 76:24]
  wire [1:0] _value_T_3 = value_1 + 2'h1; // @[Counter.scala 76:24]
  wire [3:0] _GEN_356 = 2'h1 == value_1 ? REG__1_brIdx : REG__0_brIdx; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  wire [3:0] _GEN_357 = 2'h2 == value_1 ? REG__2_brIdx : _GEN_356; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  wire  _GEN_456 = 2'h1 == value_1 ? REG__1_exceptionVec_12 : REG__0_exceptionVec_12; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  wire  _GEN_457 = 2'h2 == value_1 ? REG__2_exceptionVec_12 : _GEN_456; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  wire [38:0] _GEN_508 = 2'h1 == value_1 ? REG__1_pnpc : REG__0_pnpc; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  wire [38:0] _GEN_509 = 2'h2 == value_1 ? REG__2_pnpc : _GEN_508; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  wire [38:0] _GEN_512 = 2'h1 == value_1 ? REG__1_pc : REG__0_pc; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  wire [38:0] _GEN_513 = 2'h2 == value_1 ? REG__2_pc : _GEN_512; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  wire [63:0] _GEN_516 = 2'h1 == value_1 ? REG__1_instr : REG__0_instr; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  wire [63:0] _GEN_517 = 2'h2 == value_1 ? REG__2_instr : _GEN_516; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  assign io_enq_ready = ~_T_3; // @[FlushableQueue.scala 57:19]
  assign io_deq_valid = ~_T_2; // @[FlushableQueue.scala 56:19]
  assign io_deq_bits_instr = 2'h3 == value_1 ? REG__3_instr : _GEN_517; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  assign io_deq_bits_pc = 2'h3 == value_1 ? REG__3_pc : _GEN_513; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  assign io_deq_bits_pnpc = 2'h3 == value_1 ? REG__3_pnpc : _GEN_509; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  assign io_deq_bits_exceptionVec_12 = 2'h3 == value_1 ? REG__3_exceptionVec_12 : _GEN_457; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  assign io_deq_bits_brIdx = 2'h3 == value_1 ? REG__3_brIdx : _GEN_357; // @[FlushableQueue.scala 58:15 FlushableQueue.scala 58:15]
  always @(posedge clock) begin
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__0_instr <= 64'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h0 == value) begin // @[FlushableQueue.scala 46:24]
        REG__0_instr <= io_enq_bits_instr; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__0_pc <= 39'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h0 == value) begin // @[FlushableQueue.scala 46:24]
        REG__0_pc <= io_enq_bits_pc; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__0_pnpc <= 39'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h0 == value) begin // @[FlushableQueue.scala 46:24]
        REG__0_pnpc <= io_enq_bits_pnpc; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__0_exceptionVec_12 <= 1'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h0 == value) begin // @[FlushableQueue.scala 46:24]
        REG__0_exceptionVec_12 <= io_enq_bits_exceptionVec_12; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__0_brIdx <= 4'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h0 == value) begin // @[FlushableQueue.scala 46:24]
        REG__0_brIdx <= io_enq_bits_brIdx; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__1_instr <= 64'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h1 == value) begin // @[FlushableQueue.scala 46:24]
        REG__1_instr <= io_enq_bits_instr; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__1_pc <= 39'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h1 == value) begin // @[FlushableQueue.scala 46:24]
        REG__1_pc <= io_enq_bits_pc; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__1_pnpc <= 39'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h1 == value) begin // @[FlushableQueue.scala 46:24]
        REG__1_pnpc <= io_enq_bits_pnpc; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__1_exceptionVec_12 <= 1'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h1 == value) begin // @[FlushableQueue.scala 46:24]
        REG__1_exceptionVec_12 <= io_enq_bits_exceptionVec_12; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__1_brIdx <= 4'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h1 == value) begin // @[FlushableQueue.scala 46:24]
        REG__1_brIdx <= io_enq_bits_brIdx; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__2_instr <= 64'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h2 == value) begin // @[FlushableQueue.scala 46:24]
        REG__2_instr <= io_enq_bits_instr; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__2_pc <= 39'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h2 == value) begin // @[FlushableQueue.scala 46:24]
        REG__2_pc <= io_enq_bits_pc; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__2_pnpc <= 39'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h2 == value) begin // @[FlushableQueue.scala 46:24]
        REG__2_pnpc <= io_enq_bits_pnpc; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__2_exceptionVec_12 <= 1'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h2 == value) begin // @[FlushableQueue.scala 46:24]
        REG__2_exceptionVec_12 <= io_enq_bits_exceptionVec_12; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__2_brIdx <= 4'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h2 == value) begin // @[FlushableQueue.scala 46:24]
        REG__2_brIdx <= io_enq_bits_brIdx; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__3_instr <= 64'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h3 == value) begin // @[FlushableQueue.scala 46:24]
        REG__3_instr <= io_enq_bits_instr; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__3_pc <= 39'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h3 == value) begin // @[FlushableQueue.scala 46:24]
        REG__3_pc <= io_enq_bits_pc; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__3_pnpc <= 39'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h3 == value) begin // @[FlushableQueue.scala 46:24]
        REG__3_pnpc <= io_enq_bits_pnpc; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__3_exceptionVec_12 <= 1'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h3 == value) begin // @[FlushableQueue.scala 46:24]
        REG__3_exceptionVec_12 <= io_enq_bits_exceptionVec_12; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[FlushableQueue.scala 34:28]
      REG__3_brIdx <= 4'h0; // @[FlushableQueue.scala 34:28]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      if (2'h3 == value) begin // @[FlushableQueue.scala 46:24]
        REG__3_brIdx <= io_enq_bits_brIdx; // @[FlushableQueue.scala 46:24]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 2'h0; // @[Counter.scala 60:40]
    end else if (io_flush) begin // @[FlushableQueue.scala 73:19]
      value <= 2'h0; // @[FlushableQueue.scala 75:21]
    end else if (_T_4) begin // @[FlushableQueue.scala 45:17]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 2'h0; // @[Counter.scala 60:40]
    end else if (io_flush) begin // @[FlushableQueue.scala 73:19]
      value_1 <= 2'h0; // @[FlushableQueue.scala 76:21]
    end else if (_T_5) begin // @[FlushableQueue.scala 49:17]
      value_1 <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[FlushableQueue.scala 37:35]
      REG_1 <= 1'h0; // @[FlushableQueue.scala 37:35]
    end else if (io_flush) begin // @[FlushableQueue.scala 73:19]
      REG_1 <= 1'h0; // @[FlushableQueue.scala 78:16]
    end else if (_T_4 != _T_5) begin // @[FlushableQueue.scala 52:28]
      REG_1 <= _T_4; // @[FlushableQueue.scala 53:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  REG__0_instr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  REG__0_pc = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  REG__0_pnpc = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  REG__0_exceptionVec_12 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG__0_brIdx = _RAND_4[3:0];
  _RAND_5 = {2{`RANDOM}};
  REG__1_instr = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  REG__1_pc = _RAND_6[38:0];
  _RAND_7 = {2{`RANDOM}};
  REG__1_pnpc = _RAND_7[38:0];
  _RAND_8 = {1{`RANDOM}};
  REG__1_exceptionVec_12 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  REG__1_brIdx = _RAND_9[3:0];
  _RAND_10 = {2{`RANDOM}};
  REG__2_instr = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  REG__2_pc = _RAND_11[38:0];
  _RAND_12 = {2{`RANDOM}};
  REG__2_pnpc = _RAND_12[38:0];
  _RAND_13 = {1{`RANDOM}};
  REG__2_exceptionVec_12 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  REG__2_brIdx = _RAND_14[3:0];
  _RAND_15 = {2{`RANDOM}};
  REG__3_instr = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  REG__3_pc = _RAND_16[38:0];
  _RAND_17 = {2{`RANDOM}};
  REG__3_pnpc = _RAND_17[38:0];
  _RAND_18 = {1{`RANDOM}};
  REG__3_exceptionVec_12 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  REG__3_brIdx = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  value = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  value_1 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  REG_1 = _RAND_22[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_Frontend_inorder(
  input         clock,
  input         reset,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [63:0] io_out_0_bits_cf_instr,
  output [38:0] io_out_0_bits_cf_pc,
  output [38:0] io_out_0_bits_cf_pnpc,
  output        io_out_0_bits_cf_exceptionVec_1,
  output        io_out_0_bits_cf_exceptionVec_2,
  output        io_out_0_bits_cf_exceptionVec_12,
  output        io_out_0_bits_cf_intrVec_0,
  output        io_out_0_bits_cf_intrVec_1,
  output        io_out_0_bits_cf_intrVec_2,
  output        io_out_0_bits_cf_intrVec_3,
  output        io_out_0_bits_cf_intrVec_4,
  output        io_out_0_bits_cf_intrVec_5,
  output        io_out_0_bits_cf_intrVec_6,
  output        io_out_0_bits_cf_intrVec_7,
  output        io_out_0_bits_cf_intrVec_8,
  output        io_out_0_bits_cf_intrVec_9,
  output        io_out_0_bits_cf_intrVec_10,
  output        io_out_0_bits_cf_intrVec_11,
  output [3:0]  io_out_0_bits_cf_brIdx,
  output        io_out_0_bits_cf_crossPageIPFFix,
  output        io_out_0_bits_ctrl_src1Type,
  output        io_out_0_bits_ctrl_src2Type,
  output [2:0]  io_out_0_bits_ctrl_fuType,
  output [6:0]  io_out_0_bits_ctrl_fuOpType,
  output [4:0]  io_out_0_bits_ctrl_rfSrc1,
  output [4:0]  io_out_0_bits_ctrl_rfSrc2,
  output        io_out_0_bits_ctrl_rfWen,
  output [4:0]  io_out_0_bits_ctrl_rfDest,
  output [63:0] io_out_0_bits_data_imm,
  input         io_out_1_ready,
  output        io_out_1_valid,
  output [63:0] io_out_1_bits_cf_instr,
  output [38:0] io_out_1_bits_cf_pc,
  output [38:0] io_out_1_bits_cf_pnpc,
  output        io_out_1_bits_cf_exceptionVec_1,
  output        io_out_1_bits_cf_exceptionVec_2,
  output        io_out_1_bits_cf_exceptionVec_12,
  output        io_out_1_bits_cf_intrVec_0,
  output        io_out_1_bits_cf_intrVec_1,
  output        io_out_1_bits_cf_intrVec_2,
  output        io_out_1_bits_cf_intrVec_3,
  output        io_out_1_bits_cf_intrVec_4,
  output        io_out_1_bits_cf_intrVec_5,
  output        io_out_1_bits_cf_intrVec_6,
  output        io_out_1_bits_cf_intrVec_7,
  output        io_out_1_bits_cf_intrVec_8,
  output        io_out_1_bits_cf_intrVec_9,
  output        io_out_1_bits_cf_intrVec_10,
  output        io_out_1_bits_cf_intrVec_11,
  output [3:0]  io_out_1_bits_cf_brIdx,
  output        io_out_1_bits_cf_crossPageIPFFix,
  output        io_out_1_bits_ctrl_src1Type,
  output        io_out_1_bits_ctrl_src2Type,
  output [2:0]  io_out_1_bits_ctrl_fuType,
  output [6:0]  io_out_1_bits_ctrl_fuOpType,
  output [4:0]  io_out_1_bits_ctrl_rfSrc1,
  output [4:0]  io_out_1_bits_ctrl_rfSrc2,
  output        io_out_1_bits_ctrl_rfWen,
  output [4:0]  io_out_1_bits_ctrl_rfDest,
  output [63:0] io_out_1_bits_data_imm,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [38:0] io_imem_req_bits_addr,
  output [86:0] io_imem_req_bits_user,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input  [86:0] io_imem_resp_bits_user,
  output [3:0]  io_flushVec,
  input         io_ipf,
  input  [38:0] io_redirect_target,
  input         io_redirect_valid,
  input         flushICache,
  input         REG_6_valid,
  input  [38:0] REG_6_pc,
  input         REG_6_isMissPredict,
  input  [38:0] REG_6_actualTarget,
  input         REG_6_actualTaken,
  input  [6:0]  REG_6_fuOpType,
  input  [1:0]  REG_6_btbType,
  input         REG_6_isRVC,
  input         vmEnable,
  input  [11:0] intrVec,
  input         flushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_clock; // @[Frontend.scala 106:20]
  wire  ifu_reset; // @[Frontend.scala 106:20]
  wire  ifu_io_imem_req_ready; // @[Frontend.scala 106:20]
  wire  ifu_io_imem_req_valid; // @[Frontend.scala 106:20]
  wire [38:0] ifu_io_imem_req_bits_addr; // @[Frontend.scala 106:20]
  wire [81:0] ifu_io_imem_req_bits_user; // @[Frontend.scala 106:20]
  wire  ifu_io_imem_resp_ready; // @[Frontend.scala 106:20]
  wire  ifu_io_imem_resp_valid; // @[Frontend.scala 106:20]
  wire [63:0] ifu_io_imem_resp_bits_rdata; // @[Frontend.scala 106:20]
  wire [81:0] ifu_io_imem_resp_bits_user; // @[Frontend.scala 106:20]
  wire  ifu_io_out_ready; // @[Frontend.scala 106:20]
  wire  ifu_io_out_valid; // @[Frontend.scala 106:20]
  wire [63:0] ifu_io_out_bits_instr; // @[Frontend.scala 106:20]
  wire [38:0] ifu_io_out_bits_pc; // @[Frontend.scala 106:20]
  wire [38:0] ifu_io_out_bits_pnpc; // @[Frontend.scala 106:20]
  wire  ifu_io_out_bits_exceptionVec_12; // @[Frontend.scala 106:20]
  wire [3:0] ifu_io_out_bits_brIdx; // @[Frontend.scala 106:20]
  wire [38:0] ifu_io_redirect_target; // @[Frontend.scala 106:20]
  wire  ifu_io_redirect_valid; // @[Frontend.scala 106:20]
  wire [3:0] ifu_io_flushVec; // @[Frontend.scala 106:20]
  wire  ifu_io_ipf; // @[Frontend.scala 106:20]
  wire  ifu_flushICache; // @[Frontend.scala 106:20]
  wire  ifu_REG_6_valid; // @[Frontend.scala 106:20]
  wire [38:0] ifu_REG_6_pc; // @[Frontend.scala 106:20]
  wire  ifu_REG_6_isMissPredict; // @[Frontend.scala 106:20]
  wire [38:0] ifu_REG_6_actualTarget; // @[Frontend.scala 106:20]
  wire  ifu_REG_6_actualTaken; // @[Frontend.scala 106:20]
  wire [6:0] ifu_REG_6_fuOpType; // @[Frontend.scala 106:20]
  wire [1:0] ifu_REG_6_btbType; // @[Frontend.scala 106:20]
  wire  ifu_REG_6_isRVC; // @[Frontend.scala 106:20]
  wire  ifu_flushTLB; // @[Frontend.scala 106:20]
  wire  ibf_clock; // @[Frontend.scala 107:19]
  wire  ibf_reset; // @[Frontend.scala 107:19]
  wire  ibf_io_in_ready; // @[Frontend.scala 107:19]
  wire  ibf_io_in_valid; // @[Frontend.scala 107:19]
  wire [63:0] ibf_io_in_bits_instr; // @[Frontend.scala 107:19]
  wire [38:0] ibf_io_in_bits_pc; // @[Frontend.scala 107:19]
  wire [38:0] ibf_io_in_bits_pnpc; // @[Frontend.scala 107:19]
  wire  ibf_io_in_bits_exceptionVec_12; // @[Frontend.scala 107:19]
  wire [3:0] ibf_io_in_bits_brIdx; // @[Frontend.scala 107:19]
  wire  ibf_io_out_ready; // @[Frontend.scala 107:19]
  wire  ibf_io_out_valid; // @[Frontend.scala 107:19]
  wire [63:0] ibf_io_out_bits_instr; // @[Frontend.scala 107:19]
  wire [38:0] ibf_io_out_bits_pc; // @[Frontend.scala 107:19]
  wire [38:0] ibf_io_out_bits_pnpc; // @[Frontend.scala 107:19]
  wire  ibf_io_out_bits_exceptionVec_12; // @[Frontend.scala 107:19]
  wire [3:0] ibf_io_out_bits_brIdx; // @[Frontend.scala 107:19]
  wire  ibf_io_out_bits_crossPageIPFFix; // @[Frontend.scala 107:19]
  wire  ibf_io_flush; // @[Frontend.scala 107:19]
  wire  idu_io_in_0_ready; // @[Frontend.scala 108:20]
  wire  idu_io_in_0_valid; // @[Frontend.scala 108:20]
  wire [63:0] idu_io_in_0_bits_instr; // @[Frontend.scala 108:20]
  wire [38:0] idu_io_in_0_bits_pc; // @[Frontend.scala 108:20]
  wire [38:0] idu_io_in_0_bits_pnpc; // @[Frontend.scala 108:20]
  wire  idu_io_in_0_bits_exceptionVec_12; // @[Frontend.scala 108:20]
  wire [3:0] idu_io_in_0_bits_brIdx; // @[Frontend.scala 108:20]
  wire  idu_io_in_0_bits_crossPageIPFFix; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_ready; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_valid; // @[Frontend.scala 108:20]
  wire [63:0] idu_io_out_0_bits_cf_instr; // @[Frontend.scala 108:20]
  wire [38:0] idu_io_out_0_bits_cf_pc; // @[Frontend.scala 108:20]
  wire [38:0] idu_io_out_0_bits_cf_pnpc; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_1; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_2; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_12; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_0; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_1; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_2; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_3; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_4; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_5; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_6; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_7; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_8; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_9; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_10; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_11; // @[Frontend.scala 108:20]
  wire [3:0] idu_io_out_0_bits_cf_brIdx; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_crossPageIPFFix; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_ctrl_src1Type; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_ctrl_src2Type; // @[Frontend.scala 108:20]
  wire [2:0] idu_io_out_0_bits_ctrl_fuType; // @[Frontend.scala 108:20]
  wire [6:0] idu_io_out_0_bits_ctrl_fuOpType; // @[Frontend.scala 108:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc1; // @[Frontend.scala 108:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc2; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_ctrl_rfWen; // @[Frontend.scala 108:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfDest; // @[Frontend.scala 108:20]
  wire [63:0] idu_io_out_0_bits_data_imm; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_ready; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_valid; // @[Frontend.scala 108:20]
  wire [63:0] idu_io_out_1_bits_cf_instr; // @[Frontend.scala 108:20]
  wire [38:0] idu_io_out_1_bits_cf_pc; // @[Frontend.scala 108:20]
  wire [38:0] idu_io_out_1_bits_cf_pnpc; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_exceptionVec_1; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_exceptionVec_2; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_exceptionVec_12; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_0; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_1; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_2; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_3; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_4; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_5; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_6; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_7; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_8; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_9; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_10; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_11; // @[Frontend.scala 108:20]
  wire [3:0] idu_io_out_1_bits_cf_brIdx; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_crossPageIPFFix; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_ctrl_src1Type; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_ctrl_src2Type; // @[Frontend.scala 108:20]
  wire [2:0] idu_io_out_1_bits_ctrl_fuType; // @[Frontend.scala 108:20]
  wire [6:0] idu_io_out_1_bits_ctrl_fuOpType; // @[Frontend.scala 108:20]
  wire [4:0] idu_io_out_1_bits_ctrl_rfSrc1; // @[Frontend.scala 108:20]
  wire [4:0] idu_io_out_1_bits_ctrl_rfSrc2; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_ctrl_rfWen; // @[Frontend.scala 108:20]
  wire [4:0] idu_io_out_1_bits_ctrl_rfDest; // @[Frontend.scala 108:20]
  wire [63:0] idu_io_out_1_bits_data_imm; // @[Frontend.scala 108:20]
  wire  idu_vmEnable; // @[Frontend.scala 108:20]
  wire [11:0] idu_intrVec; // @[Frontend.scala 108:20]
  wire  FlushableQueue_clock; // @[FlushableQueue.scala 105:21]
  wire  FlushableQueue_reset; // @[FlushableQueue.scala 105:21]
  wire  FlushableQueue_io_enq_ready; // @[FlushableQueue.scala 105:21]
  wire  FlushableQueue_io_enq_valid; // @[FlushableQueue.scala 105:21]
  wire [63:0] FlushableQueue_io_enq_bits_instr; // @[FlushableQueue.scala 105:21]
  wire [38:0] FlushableQueue_io_enq_bits_pc; // @[FlushableQueue.scala 105:21]
  wire [38:0] FlushableQueue_io_enq_bits_pnpc; // @[FlushableQueue.scala 105:21]
  wire  FlushableQueue_io_enq_bits_exceptionVec_12; // @[FlushableQueue.scala 105:21]
  wire [3:0] FlushableQueue_io_enq_bits_brIdx; // @[FlushableQueue.scala 105:21]
  wire  FlushableQueue_io_deq_ready; // @[FlushableQueue.scala 105:21]
  wire  FlushableQueue_io_deq_valid; // @[FlushableQueue.scala 105:21]
  wire [63:0] FlushableQueue_io_deq_bits_instr; // @[FlushableQueue.scala 105:21]
  wire [38:0] FlushableQueue_io_deq_bits_pc; // @[FlushableQueue.scala 105:21]
  wire [38:0] FlushableQueue_io_deq_bits_pnpc; // @[FlushableQueue.scala 105:21]
  wire  FlushableQueue_io_deq_bits_exceptionVec_12; // @[FlushableQueue.scala 105:21]
  wire [3:0] FlushableQueue_io_deq_bits_brIdx; // @[FlushableQueue.scala 105:21]
  wire  FlushableQueue_io_flush; // @[FlushableQueue.scala 105:21]
  wire  _T_1 = idu_io_out_0_ready & idu_io_out_0_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T_1 ? 1'h0 : REG; // @[Pipeline.scala 25:25 Pipeline.scala 25:33 Pipeline.scala 24:24]
  wire  _T_3 = ibf_io_out_valid & idu_io_in_0_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = ibf_io_out_valid & idu_io_in_0_ready | _GEN_0; // @[Pipeline.scala 26:38 Pipeline.scala 26:46]
  reg [63:0] REG_1_instr; // @[Reg.scala 27:20]
  reg [38:0] REG_1_pc; // @[Reg.scala 27:20]
  reg [38:0] REG_1_pnpc; // @[Reg.scala 27:20]
  reg  REG_1_exceptionVec_12; // @[Reg.scala 27:20]
  reg [3:0] REG_1_brIdx; // @[Reg.scala 27:20]
  reg  REG_1_crossPageIPFFix; // @[Reg.scala 27:20]
  ysyx_210000_IFU_inorder ifu ( // @[Frontend.scala 106:20]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_imem_req_ready(ifu_io_imem_req_ready),
    .io_imem_req_valid(ifu_io_imem_req_valid),
    .io_imem_req_bits_addr(ifu_io_imem_req_bits_addr),
    .io_imem_req_bits_user(ifu_io_imem_req_bits_user),
    .io_imem_resp_ready(ifu_io_imem_resp_ready),
    .io_imem_resp_valid(ifu_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(ifu_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(ifu_io_imem_resp_bits_user),
    .io_out_ready(ifu_io_out_ready),
    .io_out_valid(ifu_io_out_valid),
    .io_out_bits_instr(ifu_io_out_bits_instr),
    .io_out_bits_pc(ifu_io_out_bits_pc),
    .io_out_bits_pnpc(ifu_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_12(ifu_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ifu_io_out_bits_brIdx),
    .io_redirect_target(ifu_io_redirect_target),
    .io_redirect_valid(ifu_io_redirect_valid),
    .io_flushVec(ifu_io_flushVec),
    .io_ipf(ifu_io_ipf),
    .flushICache(ifu_flushICache),
    .REG_6_valid(ifu_REG_6_valid),
    .REG_6_pc(ifu_REG_6_pc),
    .REG_6_isMissPredict(ifu_REG_6_isMissPredict),
    .REG_6_actualTarget(ifu_REG_6_actualTarget),
    .REG_6_actualTaken(ifu_REG_6_actualTaken),
    .REG_6_fuOpType(ifu_REG_6_fuOpType),
    .REG_6_btbType(ifu_REG_6_btbType),
    .REG_6_isRVC(ifu_REG_6_isRVC),
    .flushTLB(ifu_flushTLB)
  );
  ysyx_210000_NaiveRVCAlignBuffer ibf ( // @[Frontend.scala 107:19]
    .clock(ibf_clock),
    .reset(ibf_reset),
    .io_in_ready(ibf_io_in_ready),
    .io_in_valid(ibf_io_in_valid),
    .io_in_bits_instr(ibf_io_in_bits_instr),
    .io_in_bits_pc(ibf_io_in_bits_pc),
    .io_in_bits_pnpc(ibf_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_12(ibf_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(ibf_io_in_bits_brIdx),
    .io_out_ready(ibf_io_out_ready),
    .io_out_valid(ibf_io_out_valid),
    .io_out_bits_instr(ibf_io_out_bits_instr),
    .io_out_bits_pc(ibf_io_out_bits_pc),
    .io_out_bits_pnpc(ibf_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_12(ibf_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ibf_io_out_bits_brIdx),
    .io_out_bits_crossPageIPFFix(ibf_io_out_bits_crossPageIPFFix),
    .io_flush(ibf_io_flush)
  );
  ysyx_210000_IDU idu ( // @[Frontend.scala 108:20]
    .io_in_0_ready(idu_io_in_0_ready),
    .io_in_0_valid(idu_io_in_0_valid),
    .io_in_0_bits_instr(idu_io_in_0_bits_instr),
    .io_in_0_bits_pc(idu_io_in_0_bits_pc),
    .io_in_0_bits_pnpc(idu_io_in_0_bits_pnpc),
    .io_in_0_bits_exceptionVec_12(idu_io_in_0_bits_exceptionVec_12),
    .io_in_0_bits_brIdx(idu_io_in_0_bits_brIdx),
    .io_in_0_bits_crossPageIPFFix(idu_io_in_0_bits_crossPageIPFFix),
    .io_out_0_ready(idu_io_out_0_ready),
    .io_out_0_valid(idu_io_out_0_valid),
    .io_out_0_bits_cf_instr(idu_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(idu_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(idu_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(idu_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(idu_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(idu_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_0(idu_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(idu_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(idu_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(idu_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(idu_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(idu_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(idu_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(idu_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(idu_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(idu_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(idu_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(idu_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(idu_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossPageIPFFix(idu_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_ctrl_src1Type(idu_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(idu_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(idu_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(idu_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(idu_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(idu_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(idu_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(idu_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_data_imm(idu_io_out_0_bits_data_imm),
    .io_out_1_ready(idu_io_out_1_ready),
    .io_out_1_valid(idu_io_out_1_valid),
    .io_out_1_bits_cf_instr(idu_io_out_1_bits_cf_instr),
    .io_out_1_bits_cf_pc(idu_io_out_1_bits_cf_pc),
    .io_out_1_bits_cf_pnpc(idu_io_out_1_bits_cf_pnpc),
    .io_out_1_bits_cf_exceptionVec_1(idu_io_out_1_bits_cf_exceptionVec_1),
    .io_out_1_bits_cf_exceptionVec_2(idu_io_out_1_bits_cf_exceptionVec_2),
    .io_out_1_bits_cf_exceptionVec_12(idu_io_out_1_bits_cf_exceptionVec_12),
    .io_out_1_bits_cf_intrVec_0(idu_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(idu_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(idu_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(idu_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(idu_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(idu_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(idu_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(idu_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(idu_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(idu_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(idu_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(idu_io_out_1_bits_cf_intrVec_11),
    .io_out_1_bits_cf_brIdx(idu_io_out_1_bits_cf_brIdx),
    .io_out_1_bits_cf_crossPageIPFFix(idu_io_out_1_bits_cf_crossPageIPFFix),
    .io_out_1_bits_ctrl_src1Type(idu_io_out_1_bits_ctrl_src1Type),
    .io_out_1_bits_ctrl_src2Type(idu_io_out_1_bits_ctrl_src2Type),
    .io_out_1_bits_ctrl_fuType(idu_io_out_1_bits_ctrl_fuType),
    .io_out_1_bits_ctrl_fuOpType(idu_io_out_1_bits_ctrl_fuOpType),
    .io_out_1_bits_ctrl_rfSrc1(idu_io_out_1_bits_ctrl_rfSrc1),
    .io_out_1_bits_ctrl_rfSrc2(idu_io_out_1_bits_ctrl_rfSrc2),
    .io_out_1_bits_ctrl_rfWen(idu_io_out_1_bits_ctrl_rfWen),
    .io_out_1_bits_ctrl_rfDest(idu_io_out_1_bits_ctrl_rfDest),
    .io_out_1_bits_data_imm(idu_io_out_1_bits_data_imm),
    .vmEnable(idu_vmEnable),
    .intrVec(idu_intrVec)
  );
  ysyx_210000_FlushableQueue FlushableQueue ( // @[FlushableQueue.scala 105:21]
    .clock(FlushableQueue_clock),
    .reset(FlushableQueue_reset),
    .io_enq_ready(FlushableQueue_io_enq_ready),
    .io_enq_valid(FlushableQueue_io_enq_valid),
    .io_enq_bits_instr(FlushableQueue_io_enq_bits_instr),
    .io_enq_bits_pc(FlushableQueue_io_enq_bits_pc),
    .io_enq_bits_pnpc(FlushableQueue_io_enq_bits_pnpc),
    .io_enq_bits_exceptionVec_12(FlushableQueue_io_enq_bits_exceptionVec_12),
    .io_enq_bits_brIdx(FlushableQueue_io_enq_bits_brIdx),
    .io_deq_ready(FlushableQueue_io_deq_ready),
    .io_deq_valid(FlushableQueue_io_deq_valid),
    .io_deq_bits_instr(FlushableQueue_io_deq_bits_instr),
    .io_deq_bits_pc(FlushableQueue_io_deq_bits_pc),
    .io_deq_bits_pnpc(FlushableQueue_io_deq_bits_pnpc),
    .io_deq_bits_exceptionVec_12(FlushableQueue_io_deq_bits_exceptionVec_12),
    .io_deq_bits_brIdx(FlushableQueue_io_deq_bits_brIdx),
    .io_flush(FlushableQueue_io_flush)
  );
  assign io_out_0_valid = idu_io_out_0_valid; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_instr = idu_io_out_0_bits_cf_instr; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_pc = idu_io_out_0_bits_cf_pc; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_pnpc = idu_io_out_0_bits_cf_pnpc; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_exceptionVec_1 = idu_io_out_0_bits_cf_exceptionVec_1; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_exceptionVec_2 = idu_io_out_0_bits_cf_exceptionVec_2; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_exceptionVec_12 = idu_io_out_0_bits_cf_exceptionVec_12; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_0 = idu_io_out_0_bits_cf_intrVec_0; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_1 = idu_io_out_0_bits_cf_intrVec_1; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_2 = idu_io_out_0_bits_cf_intrVec_2; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_3 = idu_io_out_0_bits_cf_intrVec_3; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_4 = idu_io_out_0_bits_cf_intrVec_4; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_5 = idu_io_out_0_bits_cf_intrVec_5; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_6 = idu_io_out_0_bits_cf_intrVec_6; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_7 = idu_io_out_0_bits_cf_intrVec_7; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_8 = idu_io_out_0_bits_cf_intrVec_8; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_9 = idu_io_out_0_bits_cf_intrVec_9; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_10 = idu_io_out_0_bits_cf_intrVec_10; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_11 = idu_io_out_0_bits_cf_intrVec_11; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_brIdx = idu_io_out_0_bits_cf_brIdx; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_crossPageIPFFix = idu_io_out_0_bits_cf_crossPageIPFFix; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_src1Type = idu_io_out_0_bits_ctrl_src1Type; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_src2Type = idu_io_out_0_bits_ctrl_src2Type; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_fuType = idu_io_out_0_bits_ctrl_fuType; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_fuOpType = idu_io_out_0_bits_ctrl_fuOpType; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_rfSrc1 = idu_io_out_0_bits_ctrl_rfSrc1; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_rfSrc2 = idu_io_out_0_bits_ctrl_rfSrc2; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_rfWen = idu_io_out_0_bits_ctrl_rfWen; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_rfDest = idu_io_out_0_bits_ctrl_rfDest; // @[Frontend.scala 120:10]
  assign io_out_0_bits_data_imm = idu_io_out_0_bits_data_imm; // @[Frontend.scala 120:10]
  assign io_out_1_valid = idu_io_out_1_valid; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_instr = idu_io_out_1_bits_cf_instr; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_pc = idu_io_out_1_bits_cf_pc; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_pnpc = idu_io_out_1_bits_cf_pnpc; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_exceptionVec_1 = idu_io_out_1_bits_cf_exceptionVec_1; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_exceptionVec_2 = idu_io_out_1_bits_cf_exceptionVec_2; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_exceptionVec_12 = idu_io_out_1_bits_cf_exceptionVec_12; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_0 = idu_io_out_1_bits_cf_intrVec_0; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_1 = idu_io_out_1_bits_cf_intrVec_1; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_2 = idu_io_out_1_bits_cf_intrVec_2; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_3 = idu_io_out_1_bits_cf_intrVec_3; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_4 = idu_io_out_1_bits_cf_intrVec_4; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_5 = idu_io_out_1_bits_cf_intrVec_5; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_6 = idu_io_out_1_bits_cf_intrVec_6; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_7 = idu_io_out_1_bits_cf_intrVec_7; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_8 = idu_io_out_1_bits_cf_intrVec_8; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_9 = idu_io_out_1_bits_cf_intrVec_9; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_10 = idu_io_out_1_bits_cf_intrVec_10; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_11 = idu_io_out_1_bits_cf_intrVec_11; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_brIdx = idu_io_out_1_bits_cf_brIdx; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_crossPageIPFFix = idu_io_out_1_bits_cf_crossPageIPFFix; // @[Frontend.scala 120:10]
  assign io_out_1_bits_ctrl_src1Type = idu_io_out_1_bits_ctrl_src1Type; // @[Frontend.scala 120:10]
  assign io_out_1_bits_ctrl_src2Type = idu_io_out_1_bits_ctrl_src2Type; // @[Frontend.scala 120:10]
  assign io_out_1_bits_ctrl_fuType = idu_io_out_1_bits_ctrl_fuType; // @[Frontend.scala 120:10]
  assign io_out_1_bits_ctrl_fuOpType = idu_io_out_1_bits_ctrl_fuOpType; // @[Frontend.scala 120:10]
  assign io_out_1_bits_ctrl_rfSrc1 = idu_io_out_1_bits_ctrl_rfSrc1; // @[Frontend.scala 120:10]
  assign io_out_1_bits_ctrl_rfSrc2 = idu_io_out_1_bits_ctrl_rfSrc2; // @[Frontend.scala 120:10]
  assign io_out_1_bits_ctrl_rfWen = idu_io_out_1_bits_ctrl_rfWen; // @[Frontend.scala 120:10]
  assign io_out_1_bits_ctrl_rfDest = idu_io_out_1_bits_ctrl_rfDest; // @[Frontend.scala 120:10]
  assign io_out_1_bits_data_imm = idu_io_out_1_bits_data_imm; // @[Frontend.scala 120:10]
  assign io_imem_req_valid = ifu_io_imem_req_valid; // @[Frontend.scala 125:11]
  assign io_imem_req_bits_addr = ifu_io_imem_req_bits_addr; // @[Frontend.scala 125:11]
  assign io_imem_req_bits_user = {{5'd0}, ifu_io_imem_req_bits_user}; // @[Frontend.scala 125:11]
  assign io_imem_resp_ready = ifu_io_imem_resp_ready; // @[Frontend.scala 125:11]
  assign io_flushVec = ifu_io_flushVec; // @[Frontend.scala 122:15]
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_imem_req_ready = io_imem_req_ready; // @[Frontend.scala 125:11]
  assign ifu_io_imem_resp_valid = io_imem_resp_valid; // @[Frontend.scala 125:11]
  assign ifu_io_imem_resp_bits_rdata = io_imem_resp_bits_rdata; // @[Frontend.scala 125:11]
  assign ifu_io_imem_resp_bits_user = io_imem_resp_bits_user[81:0]; // @[Frontend.scala 125:11]
  assign ifu_io_out_ready = FlushableQueue_io_enq_ready; // @[FlushableQueue.scala 109:17]
  assign ifu_io_redirect_target = io_redirect_target; // @[Frontend.scala 121:15]
  assign ifu_io_redirect_valid = io_redirect_valid; // @[Frontend.scala 121:15]
  assign ifu_io_ipf = io_ipf; // @[Frontend.scala 124:10]
  assign ifu_flushICache = flushICache;
  assign ifu_REG_6_valid = REG_6_valid;
  assign ifu_REG_6_pc = REG_6_pc;
  assign ifu_REG_6_isMissPredict = REG_6_isMissPredict;
  assign ifu_REG_6_actualTarget = REG_6_actualTarget;
  assign ifu_REG_6_actualTaken = REG_6_actualTaken;
  assign ifu_REG_6_fuOpType = REG_6_fuOpType;
  assign ifu_REG_6_btbType = REG_6_btbType;
  assign ifu_REG_6_isRVC = REG_6_isRVC;
  assign ifu_flushTLB = flushTLB;
  assign ibf_clock = clock;
  assign ibf_reset = reset;
  assign ibf_io_in_valid = FlushableQueue_io_deq_valid; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_instr = FlushableQueue_io_deq_bits_instr; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_pc = FlushableQueue_io_deq_bits_pc; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_pnpc = FlushableQueue_io_deq_bits_pnpc; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_exceptionVec_12 = FlushableQueue_io_deq_bits_exceptionVec_12; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_brIdx = FlushableQueue_io_deq_bits_brIdx; // @[Frontend.scala 112:11]
  assign ibf_io_out_ready = idu_io_in_0_ready; // @[Pipeline.scala 29:16]
  assign ibf_io_flush = ifu_io_flushVec[1]; // @[Frontend.scala 119:34]
  assign idu_io_in_0_valid = REG; // @[Pipeline.scala 31:17]
  assign idu_io_in_0_bits_instr = REG_1_instr; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pc = REG_1_pc; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pnpc = REG_1_pnpc; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_exceptionVec_12 = REG_1_exceptionVec_12; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_brIdx = REG_1_brIdx; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_crossPageIPFFix = REG_1_crossPageIPFFix; // @[Pipeline.scala 30:16]
  assign idu_io_out_0_ready = io_out_0_ready; // @[Frontend.scala 120:10]
  assign idu_io_out_1_ready = io_out_1_ready; // @[Frontend.scala 120:10]
  assign idu_vmEnable = vmEnable;
  assign idu_intrVec = intrVec;
  assign FlushableQueue_clock = clock;
  assign FlushableQueue_reset = reset;
  assign FlushableQueue_io_enq_valid = ifu_io_out_valid; // @[FlushableQueue.scala 106:22]
  assign FlushableQueue_io_enq_bits_instr = ifu_io_out_bits_instr; // @[FlushableQueue.scala 107:21]
  assign FlushableQueue_io_enq_bits_pc = ifu_io_out_bits_pc; // @[FlushableQueue.scala 107:21]
  assign FlushableQueue_io_enq_bits_pnpc = ifu_io_out_bits_pnpc; // @[FlushableQueue.scala 107:21]
  assign FlushableQueue_io_enq_bits_exceptionVec_12 = ifu_io_out_bits_exceptionVec_12; // @[FlushableQueue.scala 107:21]
  assign FlushableQueue_io_enq_bits_brIdx = ifu_io_out_bits_brIdx; // @[FlushableQueue.scala 107:21]
  assign FlushableQueue_io_deq_ready = ibf_io_in_ready; // @[Frontend.scala 112:11]
  assign FlushableQueue_io_flush = ifu_io_flushVec[0]; // @[Frontend.scala 115:58]
  always @(posedge clock) begin
    if (reset) begin // @[Pipeline.scala 24:24]
      REG <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (ifu_io_flushVec[1]) begin // @[Pipeline.scala 27:20]
      REG <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG <= _GEN_1;
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_instr <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_3) begin // @[Reg.scala 28:19]
      REG_1_instr <= ibf_io_out_bits_instr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_pc <= 39'h0; // @[Reg.scala 27:20]
    end else if (_T_3) begin // @[Reg.scala 28:19]
      REG_1_pc <= ibf_io_out_bits_pc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_pnpc <= 39'h0; // @[Reg.scala 27:20]
    end else if (_T_3) begin // @[Reg.scala 28:19]
      REG_1_pnpc <= ibf_io_out_bits_pnpc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_exceptionVec_12 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_3) begin // @[Reg.scala 28:19]
      REG_1_exceptionVec_12 <= ibf_io_out_bits_exceptionVec_12; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_brIdx <= 4'h0; // @[Reg.scala 27:20]
    end else if (_T_3) begin // @[Reg.scala 28:19]
      REG_1_brIdx <= ibf_io_out_bits_brIdx; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_crossPageIPFFix <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_3) begin // @[Reg.scala 28:19]
      REG_1_crossPageIPFFix <= ibf_io_out_bits_crossPageIPFFix; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  REG_1_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  REG_1_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  REG_1_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  REG_1_exceptionVec_12 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1_brIdx = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  REG_1_crossPageIPFFix = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_ISU(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_cf_instr,
  input  [38:0] io_in_0_bits_cf_pc,
  input  [38:0] io_in_0_bits_cf_pnpc,
  input         io_in_0_bits_cf_exceptionVec_1,
  input         io_in_0_bits_cf_exceptionVec_2,
  input         io_in_0_bits_cf_exceptionVec_12,
  input         io_in_0_bits_cf_intrVec_0,
  input         io_in_0_bits_cf_intrVec_1,
  input         io_in_0_bits_cf_intrVec_2,
  input         io_in_0_bits_cf_intrVec_3,
  input         io_in_0_bits_cf_intrVec_4,
  input         io_in_0_bits_cf_intrVec_5,
  input         io_in_0_bits_cf_intrVec_6,
  input         io_in_0_bits_cf_intrVec_7,
  input         io_in_0_bits_cf_intrVec_8,
  input         io_in_0_bits_cf_intrVec_9,
  input         io_in_0_bits_cf_intrVec_10,
  input         io_in_0_bits_cf_intrVec_11,
  input  [3:0]  io_in_0_bits_cf_brIdx,
  input         io_in_0_bits_cf_crossPageIPFFix,
  input         io_in_0_bits_ctrl_src1Type,
  input         io_in_0_bits_ctrl_src2Type,
  input  [2:0]  io_in_0_bits_ctrl_fuType,
  input  [6:0]  io_in_0_bits_ctrl_fuOpType,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2,
  input         io_in_0_bits_ctrl_rfWen,
  input  [4:0]  io_in_0_bits_ctrl_rfDest,
  input  [63:0] io_in_0_bits_data_imm,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_cf_instr,
  output [38:0] io_out_bits_cf_pc,
  output [38:0] io_out_bits_cf_pnpc,
  output        io_out_bits_cf_exceptionVec_1,
  output        io_out_bits_cf_exceptionVec_2,
  output        io_out_bits_cf_exceptionVec_12,
  output        io_out_bits_cf_intrVec_0,
  output        io_out_bits_cf_intrVec_1,
  output        io_out_bits_cf_intrVec_2,
  output        io_out_bits_cf_intrVec_3,
  output        io_out_bits_cf_intrVec_4,
  output        io_out_bits_cf_intrVec_5,
  output        io_out_bits_cf_intrVec_6,
  output        io_out_bits_cf_intrVec_7,
  output        io_out_bits_cf_intrVec_8,
  output        io_out_bits_cf_intrVec_9,
  output        io_out_bits_cf_intrVec_10,
  output        io_out_bits_cf_intrVec_11,
  output [3:0]  io_out_bits_cf_brIdx,
  output        io_out_bits_cf_crossPageIPFFix,
  output [2:0]  io_out_bits_ctrl_fuType,
  output [6:0]  io_out_bits_ctrl_fuOpType,
  output        io_out_bits_ctrl_rfWen,
  output [4:0]  io_out_bits_ctrl_rfDest,
  output        io_out_bits_ctrl_permitLibLoad,
  output        io_out_bits_ctrl_permitLibStore,
  output        io_out_bits_ctrl_lsuIsLoad,
  output [63:0] io_out_bits_data_src1,
  output [63:0] io_out_bits_data_src2,
  output [63:0] io_out_bits_data_imm,
  output [63:0] io_out_bits_data_addr,
  input         io_wb_rfWen,
  input  [4:0]  io_wb_rfDest,
  input  [63:0] io_wb_rfData,
  input         io_forward_valid,
  input         io_forward_wb_rfWen,
  input  [4:0]  io_forward_wb_rfDest,
  input  [63:0] io_forward_wb_rfData,
  input  [2:0]  io_forward_fuType,
  input         io_flush,
  output [63:0] isuAddr_0,
  input         isu_perm_lib_ld,
  input         isu_perm_lib_st
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  wire  forwardRfWen = io_forward_wb_rfWen & io_forward_valid; // @[ISU.scala 42:42]
  wire  dontForward1 = io_forward_fuType != 3'h0 & io_forward_fuType != 3'h1; // @[ISU.scala 43:57]
  wire  src1DependEX = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_forward_wb_rfDest &
    forwardRfWen; // @[ISU.scala 40:100]
  wire  src2DependEX = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_forward_wb_rfDest &
    forwardRfWen; // @[ISU.scala 40:100]
  wire  src1DependWB = io_in_0_bits_ctrl_rfSrc1 != 5'h0 & io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest & io_wb_rfWen; // @[ISU.scala 40:100]
  wire  src2DependWB = io_in_0_bits_ctrl_rfSrc2 != 5'h0 & io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest & io_wb_rfWen; // @[ISU.scala 40:100]
  wire  _T_14 = ~dontForward1; // @[ISU.scala 49:46]
  wire  src1ForwardNextCycle = src1DependEX & ~dontForward1; // @[ISU.scala 49:43]
  wire  src2ForwardNextCycle = src2DependEX & _T_14; // @[ISU.scala 50:43]
  wire  _T_17 = dontForward1 ? ~src1DependEX : 1'h1; // @[ISU.scala 51:40]
  wire  src1Forward = src1DependWB & _T_17; // @[ISU.scala 51:34]
  wire  _T_19 = dontForward1 ? ~src2DependEX : 1'h1; // @[ISU.scala 52:40]
  wire  src2Forward = src2DependWB & _T_19; // @[ISU.scala 52:34]
  reg [31:0] REG; // @[RF.scala 37:21]
  wire [31:0] _T_20 = REG >> io_in_0_bits_ctrl_rfSrc1; // @[RF.scala 38:37]
  wire  src1Ready = ~_T_20[0] | src1ForwardNextCycle | src1Forward; // @[ISU.scala 55:62]
  wire [31:0] _T_24 = REG >> io_in_0_bits_ctrl_rfSrc2; // @[RF.scala 38:37]
  wire  src2Ready = ~_T_24[0] | src2ForwardNextCycle | src2Forward; // @[ISU.scala 56:62]
  reg [63:0] REG_1_0; // @[RF.scala 31:19]
  reg [63:0] REG_1_1; // @[RF.scala 31:19]
  reg [63:0] REG_1_2; // @[RF.scala 31:19]
  reg [63:0] REG_1_3; // @[RF.scala 31:19]
  reg [63:0] REG_1_4; // @[RF.scala 31:19]
  reg [63:0] REG_1_5; // @[RF.scala 31:19]
  reg [63:0] REG_1_6; // @[RF.scala 31:19]
  reg [63:0] REG_1_7; // @[RF.scala 31:19]
  reg [63:0] REG_1_8; // @[RF.scala 31:19]
  reg [63:0] REG_1_9; // @[RF.scala 31:19]
  reg [63:0] REG_1_10; // @[RF.scala 31:19]
  reg [63:0] REG_1_11; // @[RF.scala 31:19]
  reg [63:0] REG_1_12; // @[RF.scala 31:19]
  reg [63:0] REG_1_13; // @[RF.scala 31:19]
  reg [63:0] REG_1_14; // @[RF.scala 31:19]
  reg [63:0] REG_1_15; // @[RF.scala 31:19]
  reg [63:0] REG_1_16; // @[RF.scala 31:19]
  reg [63:0] REG_1_17; // @[RF.scala 31:19]
  reg [63:0] REG_1_18; // @[RF.scala 31:19]
  reg [63:0] REG_1_19; // @[RF.scala 31:19]
  reg [63:0] REG_1_20; // @[RF.scala 31:19]
  reg [63:0] REG_1_21; // @[RF.scala 31:19]
  reg [63:0] REG_1_22; // @[RF.scala 31:19]
  reg [63:0] REG_1_23; // @[RF.scala 31:19]
  reg [63:0] REG_1_24; // @[RF.scala 31:19]
  reg [63:0] REG_1_25; // @[RF.scala 31:19]
  reg [63:0] REG_1_26; // @[RF.scala 31:19]
  reg [63:0] REG_1_27; // @[RF.scala 31:19]
  reg [63:0] REG_1_28; // @[RF.scala 31:19]
  reg [63:0] REG_1_29; // @[RF.scala 31:19]
  reg [63:0] REG_1_30; // @[RF.scala 31:19]
  reg [63:0] REG_1_31; // @[RF.scala 31:19]
  wire [24:0] hi = io_in_0_bits_cf_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_33 = {hi,io_in_0_bits_cf_pc}; // @[Cat.scala 30:58]
  wire  _T_34 = ~src1ForwardNextCycle; // @[ISU.scala 65:21]
  wire  _T_35 = src1Forward & ~src1ForwardNextCycle; // @[ISU.scala 65:18]
  wire  _T_40 = ~io_in_0_bits_ctrl_src1Type & _T_34 & ~src1Forward; // @[ISU.scala 66:76]
  wire [63:0] _GEN_1 = 5'h1 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_1 : REG_1_0; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_2 = 5'h2 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_2 : _GEN_1; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_3 = 5'h3 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_3 : _GEN_2; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_4 = 5'h4 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_4 : _GEN_3; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_5 = 5'h5 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_5 : _GEN_4; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_6 = 5'h6 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_6 : _GEN_5; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_7 = 5'h7 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_7 : _GEN_6; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_8 = 5'h8 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_8 : _GEN_7; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_9 = 5'h9 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_9 : _GEN_8; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_10 = 5'ha == io_in_0_bits_ctrl_rfSrc1 ? REG_1_10 : _GEN_9; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_11 = 5'hb == io_in_0_bits_ctrl_rfSrc1 ? REG_1_11 : _GEN_10; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_12 = 5'hc == io_in_0_bits_ctrl_rfSrc1 ? REG_1_12 : _GEN_11; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_13 = 5'hd == io_in_0_bits_ctrl_rfSrc1 ? REG_1_13 : _GEN_12; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_14 = 5'he == io_in_0_bits_ctrl_rfSrc1 ? REG_1_14 : _GEN_13; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_15 = 5'hf == io_in_0_bits_ctrl_rfSrc1 ? REG_1_15 : _GEN_14; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_16 = 5'h10 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_16 : _GEN_15; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_17 = 5'h11 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_17 : _GEN_16; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_18 = 5'h12 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_18 : _GEN_17; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_19 = 5'h13 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_19 : _GEN_18; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_20 = 5'h14 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_20 : _GEN_19; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_21 = 5'h15 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_21 : _GEN_20; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_22 = 5'h16 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_22 : _GEN_21; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_23 = 5'h17 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_23 : _GEN_22; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_24 = 5'h18 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_24 : _GEN_23; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_25 = 5'h19 == io_in_0_bits_ctrl_rfSrc1 ? REG_1_25 : _GEN_24; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_26 = 5'h1a == io_in_0_bits_ctrl_rfSrc1 ? REG_1_26 : _GEN_25; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_27 = 5'h1b == io_in_0_bits_ctrl_rfSrc1 ? REG_1_27 : _GEN_26; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_28 = 5'h1c == io_in_0_bits_ctrl_rfSrc1 ? REG_1_28 : _GEN_27; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_29 = 5'h1d == io_in_0_bits_ctrl_rfSrc1 ? REG_1_29 : _GEN_28; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_30 = 5'h1e == io_in_0_bits_ctrl_rfSrc1 ? REG_1_30 : _GEN_29; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_31 = 5'h1f == io_in_0_bits_ctrl_rfSrc1 ? REG_1_31 : _GEN_30; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _T_42 = io_in_0_bits_ctrl_rfSrc1 == 5'h0 ? 64'h0 : _GEN_31; // @[RF.scala 32:36]
  wire [63:0] _T_43 = io_in_0_bits_ctrl_src1Type ? _T_33 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_44 = src1ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = _T_35 ? io_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = _T_40 ? _T_42 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_47 = _T_43 | _T_44; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = _T_47 | _T_45; // @[Mux.scala 27:72]
  wire  _T_51 = ~src2ForwardNextCycle; // @[ISU.scala 71:21]
  wire  _T_52 = src2Forward & ~src2ForwardNextCycle; // @[ISU.scala 71:18]
  wire  _T_57 = ~io_in_0_bits_ctrl_src2Type & _T_51 & ~src2Forward; // @[ISU.scala 72:77]
  wire [63:0] _GEN_33 = 5'h1 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_1 : REG_1_0; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_34 = 5'h2 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_2 : _GEN_33; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_35 = 5'h3 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_3 : _GEN_34; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_36 = 5'h4 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_4 : _GEN_35; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_37 = 5'h5 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_5 : _GEN_36; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_38 = 5'h6 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_6 : _GEN_37; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_39 = 5'h7 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_7 : _GEN_38; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_40 = 5'h8 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_8 : _GEN_39; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_41 = 5'h9 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_9 : _GEN_40; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_42 = 5'ha == io_in_0_bits_ctrl_rfSrc2 ? REG_1_10 : _GEN_41; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_43 = 5'hb == io_in_0_bits_ctrl_rfSrc2 ? REG_1_11 : _GEN_42; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_44 = 5'hc == io_in_0_bits_ctrl_rfSrc2 ? REG_1_12 : _GEN_43; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_45 = 5'hd == io_in_0_bits_ctrl_rfSrc2 ? REG_1_13 : _GEN_44; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_46 = 5'he == io_in_0_bits_ctrl_rfSrc2 ? REG_1_14 : _GEN_45; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_47 = 5'hf == io_in_0_bits_ctrl_rfSrc2 ? REG_1_15 : _GEN_46; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_48 = 5'h10 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_16 : _GEN_47; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_49 = 5'h11 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_17 : _GEN_48; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_50 = 5'h12 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_18 : _GEN_49; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_51 = 5'h13 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_19 : _GEN_50; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_52 = 5'h14 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_20 : _GEN_51; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_53 = 5'h15 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_21 : _GEN_52; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_54 = 5'h16 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_22 : _GEN_53; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_55 = 5'h17 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_23 : _GEN_54; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_56 = 5'h18 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_24 : _GEN_55; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_57 = 5'h19 == io_in_0_bits_ctrl_rfSrc2 ? REG_1_25 : _GEN_56; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_58 = 5'h1a == io_in_0_bits_ctrl_rfSrc2 ? REG_1_26 : _GEN_57; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_59 = 5'h1b == io_in_0_bits_ctrl_rfSrc2 ? REG_1_27 : _GEN_58; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_60 = 5'h1c == io_in_0_bits_ctrl_rfSrc2 ? REG_1_28 : _GEN_59; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_61 = 5'h1d == io_in_0_bits_ctrl_rfSrc2 ? REG_1_29 : _GEN_60; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_62 = 5'h1e == io_in_0_bits_ctrl_rfSrc2 ? REG_1_30 : _GEN_61; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _GEN_63 = 5'h1f == io_in_0_bits_ctrl_rfSrc2 ? REG_1_31 : _GEN_62; // @[RF.scala 32:36 RF.scala 32:36]
  wire [63:0] _T_59 = io_in_0_bits_ctrl_rfSrc2 == 5'h0 ? 64'h0 : _GEN_63; // @[RF.scala 32:36]
  wire [63:0] _T_60 = io_in_0_bits_ctrl_src2Type ? io_in_0_bits_data_imm : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_61 = src2ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_62 = _T_52 ? io_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_63 = _T_57 ? _T_59 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_64 = _T_60 | _T_61; // @[Mux.scala 27:72]
  wire [63:0] _T_65 = _T_64 | _T_62; // @[Mux.scala 27:72]
  wire  _T_73 = ~io_in_0_bits_ctrl_fuOpType[3] & ~io_in_0_bits_ctrl_fuOpType[5]; // @[LSU.scala 56:49]
  wire [63:0] isuAddr = _T_73 | io_in_0_bits_ctrl_fuOpType[3] ? io_out_bits_data_addr : io_out_bits_data_src1; // @[ISU.scala 80:20]
  wire  _T_81 = io_in_0_bits_ctrl_fuOpType == 7'h20; // @[LSU.scala 57:37]
  wire  _T_87 = io_wb_rfDest != 5'h0 & io_wb_rfDest == io_forward_wb_rfDest & forwardRfWen; // @[ISU.scala 40:100]
  wire [62:0] _T_90 = 63'h1 << io_wb_rfDest; // @[RF.scala 39:39]
  wire [31:0] wbClearMask = io_wb_rfWen & ~_T_87 ? _T_90[31:0] : 32'h0; // @[ISU.scala 94:24]
  wire  _T_92 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [62:0] _T_93 = 63'h1 << io_in_0_bits_ctrl_rfDest; // @[RF.scala 39:39]
  wire [31:0] isuFireSetMask = _T_92 ? _T_93[31:0] : 32'h0; // @[ISU.scala 96:27]
  wire [31:0] _T_100 = ~wbClearMask; // @[RF.scala 45:26]
  wire [31:0] _T_101 = REG & _T_100; // @[RF.scala 45:24]
  wire [31:0] _T_102 = _T_101 | isuFireSetMask; // @[RF.scala 45:38]
  wire [30:0] hi_2 = _T_102[31:1]; // @[RF.scala 45:48]
  wire [31:0] _T_103 = {hi_2,1'h0}; // @[Cat.scala 30:58]
  wire  _T_112 = io_in_0_valid & ~io_out_valid; // @[ISU.scala 106:40]
  wire  _T_115 = io_out_valid & ~_T_92; // @[ISU.scala 107:38]
  wire  _T_116 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_0_ready = ~io_in_0_valid | _T_92; // @[ISU.scala 100:37]
  assign io_out_valid = io_in_0_valid & src1Ready & src2Ready; // @[ISU.scala 57:47]
  assign io_out_bits_cf_instr = io_in_0_bits_cf_instr; // @[ISU.scala 83:18]
  assign io_out_bits_cf_pc = io_in_0_bits_cf_pc; // @[ISU.scala 83:18]
  assign io_out_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[ISU.scala 83:18]
  assign io_out_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[ISU.scala 83:18]
  assign io_out_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[ISU.scala 83:18]
  assign io_out_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[ISU.scala 83:18]
  assign io_out_bits_cf_intrVec_0 = io_in_0_bits_cf_intrVec_0; // @[ISU.scala 83:18]
  assign io_out_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[ISU.scala 83:18]
  assign io_out_bits_cf_intrVec_2 = io_in_0_bits_cf_intrVec_2; // @[ISU.scala 83:18]
  assign io_out_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[ISU.scala 83:18]
  assign io_out_bits_cf_intrVec_4 = io_in_0_bits_cf_intrVec_4; // @[ISU.scala 83:18]
  assign io_out_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[ISU.scala 83:18]
  assign io_out_bits_cf_intrVec_6 = io_in_0_bits_cf_intrVec_6; // @[ISU.scala 83:18]
  assign io_out_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[ISU.scala 83:18]
  assign io_out_bits_cf_intrVec_8 = io_in_0_bits_cf_intrVec_8; // @[ISU.scala 83:18]
  assign io_out_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[ISU.scala 83:18]
  assign io_out_bits_cf_intrVec_10 = io_in_0_bits_cf_intrVec_10; // @[ISU.scala 83:18]
  assign io_out_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[ISU.scala 83:18]
  assign io_out_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[ISU.scala 83:18]
  assign io_out_bits_cf_crossPageIPFFix = io_in_0_bits_cf_crossPageIPFFix; // @[ISU.scala 83:18]
  assign io_out_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[ISU.scala 84:20]
  assign io_out_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[ISU.scala 84:20]
  assign io_out_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[ISU.scala 84:20]
  assign io_out_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[ISU.scala 84:20]
  assign io_out_bits_ctrl_permitLibLoad = isu_perm_lib_ld;
  assign io_out_bits_ctrl_permitLibStore = isu_perm_lib_st;
  assign io_out_bits_ctrl_lsuIsLoad = _T_73 | _T_81; // @[ISU.scala 89:59]
  assign io_out_bits_data_src1 = _T_48 | _T_46; // @[Mux.scala 27:72]
  assign io_out_bits_data_src2 = _T_65 | _T_63; // @[Mux.scala 27:72]
  assign io_out_bits_data_imm = io_in_0_bits_data_imm; // @[ISU.scala 74:25]
  assign io_out_bits_data_addr = io_out_bits_data_src1 + io_out_bits_data_imm; // @[ISU.scala 75:50]
  assign isuAddr_0 = isuAddr;
  always @(posedge clock) begin
    if (reset) begin // @[RF.scala 37:21]
      REG <= 32'h0; // @[RF.scala 37:21]
    end else if (io_flush) begin // @[ISU.scala 97:19]
      REG <= 32'h0; // @[RF.scala 45:10]
    end else begin
      REG <= _T_103; // @[RF.scala 45:10]
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_0 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h0 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_0 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_1 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h1 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_1 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_2 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h2 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_2 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_3 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h3 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_3 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_4 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h4 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_4 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_5 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h5 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_5 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_6 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h6 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_6 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_7 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h7 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_7 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_8 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h8 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_8 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_9 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h9 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_9 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_10 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'ha == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_10 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_11 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'hb == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_11 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_12 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'hc == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_12 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_13 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'hd == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_13 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_14 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'he == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_14 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_15 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'hf == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_15 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_16 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h10 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_16 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_17 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h11 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_17 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_18 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h12 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_18 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_19 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h13 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_19 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_20 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h14 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_20 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_21 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h15 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_21 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_22 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h16 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_22 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_23 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h17 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_23 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_24 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h18 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_24 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_25 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h19 == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_25 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_26 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h1a == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_26 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_27 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h1b == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_27 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_28 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h1c == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_28 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_29 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h1d == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_29 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_30 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h1e == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_30 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
    if (reset) begin // @[RF.scala 31:19]
      REG_1_31 <= 64'h0; // @[RF.scala 31:19]
    end else if (io_wb_rfWen) begin // @[ISU.scala 92:22]
      if (5'h1f == io_wb_rfDest) begin // @[RF.scala 33:50]
        REG_1_31 <= io_wb_rfData; // @[RF.scala 33:50]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  REG_1_0 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  REG_1_1 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  REG_1_2 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  REG_1_3 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  REG_1_4 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  REG_1_5 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  REG_1_6 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  REG_1_7 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  REG_1_8 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  REG_1_9 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  REG_1_10 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  REG_1_11 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  REG_1_12 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  REG_1_13 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  REG_1_14 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  REG_1_15 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  REG_1_16 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  REG_1_17 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  REG_1_18 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  REG_1_19 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  REG_1_20 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  REG_1_21 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  REG_1_22 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  REG_1_23 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  REG_1_24 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  REG_1_25 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  REG_1_26 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  REG_1_27 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  REG_1_28 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  REG_1_29 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  REG_1_30 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  REG_1_31 = _RAND_32[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_ALU(
  input         clock,
  input         reset,
  input         io__in_valid,
  input  [63:0] io__in_bits_src1,
  input  [63:0] io__in_bits_src2,
  input  [6:0]  io__in_bits_func,
  input         io__out_ready,
  output        io__out_valid,
  output [63:0] io__out_bits,
  input  [63:0] io__cfIn_instr,
  input  [38:0] io__cfIn_pc,
  input  [38:0] io__cfIn_pnpc,
  input  [3:0]  io__cfIn_brIdx,
  output [38:0] io__redirect_target,
  output        io__redirect_valid,
  input  [63:0] io__offset,
  output        _T_113_0,
  output        REG_6_0_valid,
  output [38:0] REG_6_0_pc,
  output        REG_6_0_isMissPredict,
  output [38:0] REG_6_0_actualTarget,
  output        REG_6_0_actualTaken,
  output [6:0]  REG_6_0_fuOpType,
  output [1:0]  REG_6_0_btbType,
  output        REG_6_0_isRVC,
  output        io_redirect_valid,
  output [38:0] io_redirect_target
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  isAdderSub = ~io__in_bits_func[6]; // @[ALU.scala 89:20]
  wire [63:0] _T_2 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_3 = io__in_bits_src2 ^ _T_2; // @[ALU.scala 90:33]
  wire [64:0] _T_4 = io__in_bits_src1 + _T_3; // @[ALU.scala 90:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[ALU.scala 90:60]
  wire [64:0] adderRes = _T_4 + _GEN_0; // @[ALU.scala 90:60]
  wire [63:0] xorRes = io__in_bits_src1 ^ io__in_bits_src2; // @[ALU.scala 91:21]
  wire  sltu = ~adderRes[64]; // @[ALU.scala 92:14]
  wire  slt = xorRes[63] ^ sltu; // @[ALU.scala 93:28]
  wire [31:0] lo = io__in_bits_src1[31:0]; // @[ALU.scala 96:35]
  wire [63:0] _T_9 = {32'h0,lo}; // @[Cat.scala 30:58]
  wire [31:0] hi = lo[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_12 = {hi,lo}; // @[Cat.scala 30:58]
  wire [63:0] _T_14 = 7'h25 == io__in_bits_func ? _T_9 : io__in_bits_src1; // @[Mux.scala 80:57]
  wire [63:0] shsrc1 = 7'h2d == io__in_bits_func ? _T_12 : _T_14; // @[Mux.scala 80:57]
  wire [5:0] shamt = io__in_bits_func[5] ? {{1'd0}, io__in_bits_src2[4:0]} : io__in_bits_src2[5:0]; // @[ALU.scala 99:18]
  wire [126:0] _GEN_1 = {{63'd0}, shsrc1}; // @[ALU.scala 101:33]
  wire [126:0] _T_20 = _GEN_1 << shamt; // @[ALU.scala 101:33]
  wire [63:0] _T_22 = {63'h0,slt}; // @[Cat.scala 30:58]
  wire [63:0] _T_23 = {63'h0,sltu}; // @[Cat.scala 30:58]
  wire [63:0] _T_24 = shsrc1 >> shamt; // @[ALU.scala 105:32]
  wire [63:0] _T_25 = io__in_bits_src1 | io__in_bits_src2; // @[ALU.scala 106:30]
  wire [63:0] _T_26 = io__in_bits_src1 & io__in_bits_src2; // @[ALU.scala 107:30]
  wire [63:0] _T_27 = 7'h2d == io__in_bits_func ? _T_12 : _T_14; // @[ALU.scala 108:32]
  wire [63:0] _T_29 = $signed(_T_27) >>> shamt; // @[ALU.scala 108:49]
  wire [64:0] _T_31 = 4'h1 == io__in_bits_func[3:0] ? {{1'd0}, _T_20[63:0]} : adderRes; // @[Mux.scala 80:57]
  wire [64:0] _T_33 = 4'h2 == io__in_bits_func[3:0] ? {{1'd0}, _T_22} : _T_31; // @[Mux.scala 80:57]
  wire [64:0] _T_35 = 4'h3 == io__in_bits_func[3:0] ? {{1'd0}, _T_23} : _T_33; // @[Mux.scala 80:57]
  wire [64:0] _T_37 = 4'h4 == io__in_bits_func[3:0] ? {{1'd0}, xorRes} : _T_35; // @[Mux.scala 80:57]
  wire [64:0] _T_39 = 4'h5 == io__in_bits_func[3:0] ? {{1'd0}, _T_24} : _T_37; // @[Mux.scala 80:57]
  wire [64:0] _T_41 = 4'h6 == io__in_bits_func[3:0] ? {{1'd0}, _T_25} : _T_39; // @[Mux.scala 80:57]
  wire [64:0] _T_43 = 4'h7 == io__in_bits_func[3:0] ? {{1'd0}, _T_26} : _T_41; // @[Mux.scala 80:57]
  wire [64:0] res = 4'hd == io__in_bits_func[3:0] ? {{1'd0}, _T_29} : _T_43; // @[Mux.scala 80:57]
  wire [31:0] lo_2 = res[31:0]; // @[ALU.scala 110:57]
  wire [31:0] hi_1 = lo_2[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_48 = {hi_1,lo_2}; // @[Cat.scala 30:58]
  wire [64:0] aluRes = io__in_bits_func[5] ? {{1'd0}, _T_48} : res; // @[ALU.scala 110:19]
  wire  _T_50 = ~(|xorRes); // @[ALU.scala 113:48]
  wire  isBranch = ~io__in_bits_func[3]; // @[ALU.scala 65:30]
  wire  isBru = io__in_bits_func[4]; // @[ALU.scala 64:31]
  wire  _T_53 = 2'h0 == io__in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_54 = 2'h2 == io__in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_55 = 2'h3 == io__in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_60 = _T_53 & _T_50 | _T_54 & slt | _T_55 & sltu; // @[Mux.scala 27:72]
  wire  taken = _T_60 ^ io__in_bits_func[0]; // @[ALU.scala 120:72]
  wire [63:0] _GEN_2 = {{25'd0}, io__cfIn_pc}; // @[ALU.scala 121:41]
  wire [63:0] _T_63 = _GEN_2 + io__offset; // @[ALU.scala 121:41]
  wire [64:0] _T_64 = isBranch ? {{1'd0}, _T_63} : adderRes; // @[ALU.scala 121:19]
  wire [38:0] target = _T_64[38:0]; // @[ALU.scala 121:63]
  wire  _T_66 = ~taken & isBranch; // @[ALU.scala 122:33]
  wire  predictWrong = ~taken & isBranch ? io__cfIn_brIdx[0] : ~io__cfIn_brIdx[0] | io__redirect_target != io__cfIn_pnpc
    ; // @[ALU.scala 122:25]
  wire  isRVC = io__cfIn_instr[1:0] != 2'h3; // @[ALU.scala 123:35]
  wire  _T_83 = ~isRVC; // @[ALU.scala 125:55]
  wire [38:0] _T_92 = io__cfIn_pc + 39'h2; // @[ALU.scala 126:71]
  wire [38:0] _T_94 = io__cfIn_pc + 39'h4; // @[ALU.scala 126:89]
  wire [38:0] _T_95 = isRVC ? _T_92 : _T_94; // @[ALU.scala 126:52]
  wire  _T_97 = io__in_valid & isBru; // @[ALU.scala 128:30]
  wire  _T_98 = io__in_valid & isBru & predictWrong; // @[ALU.scala 128:39]
  wire [24:0] hi_2 = io__cfIn_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_102 = {hi_2,io__cfIn_pc}; // @[Cat.scala 30:58]
  wire [63:0] _T_104 = _T_102 + 64'h4; // @[ALU.scala 134:71]
  wire [63:0] _T_109 = _T_102 + 64'h2; // @[ALU.scala 134:108]
  wire [63:0] _T_110 = _T_83 ? _T_104 : _T_109; // @[ALU.scala 134:32]
  wire [64:0] _T_111 = isBru ? {{1'd0}, _T_110} : aluRes; // @[ALU.scala 134:21]
  wire  _T_113 = io__in_valid & io__in_bits_func == 7'h7e; // @[ALU.scala 139:31]
  wire  _T_125 = io__in_bits_func == 7'h58 | io__in_bits_func == 7'h5c; // @[ALU.scala 143:180]
  wire  _T_126 = io__in_bits_func == 7'h5a; // @[ALU.scala 143:214]
  wire  _T_127 = io__in_bits_func == 7'h5e; // @[ALU.scala 143:239]
  wire  _T_142 = 7'h5c == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_143 = 7'h5e == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_144 = 7'h58 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_145 = 7'h5a == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire [1:0] _T_153 = _T_143 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_155 = _T_145 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_3 = {{1'd0}, _T_142}; // @[Mux.scala 27:72]
  wire [1:0] _T_162 = _GEN_3 | _T_153; // @[Mux.scala 27:72]
  wire [1:0] _GEN_4 = {{1'd0}, _T_144}; // @[Mux.scala 27:72]
  wire [1:0] _T_163 = _T_162 | _GEN_4; // @[Mux.scala 27:72]
  wire [1:0] _T_164 = _T_163 | _T_155; // @[Mux.scala 27:72]
  reg  REG_6_valid; // @[ALU.scala 166:34]
  reg [38:0] REG_6_pc; // @[ALU.scala 166:34]
  reg  REG_6_isMissPredict; // @[ALU.scala 166:34]
  reg [38:0] REG_6_actualTarget; // @[ALU.scala 166:34]
  reg  REG_6_actualTaken; // @[ALU.scala 166:34]
  reg [6:0] REG_6_fuOpType; // @[ALU.scala 166:34]
  reg [1:0] REG_6_btbType; // @[ALU.scala 166:34]
  reg  REG_6_isRVC; // @[ALU.scala 166:34]
  wire  _T_200 = _T_97 & ~predictWrong; // @[ALU.scala 168:32]
  wire  _T_203 = _T_200 & isBranch; // @[ALU.scala 170:33]
  wire  _T_204 = _T_98 & isBranch; // @[ALU.scala 171:33]
  wire  _T_208 = _T_204 & io__cfIn_pc[2:0] == 3'h0; // @[ALU.scala 172:45]
  wire  _T_209 = _T_204 & io__cfIn_pc[2:0] == 3'h0 & isRVC; // @[ALU.scala 172:73]
  wire  _T_215 = _T_208 & _T_83; // @[ALU.scala 173:73]
  wire  _T_219 = _T_204 & io__cfIn_pc[2:0] == 3'h2; // @[ALU.scala 174:45]
  wire  _T_220 = _T_204 & io__cfIn_pc[2:0] == 3'h2 & isRVC; // @[ALU.scala 174:73]
  wire  _T_226 = _T_219 & _T_83; // @[ALU.scala 175:73]
  wire  _T_230 = _T_204 & io__cfIn_pc[2:0] == 3'h4; // @[ALU.scala 176:45]
  wire  _T_231 = _T_204 & io__cfIn_pc[2:0] == 3'h4 & isRVC; // @[ALU.scala 176:73]
  wire  _T_237 = _T_230 & _T_83; // @[ALU.scala 177:73]
  wire  _T_241 = _T_204 & io__cfIn_pc[2:0] == 3'h6; // @[ALU.scala 178:45]
  wire  _T_242 = _T_204 & io__cfIn_pc[2:0] == 3'h6 & isRVC; // @[ALU.scala 178:73]
  wire  _T_248 = _T_241 & _T_83; // @[ALU.scala 179:73]
  wire  _T_252 = _T_200 & _T_125; // @[ALU.scala 180:33]
  wire  _T_256 = _T_98 & _T_125; // @[ALU.scala 181:33]
  wire  _T_258 = _T_200 & _T_126; // @[ALU.scala 182:33]
  wire  _T_260 = _T_98 & _T_126; // @[ALU.scala 183:33]
  wire  _T_262 = _T_200 & _T_127; // @[ALU.scala 184:33]
  wire  _T_264 = _T_98 & _T_127; // @[ALU.scala 185:33]
  assign io__out_valid = io__in_valid; // @[ALU.scala 153:16]
  assign io__out_bits = _T_111[63:0]; // @[ALU.scala 134:15]
  assign io__redirect_target = _T_66 ? _T_95 : target; // @[ALU.scala 126:28]
  assign io__redirect_valid = io__in_valid & isBru & predictWrong; // @[ALU.scala 128:39]
  assign _T_113_0 = _T_113;
  assign REG_6_0_valid = REG_6_valid;
  assign REG_6_0_pc = REG_6_pc;
  assign REG_6_0_isMissPredict = REG_6_isMissPredict;
  assign REG_6_0_actualTarget = REG_6_actualTarget;
  assign REG_6_0_actualTaken = REG_6_actualTaken;
  assign REG_6_0_fuOpType = REG_6_fuOpType;
  assign REG_6_0_btbType = REG_6_btbType;
  assign REG_6_0_isRVC = REG_6_isRVC;
  assign io_redirect_valid = io__redirect_valid;
  assign io_redirect_target = io__redirect_target;
  always @(posedge clock) begin
    if (reset) begin // @[ALU.scala 166:34]
      REG_6_valid <= 1'h0; // @[ALU.scala 166:34]
    end else begin
      REG_6_valid <= _T_97; // @[ALU.scala 166:34]
    end
    if (reset) begin // @[ALU.scala 166:34]
      REG_6_pc <= 39'h0; // @[ALU.scala 166:34]
    end else begin
      REG_6_pc <= io__cfIn_pc; // @[ALU.scala 166:34]
    end
    if (reset) begin // @[ALU.scala 166:34]
      REG_6_isMissPredict <= 1'h0; // @[ALU.scala 166:34]
    end else if (~taken & isBranch) begin // @[ALU.scala 122:25]
      REG_6_isMissPredict <= io__cfIn_brIdx[0];
    end else begin
      REG_6_isMissPredict <= ~io__cfIn_brIdx[0] | io__redirect_target != io__cfIn_pnpc;
    end
    if (reset) begin // @[ALU.scala 166:34]
      REG_6_actualTarget <= 39'h0; // @[ALU.scala 166:34]
    end else begin
      REG_6_actualTarget <= target; // @[ALU.scala 166:34]
    end
    if (reset) begin // @[ALU.scala 166:34]
      REG_6_actualTaken <= 1'h0; // @[ALU.scala 166:34]
    end else begin
      REG_6_actualTaken <= taken; // @[ALU.scala 166:34]
    end
    if (reset) begin // @[ALU.scala 166:34]
      REG_6_fuOpType <= 7'h0; // @[ALU.scala 166:34]
    end else begin
      REG_6_fuOpType <= io__in_bits_func; // @[ALU.scala 166:34]
    end
    if (reset) begin // @[ALU.scala 166:34]
      REG_6_btbType <= 2'h0; // @[ALU.scala 166:34]
    end else begin
      REG_6_btbType <= _T_164; // @[ALU.scala 166:34]
    end
    if (reset) begin // @[ALU.scala 166:34]
      REG_6_isRVC <= 1'h0; // @[ALU.scala 166:34]
    end else begin
      REG_6_isRVC <= isRVC; // @[ALU.scala 166:34]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(io__cfIn_instr[1:0] == 2'h3 | isRVC | ~io__in_valid | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ALU.scala:124 assert(io.cfIn.instr(1,0) === \"b11\".U || isRVC || !valid)\n"); // @[ALU.scala 124:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(io__cfIn_instr[1:0] == 2'h3 | isRVC | ~io__in_valid | reset)) begin
          $fatal; // @[ALU.scala 124:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG_6_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  REG_6_pc = _RAND_1[38:0];
  _RAND_2 = {1{`RANDOM}};
  REG_6_isMissPredict = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  REG_6_actualTarget = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  REG_6_actualTaken = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG_6_fuOpType = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  REG_6_btbType = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  REG_6_isRVC = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_LSExecUnit(
  input         clock,
  input         reset,
  input         io__in_valid,
  input  [63:0] io__in_bits_src1,
  input  [6:0]  io__in_bits_func,
  input         io__out_ready,
  output        io__out_valid,
  output [63:0] io__out_bits,
  input  [63:0] io__wdata,
  input         io__dmem_req_ready,
  output        io__dmem_req_valid,
  output [38:0] io__dmem_req_bits_addr,
  output [2:0]  io__dmem_req_bits_size,
  output [3:0]  io__dmem_req_bits_cmd,
  output [7:0]  io__dmem_req_bits_wmask,
  output [63:0] io__dmem_req_bits_wdata,
  output        io__dmem_resp_ready,
  input         io__dmem_resp_valid,
  input  [63:0] io__dmem_resp_bits_rdata,
  output        io__isMMIO,
  output        io__dtlbPF,
  output        io__loadAddrMisaligned,
  output        io__storeAddrMisaligned,
  input         DTLBPF,
  input         DTLBENABLE,
  input         ISAMO2,
  output [63:0] io_in_bits_src1,
  input         DTLBFINISH
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] addrLatch; // @[UnpipelinedLSU.scala 342:26]
  wire  isStore = io__in_valid & io__in_bits_func[3]; // @[UnpipelinedLSU.scala 343:23]
  wire  _T_1 = ~isStore; // @[UnpipelinedLSU.scala 344:21]
  wire  partialLoad = ~isStore & io__in_bits_func != 7'h3; // @[UnpipelinedLSU.scala 344:30]
  reg [1:0] state; // @[UnpipelinedLSU.scala 347:22]
  wire  _T_3 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = io__dmem_req_ready & io__dmem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_9 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_2 = DTLBFINISH & DTLBPF ? 2'h0 : state; // @[UnpipelinedLSU.scala 367:36 UnpipelinedLSU.scala 367:44 UnpipelinedLSU.scala 347:22]
  wire  _T_13 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_14 = io__dmem_resp_ready & io__dmem_resp_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_15 = partialLoad ? 2'h3 : 2'h0; // @[UnpipelinedLSU.scala 370:62]
  wire [1:0] _GEN_4 = _T_14 ? _T_15 : state; // @[UnpipelinedLSU.scala 370:48 UnpipelinedLSU.scala 370:56 UnpipelinedLSU.scala 347:22]
  wire  _T_16 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_5 = _T_16 ? 2'h0 : state; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 371:32 UnpipelinedLSU.scala 347:22]
  wire [7:0] hi = io__wdata[7:0]; // @[UnpipelinedLSU.scala 319:30]
  wire [63:0] _T_34 = {hi,hi,hi,hi,hi,hi,hi,hi}; // @[Cat.scala 30:58]
  wire [15:0] hi_3 = io__wdata[15:0]; // @[UnpipelinedLSU.scala 320:30]
  wire [63:0] _T_35 = {hi_3,hi_3,hi_3,hi_3}; // @[Cat.scala 30:58]
  wire [31:0] hi_5 = io__wdata[31:0]; // @[UnpipelinedLSU.scala 321:30]
  wire [63:0] _T_36 = {hi_5,hi_5}; // @[Cat.scala 30:58]
  wire  _T_37 = 2'h0 == io__in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_38 = 2'h1 == io__in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_39 = 2'h2 == io__in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_40 = 2'h3 == io__in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_41 = _T_37 ? _T_34 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_42 = _T_38 ? _T_35 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_43 = _T_39 ? _T_36 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_44 = _T_40 ? io__wdata : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = _T_41 | _T_42; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = _T_45 | _T_43; // @[Mux.scala 27:72]
  wire [1:0] _T_53 = _T_38 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_54 = _T_39 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_55 = _T_40 ? 8'hff : 8'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_13 = {{1'd0}, _T_37}; // @[Mux.scala 27:72]
  wire [1:0] _T_56 = _GEN_13 | _T_53; // @[Mux.scala 27:72]
  wire [3:0] _GEN_14 = {{2'd0}, _T_56}; // @[Mux.scala 27:72]
  wire [3:0] _T_57 = _GEN_14 | _T_54; // @[Mux.scala 27:72]
  wire [7:0] _GEN_15 = {{4'd0}, _T_57}; // @[Mux.scala 27:72]
  wire [7:0] _T_58 = _GEN_15 | _T_55; // @[Mux.scala 27:72]
  wire [14:0] _GEN_16 = {{7'd0}, _T_58}; // @[UnpipelinedLSU.scala 315:8]
  wire [14:0] reqWmask = _GEN_16 << io__in_bits_src1[2:0]; // @[UnpipelinedLSU.scala 315:8]
  wire  _T_75 = partialLoad ? state == 2'h3 : _T_14 & state == 2'h2; // @[UnpipelinedLSU.scala 391:114]
  reg [63:0] rdataLatch; // @[UnpipelinedLSU.scala 397:27]
  wire  _T_93 = 3'h0 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_94 = 3'h1 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_95 = 3'h2 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_96 = 3'h3 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_97 = 3'h4 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_98 = 3'h5 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_99 = 3'h6 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_100 = 3'h7 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_101 = _T_93 ? rdataLatch : 64'h0; // @[Mux.scala 27:72]
  wire [55:0] _T_102 = _T_94 ? rdataLatch[63:8] : 56'h0; // @[Mux.scala 27:72]
  wire [47:0] _T_103 = _T_95 ? rdataLatch[63:16] : 48'h0; // @[Mux.scala 27:72]
  wire [39:0] _T_104 = _T_96 ? rdataLatch[63:24] : 40'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_105 = _T_97 ? rdataLatch[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [23:0] _T_106 = _T_98 ? rdataLatch[63:40] : 24'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_107 = _T_99 ? rdataLatch[63:48] : 16'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_108 = _T_100 ? rdataLatch[63:56] : 8'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_17 = {{8'd0}, _T_102}; // @[Mux.scala 27:72]
  wire [63:0] _T_109 = _T_101 | _GEN_17; // @[Mux.scala 27:72]
  wire [63:0] _GEN_18 = {{16'd0}, _T_103}; // @[Mux.scala 27:72]
  wire [63:0] _T_110 = _T_109 | _GEN_18; // @[Mux.scala 27:72]
  wire [63:0] _GEN_19 = {{24'd0}, _T_104}; // @[Mux.scala 27:72]
  wire [63:0] _T_111 = _T_110 | _GEN_19; // @[Mux.scala 27:72]
  wire [63:0] _GEN_20 = {{32'd0}, _T_105}; // @[Mux.scala 27:72]
  wire [63:0] _T_112 = _T_111 | _GEN_20; // @[Mux.scala 27:72]
  wire [63:0] _GEN_21 = {{40'd0}, _T_106}; // @[Mux.scala 27:72]
  wire [63:0] _T_113 = _T_112 | _GEN_21; // @[Mux.scala 27:72]
  wire [63:0] _GEN_22 = {{48'd0}, _T_107}; // @[Mux.scala 27:72]
  wire [63:0] _T_114 = _T_113 | _GEN_22; // @[Mux.scala 27:72]
  wire [63:0] _GEN_23 = {{56'd0}, _T_108}; // @[Mux.scala 27:72]
  wire [63:0] rdataSel = _T_114 | _GEN_23; // @[Mux.scala 27:72]
  wire [7:0] lo = rdataSel[7:0]; // @[UnpipelinedLSU.scala 416:41]
  wire [55:0] hi_6 = lo[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_134 = {hi_6,lo}; // @[Cat.scala 30:58]
  wire [15:0] lo_1 = rdataSel[15:0]; // @[UnpipelinedLSU.scala 417:41]
  wire [47:0] hi_7 = lo_1[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_137 = {hi_7,lo_1}; // @[Cat.scala 30:58]
  wire [31:0] lo_2 = rdataSel[31:0]; // @[UnpipelinedLSU.scala 418:41]
  wire [31:0] hi_8 = lo_2[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_140 = {hi_8,lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _T_141 = {56'h0,lo}; // @[Cat.scala 30:58]
  wire [63:0] _T_142 = {48'h0,lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _T_143 = {32'h0,lo_2}; // @[Cat.scala 30:58]
  wire  _T_144 = 7'h0 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_145 = 7'h1 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_146 = 7'h2 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_147 = 7'h4 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_148 = 7'h5 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_149 = 7'h6 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire [63:0] _T_150 = _T_144 ? _T_134 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_151 = _T_145 ? _T_137 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_152 = _T_146 ? _T_140 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_153 = _T_147 ? _T_141 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_154 = _T_148 ? _T_142 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_155 = _T_149 ? _T_143 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_156 = _T_150 | _T_151; // @[Mux.scala 27:72]
  wire [63:0] _T_157 = _T_156 | _T_152; // @[Mux.scala 27:72]
  wire [63:0] _T_158 = _T_157 | _T_153; // @[Mux.scala 27:72]
  wire [63:0] _T_159 = _T_158 | _T_154; // @[Mux.scala 27:72]
  wire [63:0] rdataPartialLoad = _T_159 | _T_155; // @[Mux.scala 27:72]
  wire  _T_163 = ~io__in_bits_src1[0]; // @[UnpipelinedLSU.scala 425:27]
  wire  _T_165 = io__in_bits_src1[1:0] == 2'h0; // @[UnpipelinedLSU.scala 426:29]
  wire  _T_167 = io__in_bits_src1[2:0] == 3'h0; // @[UnpipelinedLSU.scala 427:29]
  wire  addrAligned = _T_37 | _T_38 & _T_163 | _T_39 & _T_165 | _T_40 & _T_167; // @[Mux.scala 27:72]
  wire  _T_185 = ~addrAligned; // @[UnpipelinedLSU.scala 438:60]
  wire  _T_199 = ~io__dmem_req_bits_cmd[0] & ~io__dmem_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_200 = io__dmem_req_valid & _T_199; // @[SimpleBus.scala 104:29]
  wire  _T_202 = _T_200 & _T_4; // @[UnpipelinedLSU.scala 443:39]
  reg  REG_5; // @[StopWatch.scala 24:20]
  wire  _GEN_9 = _T_200 | REG_5; // @[StopWatch.scala 30:20 StopWatch.scala 30:24 StopWatch.scala 24:20]
  wire  _T_211 = io__dmem_req_valid & io__dmem_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  reg  REG_6; // @[StopWatch.scala 24:20]
  wire  _GEN_11 = _T_211 | REG_6; // @[StopWatch.scala 30:20 StopWatch.scala 30:24 StopWatch.scala 24:20]
  assign io__out_valid = DTLBPF & state != 2'h0 | io__loadAddrMisaligned | io__storeAddrMisaligned | _T_75; // @[UnpipelinedLSU.scala 391:22]
  assign io__out_bits = partialLoad ? rdataPartialLoad : io__dmem_resp_bits_rdata; // @[UnpipelinedLSU.scala 430:21]
  assign io__dmem_req_valid = io__in_valid & state == 2'h0 & ~io__loadAddrMisaligned & ~io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 388:75]
  assign io__dmem_req_bits_addr = io__in_bits_src1[38:0]; // @[UnpipelinedLSU.scala 379:68]
  assign io__dmem_req_bits_size = {{1'd0}, io__in_bits_func[1:0]}; // @[UnpipelinedLSU.scala 378:18]
  assign io__dmem_req_bits_cmd = {{3'd0}, isStore}; // @[UnpipelinedLSU.scala 343:23]
  assign io__dmem_req_bits_wmask = reqWmask[7:0]; // @[SimpleBus.scala 68:16]
  assign io__dmem_req_bits_wdata = _T_46 | _T_44; // @[Mux.scala 27:72]
  assign io__dmem_resp_ready = 1'h1; // @[UnpipelinedLSU.scala 389:19]
  assign io__isMMIO = 1'h0;
  assign io__dtlbPF = DTLBPF; // @[UnpipelinedLSU.scala 358:13]
  assign io__loadAddrMisaligned = io__in_valid & _T_1 & ~ISAMO2 & ~addrAligned; // @[UnpipelinedLSU.scala 438:57]
  assign io__storeAddrMisaligned = io__in_valid & (isStore | ISAMO2) & _T_185; // @[UnpipelinedLSU.scala 439:57]
  assign io_in_bits_src1 = io__in_bits_src1;
  always @(posedge clock) begin
    if (reset) begin // @[UnpipelinedLSU.scala 342:26]
      addrLatch <= 64'h0; // @[UnpipelinedLSU.scala 342:26]
    end else begin
      addrLatch <= io__in_bits_src1; // @[UnpipelinedLSU.scala 342:26]
    end
    if (reset) begin // @[UnpipelinedLSU.scala 347:22]
      state <= 2'h0; // @[UnpipelinedLSU.scala 347:22]
    end else if (_T_3) begin // @[Conditional.scala 40:58]
      if (_T_4 & ~DTLBENABLE) begin // @[UnpipelinedLSU.scala 363:45]
        state <= 2'h2; // @[UnpipelinedLSU.scala 363:53]
      end else if (_T_4 & DTLBENABLE) begin // @[UnpipelinedLSU.scala 362:45]
        state <= 2'h1; // @[UnpipelinedLSU.scala 362:53]
      end
    end else if (_T_9) begin // @[Conditional.scala 39:67]
      if (DTLBFINISH & ~DTLBPF) begin // @[UnpipelinedLSU.scala 368:36]
        state <= 2'h2; // @[UnpipelinedLSU.scala 368:44]
      end else begin
        state <= _GEN_2;
      end
    end else if (_T_13) begin // @[Conditional.scala 39:67]
      state <= _GEN_4;
    end else begin
      state <= _GEN_5;
    end
    if (reset) begin // @[UnpipelinedLSU.scala 397:27]
      rdataLatch <= 64'h0; // @[UnpipelinedLSU.scala 397:27]
    end else begin
      rdataLatch <= io__dmem_resp_bits_rdata; // @[UnpipelinedLSU.scala 397:27]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_5 <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (_T_14) begin // @[StopWatch.scala 31:19]
      REG_5 <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      REG_5 <= _GEN_9;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_6 <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (_T_14) begin // @[StopWatch.scala 31:19]
      REG_6 <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      REG_6 <= _GEN_11;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  addrLatch = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
  _RAND_2 = {2{`RANDOM}};
  rdataLatch = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  REG_5 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_6 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_AtomALU(
  input  [63:0] io_src1,
  input  [63:0] io_src2,
  input  [6:0]  io_func,
  input         io_isWordOp,
  output [63:0] io_result
);
  wire  isAdderSub = ~io_func[6]; // @[LSU.scala 184:20]
  wire [63:0] _T_2 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_3 = io_src2 ^ _T_2; // @[LSU.scala 185:33]
  wire [64:0] _T_4 = io_src1 + _T_3; // @[LSU.scala 185:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[LSU.scala 185:60]
  wire [64:0] adderRes = _T_4 + _GEN_0; // @[LSU.scala 185:60]
  wire [63:0] xorRes = io_src1 ^ io_src2; // @[LSU.scala 186:21]
  wire  sltu = ~adderRes[64]; // @[LSU.scala 187:14]
  wire  slt = xorRes[63] ^ sltu; // @[LSU.scala 188:28]
  wire [63:0] _T_9 = io_src1 & io_src2; // @[LSU.scala 194:32]
  wire [63:0] _T_10 = io_src1 | io_src2; // @[LSU.scala 195:32]
  wire [63:0] _T_12 = slt ? io_src1 : io_src2; // @[LSU.scala 196:29]
  wire [63:0] _T_14 = slt ? io_src2 : io_src1; // @[LSU.scala 197:29]
  wire [63:0] _T_16 = sltu ? io_src1 : io_src2; // @[LSU.scala 198:29]
  wire [63:0] _T_18 = sltu ? io_src2 : io_src1; // @[LSU.scala 199:29]
  wire [64:0] _T_20 = 6'h22 == io_func[5:0] ? {{1'd0}, io_src2} : adderRes; // @[Mux.scala 80:57]
  wire [64:0] _T_22 = 6'h24 == io_func[5:0] ? {{1'd0}, xorRes} : _T_20; // @[Mux.scala 80:57]
  wire [64:0] _T_24 = 6'h25 == io_func[5:0] ? {{1'd0}, _T_9} : _T_22; // @[Mux.scala 80:57]
  wire [64:0] _T_26 = 6'h26 == io_func[5:0] ? {{1'd0}, _T_10} : _T_24; // @[Mux.scala 80:57]
  wire [64:0] _T_28 = 6'h37 == io_func[5:0] ? {{1'd0}, _T_12} : _T_26; // @[Mux.scala 80:57]
  wire [64:0] _T_30 = 6'h30 == io_func[5:0] ? {{1'd0}, _T_14} : _T_28; // @[Mux.scala 80:57]
  wire [64:0] _T_32 = 6'h31 == io_func[5:0] ? {{1'd0}, _T_16} : _T_30; // @[Mux.scala 80:57]
  wire [64:0] res = 6'h32 == io_func[5:0] ? {{1'd0}, _T_18} : _T_32; // @[Mux.scala 80:57]
  wire [31:0] lo = res[31:0]; // @[LSU.scala 202:45]
  wire [31:0] hi = lo[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_36 = {hi,lo}; // @[Cat.scala 30:58]
  assign io_result = io_isWordOp ? _T_36 : res[63:0]; // @[LSU.scala 202:20]
endmodule
module ysyx_210000_UnpipelinedLSU(
  input         clock,
  input         reset,
  input         io__in_valid,
  input  [63:0] io__in_bits_src1,
  input  [6:0]  io__in_bits_func,
  input         io__out_ready,
  output        io__out_valid,
  output [63:0] io__out_bits,
  input  [63:0] io__srcSum,
  input  [63:0] io__wdata,
  input  [31:0] io__instr,
  input         io__dmem_req_ready,
  output        io__dmem_req_valid,
  output [38:0] io__dmem_req_bits_addr,
  output [2:0]  io__dmem_req_bits_size,
  output [3:0]  io__dmem_req_bits_cmd,
  output [7:0]  io__dmem_req_bits_wmask,
  output [63:0] io__dmem_req_bits_wdata,
  input         io__dmem_resp_valid,
  input  [63:0] io__dmem_resp_bits_rdata,
  output        io__dtlbPF,
  output        io__loadAddrMisaligned,
  output        io__storeAddrMisaligned,
  output        setLr_0,
  input         DTLBPF,
  output        amoReq_0,
  input         cannot_access_memory,
  input         DTLBENABLE,
  output [63:0] io_in_bits_src1,
  input         DTLBFINISH,
  output        _T_20_0,
  output [63:0] setLrAddr_0,
  output [63:0] _T_28_0,
  output        setLrVal_0,
  input  [63:0] lr_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  lsExecUnit_clock; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_reset; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_io__in_valid; // @[UnpipelinedLSU.scala 48:28]
  wire [63:0] lsExecUnit_io__in_bits_src1; // @[UnpipelinedLSU.scala 48:28]
  wire [6:0] lsExecUnit_io__in_bits_func; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_io__out_ready; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_io__out_valid; // @[UnpipelinedLSU.scala 48:28]
  wire [63:0] lsExecUnit_io__out_bits; // @[UnpipelinedLSU.scala 48:28]
  wire [63:0] lsExecUnit_io__wdata; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_io__dmem_req_ready; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_io__dmem_req_valid; // @[UnpipelinedLSU.scala 48:28]
  wire [38:0] lsExecUnit_io__dmem_req_bits_addr; // @[UnpipelinedLSU.scala 48:28]
  wire [2:0] lsExecUnit_io__dmem_req_bits_size; // @[UnpipelinedLSU.scala 48:28]
  wire [3:0] lsExecUnit_io__dmem_req_bits_cmd; // @[UnpipelinedLSU.scala 48:28]
  wire [7:0] lsExecUnit_io__dmem_req_bits_wmask; // @[UnpipelinedLSU.scala 48:28]
  wire [63:0] lsExecUnit_io__dmem_req_bits_wdata; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_io__dmem_resp_ready; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_io__dmem_resp_valid; // @[UnpipelinedLSU.scala 48:28]
  wire [63:0] lsExecUnit_io__dmem_resp_bits_rdata; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_io__isMMIO; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_io__dtlbPF; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_io__loadAddrMisaligned; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_DTLBPF; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_DTLBENABLE; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_ISAMO2; // @[UnpipelinedLSU.scala 48:28]
  wire [63:0] lsExecUnit_io_in_bits_src1; // @[UnpipelinedLSU.scala 48:28]
  wire  lsExecUnit_DTLBFINISH; // @[UnpipelinedLSU.scala 48:28]
  wire [63:0] atomALU_io_src1; // @[UnpipelinedLSU.scala 100:25]
  wire [63:0] atomALU_io_src2; // @[UnpipelinedLSU.scala 100:25]
  wire [6:0] atomALU_io_func; // @[UnpipelinedLSU.scala 100:25]
  wire  atomALU_io_isWordOp; // @[UnpipelinedLSU.scala 100:25]
  wire [63:0] atomALU_io_result; // @[UnpipelinedLSU.scala 100:25]
  wire  _T_5 = ~io__in_bits_func[3] & ~io__in_bits_func[5]; // @[LSU.scala 56:49]
  wire  atomReq = io__in_valid & io__in_bits_func[5]; // @[UnpipelinedLSU.scala 55:26]
  wire  _T_8 = io__in_bits_func == 7'h20; // @[LSU.scala 57:37]
  wire  _T_11 = io__in_bits_func == 7'h21; // @[LSU.scala 58:37]
  wire  _T_13 = io__in_bits_func[5] & ~_T_8 & ~_T_11; // @[LSU.scala 59:61]
  wire  amoReq = io__in_valid & _T_13; // @[UnpipelinedLSU.scala 56:26]
  wire  lrReq = io__in_valid & _T_8; // @[UnpipelinedLSU.scala 57:25]
  wire  scReq = io__in_valid & _T_11; // @[UnpipelinedLSU.scala 58:25]
  wire [2:0] funct3 = io__instr[14:12]; // @[UnpipelinedLSU.scala 66:26]
  wire  scInvalid = ~(io__in_bits_src1 == lr_addr) & scReq; // @[UnpipelinedLSU.scala 83:40]
  reg [2:0] state; // @[UnpipelinedLSU.scala 97:24]
  reg [63:0] atomMemReg; // @[UnpipelinedLSU.scala 98:29]
  reg [63:0] atomRegReg; // @[UnpipelinedLSU.scala 99:29]
  wire  _T_20 = io__in_valid & ~scInvalid; // @[UnpipelinedLSU.scala 111:33]
  wire [63:0] _T_28 = _T_5 | io__in_bits_func[3] ? io__srcSum : io__in_bits_src1; // @[UnpipelinedLSU.scala 113:30]
  wire  _T_29 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_34 = ~cannot_access_memory; // @[UnpipelinedLSU.scala 147:23]
  wire  _T_36 = ~atomReq; // @[UnpipelinedLSU.scala 150:56]
  wire  _T_40 = lsExecUnit_io__out_ready & lsExecUnit_io__out_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_1 = amoReq & _T_34 ? 3'h5 : 3'h0; // @[UnpipelinedLSU.scala 161:44 UnpipelinedLSU.scala 161:51 UnpipelinedLSU.scala 158:17]
  wire [2:0] _GEN_2 = lrReq & _T_34 ? 3'h3 : _GEN_1; // @[UnpipelinedLSU.scala 162:43 UnpipelinedLSU.scala 162:50]
  wire [2:0] _T_51 = scInvalid ? 3'h0 : 3'h4; // @[UnpipelinedLSU.scala 163:56]
  wire  _T_52 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_4 = io__out_valid ? 3'h0 : state; // @[UnpipelinedLSU.scala 177:28 UnpipelinedLSU.scala 177:35 UnpipelinedLSU.scala 97:24]
  wire  _T_65 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [1:0] _T_66 = funct3[0] ? 2'h3 : 2'h2; // @[UnpipelinedLSU.scala 197:42]
  wire [2:0] _GEN_5 = _T_40 ? 3'h6 : state; // @[UnpipelinedLSU.scala 201:39 UnpipelinedLSU.scala 202:17 UnpipelinedLSU.scala 97:24]
  wire  _T_71 = 3'h6 == state; // @[Conditional.scala 37:30]
  wire  _T_75 = 3'h7 == state; // @[Conditional.scala 37:30]
  wire [3:0] _T_76 = funct3[0] ? 4'hb : 4'ha; // @[UnpipelinedLSU.scala 228:42]
  wire [2:0] _GEN_6 = _T_40 ? 3'h0 : state; // @[UnpipelinedLSU.scala 232:39 UnpipelinedLSU.scala 233:17 UnpipelinedLSU.scala 97:24]
  wire  _T_83 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_91 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [63:0] _GEN_11 = io__in_bits_src1; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 254:36]
  wire  _GEN_14 = _T_91 & _T_40; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 258:36 UnpipelinedLSU.scala 135:32]
  wire [2:0] _GEN_16 = _T_91 ? _GEN_6 : state; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 97:24]
  wire  _GEN_17 = _T_83 | _T_91; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 238:36]
  wire [3:0] _GEN_20 = _T_83 ? {{2'd0}, _T_66} : _T_76; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 242:36]
  wire  _GEN_22 = _T_83 ? _T_40 : _GEN_14; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 244:36]
  wire [2:0] _GEN_24 = _T_83 ? _GEN_6 : _GEN_16; // @[Conditional.scala 39:67]
  wire  _GEN_25 = _T_75 | _GEN_17; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 224:36]
  wire [3:0] _GEN_28 = _T_75 ? _T_76 : _GEN_20; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 228:36]
  wire [63:0] _GEN_29 = _T_75 ? atomMemReg : io__wdata; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 229:36]
  wire  _GEN_30 = _T_75 ? _T_40 : _GEN_22; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 230:36]
  wire [2:0] _GEN_32 = _T_75 ? _GEN_6 : _GEN_24; // @[Conditional.scala 39:67]
  wire  _GEN_33 = _T_71 ? 1'h0 : _GEN_25; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 210:36]
  wire  _GEN_34 = _T_71 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 211:36]
  wire  _GEN_38 = _T_71 ? 1'h0 : _GEN_30; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 216:36]
  wire [2:0] _GEN_40 = _T_71 ? 3'h7 : _GEN_32; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 218:15]
  wire [63:0] _GEN_41 = _T_71 ? atomALU_io_result : atomMemReg; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 219:20 UnpipelinedLSU.scala 98:29]
  wire  _GEN_42 = _T_65 | _GEN_33; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 193:36]
  wire  _GEN_43 = _T_65 | _GEN_34; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 194:36]
  wire [3:0] _GEN_45 = _T_65 ? {{2'd0}, _T_66} : _GEN_28; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 197:36]
  wire  _GEN_47 = _T_65 ? 1'h0 : _GEN_38; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 199:36]
  wire [2:0] _GEN_49 = _T_65 ? _GEN_5 : _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_52 = _T_52 | _GEN_42; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 168:36]
  wire  _GEN_53 = _T_52 | _GEN_43; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 169:36]
  wire [6:0] _GEN_55 = _T_52 ? io__in_bits_func : {{3'd0}, _GEN_45}; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 172:36]
  wire [63:0] _GEN_56 = _T_52 ? io__wdata : _GEN_29; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 173:36]
  wire  _GEN_58 = _T_52 ? lsExecUnit_io__out_valid : _GEN_47; // @[Conditional.scala 39:67 UnpipelinedLSU.scala 175:36]
  wire  _GEN_68 = _T_29 ? lsExecUnit_io__out_valid | scInvalid | cannot_access_memory : _GEN_58; // @[Conditional.scala 40:58 UnpipelinedLSU.scala 157:38]
  wire [63:0] _T_109 = state == 3'h7 ? atomRegReg : lsExecUnit_io__out_bits; // @[UnpipelinedLSU.scala 284:45]
  wire  setLr = io__out_valid & (lrReq | scReq); // @[UnpipelinedLSU.scala 279:28]
  wire  setLrVal = lrReq; // @[UnpipelinedLSU.scala 57:25]
  wire [63:0] setLrAddr = io__in_bits_src1; // @[UnpipelinedLSU.scala 74:25 UnpipelinedLSU.scala 281:15]
  ysyx_210000_LSExecUnit lsExecUnit ( // @[UnpipelinedLSU.scala 48:28]
    .clock(lsExecUnit_clock),
    .reset(lsExecUnit_reset),
    .io__in_valid(lsExecUnit_io__in_valid),
    .io__in_bits_src1(lsExecUnit_io__in_bits_src1),
    .io__in_bits_func(lsExecUnit_io__in_bits_func),
    .io__out_ready(lsExecUnit_io__out_ready),
    .io__out_valid(lsExecUnit_io__out_valid),
    .io__out_bits(lsExecUnit_io__out_bits),
    .io__wdata(lsExecUnit_io__wdata),
    .io__dmem_req_ready(lsExecUnit_io__dmem_req_ready),
    .io__dmem_req_valid(lsExecUnit_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsExecUnit_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsExecUnit_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsExecUnit_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsExecUnit_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsExecUnit_io__dmem_req_bits_wdata),
    .io__dmem_resp_ready(lsExecUnit_io__dmem_resp_ready),
    .io__dmem_resp_valid(lsExecUnit_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsExecUnit_io__dmem_resp_bits_rdata),
    .io__isMMIO(lsExecUnit_io__isMMIO),
    .io__dtlbPF(lsExecUnit_io__dtlbPF),
    .io__loadAddrMisaligned(lsExecUnit_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsExecUnit_io__storeAddrMisaligned),
    .DTLBPF(lsExecUnit_DTLBPF),
    .DTLBENABLE(lsExecUnit_DTLBENABLE),
    .ISAMO2(lsExecUnit_ISAMO2),
    .io_in_bits_src1(lsExecUnit_io_in_bits_src1),
    .DTLBFINISH(lsExecUnit_DTLBFINISH)
  );
  ysyx_210000_AtomALU atomALU ( // @[UnpipelinedLSU.scala 100:25]
    .io_src1(atomALU_io_src1),
    .io_src2(atomALU_io_src2),
    .io_func(atomALU_io_func),
    .io_isWordOp(atomALU_io_isWordOp),
    .io_result(atomALU_io_result)
  );
  assign io__out_valid = DTLBPF | io__loadAddrMisaligned | io__storeAddrMisaligned | _GEN_68; // @[UnpipelinedLSU.scala 266:68 UnpipelinedLSU.scala 268:20]
  assign io__out_bits = scReq ? {{63'd0}, scInvalid} : _T_109; // @[UnpipelinedLSU.scala 284:23]
  assign io__dmem_req_valid = lsExecUnit_io__dmem_req_valid; // @[UnpipelinedLSU.scala 283:13]
  assign io__dmem_req_bits_addr = lsExecUnit_io__dmem_req_bits_addr; // @[UnpipelinedLSU.scala 283:13]
  assign io__dmem_req_bits_size = lsExecUnit_io__dmem_req_bits_size; // @[UnpipelinedLSU.scala 283:13]
  assign io__dmem_req_bits_cmd = lsExecUnit_io__dmem_req_bits_cmd; // @[UnpipelinedLSU.scala 283:13]
  assign io__dmem_req_bits_wmask = lsExecUnit_io__dmem_req_bits_wmask; // @[UnpipelinedLSU.scala 283:13]
  assign io__dmem_req_bits_wdata = lsExecUnit_io__dmem_req_bits_wdata; // @[UnpipelinedLSU.scala 283:13]
  assign io__dtlbPF = lsExecUnit_io__dtlbPF; // @[UnpipelinedLSU.scala 51:15]
  assign io__loadAddrMisaligned = lsExecUnit_io__loadAddrMisaligned; // @[UnpipelinedLSU.scala 294:27]
  assign io__storeAddrMisaligned = lsExecUnit_io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 295:28]
  assign setLr_0 = setLr;
  assign amoReq_0 = amoReq;
  assign io_in_bits_src1 = lsExecUnit_io_in_bits_src1;
  assign _T_20_0 = _T_20;
  assign setLrAddr_0 = _GEN_11;
  assign _T_28_0 = _T_28;
  assign setLrVal_0 = setLrVal;
  assign lsExecUnit_clock = clock;
  assign lsExecUnit_reset = reset;
  assign lsExecUnit_io__in_valid = _T_29 ? io__in_valid & ~atomReq & _T_34 : _GEN_52; // @[Conditional.scala 40:58 UnpipelinedLSU.scala 150:38]
  assign lsExecUnit_io__in_bits_src1 = _T_29 ? io__srcSum : io__in_bits_src1; // @[Conditional.scala 40:58 UnpipelinedLSU.scala 152:38]
  assign lsExecUnit_io__in_bits_func = _T_29 ? io__in_bits_func : _GEN_55; // @[Conditional.scala 40:58 UnpipelinedLSU.scala 154:38]
  assign lsExecUnit_io__out_ready = _T_29 | _GEN_53; // @[Conditional.scala 40:58 UnpipelinedLSU.scala 151:38]
  assign lsExecUnit_io__wdata = _T_29 ? io__wdata : _GEN_56; // @[Conditional.scala 40:58 UnpipelinedLSU.scala 155:38]
  assign lsExecUnit_io__dmem_req_ready = io__dmem_req_ready; // @[UnpipelinedLSU.scala 283:13]
  assign lsExecUnit_io__dmem_resp_valid = io__dmem_resp_valid; // @[UnpipelinedLSU.scala 283:13]
  assign lsExecUnit_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[UnpipelinedLSU.scala 283:13]
  assign lsExecUnit_DTLBPF = DTLBPF;
  assign lsExecUnit_DTLBENABLE = DTLBENABLE;
  assign lsExecUnit_ISAMO2 = amoReq;
  assign lsExecUnit_DTLBFINISH = DTLBFINISH;
  assign atomALU_io_src1 = atomMemReg; // @[UnpipelinedLSU.scala 101:21]
  assign atomALU_io_src2 = io__wdata; // @[UnpipelinedLSU.scala 102:21]
  assign atomALU_io_func = io__in_bits_func; // @[UnpipelinedLSU.scala 103:21]
  assign atomALU_io_isWordOp = ~funct3[0]; // @[UnpipelinedLSU.scala 68:22]
  always @(posedge clock) begin
    if (reset) begin // @[UnpipelinedLSU.scala 97:24]
      state <= 3'h0; // @[UnpipelinedLSU.scala 97:24]
    end else if (DTLBPF | io__loadAddrMisaligned | io__storeAddrMisaligned) begin // @[UnpipelinedLSU.scala 266:68]
      state <= 3'h0; // @[UnpipelinedLSU.scala 267:13]
    end else if (_T_29) begin // @[Conditional.scala 40:58]
      if (scReq & _T_34) begin // @[UnpipelinedLSU.scala 163:43]
        state <= _T_51; // @[UnpipelinedLSU.scala 163:50]
      end else begin
        state <= _GEN_2;
      end
    end else if (_T_52) begin // @[Conditional.scala 39:67]
      state <= _GEN_4;
    end else begin
      state <= _GEN_49;
    end
    if (reset) begin // @[UnpipelinedLSU.scala 98:29]
      atomMemReg <= 64'h0; // @[UnpipelinedLSU.scala 98:29]
    end else if (!(_T_29)) begin // @[Conditional.scala 40:58]
      if (!(_T_52)) begin // @[Conditional.scala 39:67]
        if (_T_65) begin // @[Conditional.scala 39:67]
          atomMemReg <= lsExecUnit_io__out_bits; // @[UnpipelinedLSU.scala 205:20]
        end else begin
          atomMemReg <= _GEN_41;
        end
      end
    end
    if (reset) begin // @[UnpipelinedLSU.scala 99:29]
      atomRegReg <= 64'h0; // @[UnpipelinedLSU.scala 99:29]
    end else if (!(_T_29)) begin // @[Conditional.scala 40:58]
      if (!(_T_52)) begin // @[Conditional.scala 39:67]
        if (_T_65) begin // @[Conditional.scala 39:67]
          atomRegReg <= lsExecUnit_io__out_bits; // @[UnpipelinedLSU.scala 206:20]
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_29 & _T_52 & ~(_T_36 | ~amoReq | ~lrReq | ~scReq | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at UnpipelinedLSU.scala:176 assert(!atomReq || !amoReq || !lrReq || !scReq)\n"); // @[UnpipelinedLSU.scala 176:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~_T_29 & _T_52 & ~(_T_36 | ~amoReq | ~lrReq | ~scReq | reset)) begin
          $fatal; // @[UnpipelinedLSU.scala 176:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  atomMemReg = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  atomRegReg = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_PipedMultiplier(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [64:0]  io_in_bits_0,
  input  [64:0]  io_in_bits_1,
  input          io_out_ready,
  output         io_out_valid,
  output [129:0] io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [64:0] REG; // @[PipedMultiplier.scala 25:43]
  reg [64:0] REG_1; // @[PipedMultiplier.scala 25:43]
  wire [129:0] mulRes = $signed(REG) * $signed(REG_1); // @[PipedMultiplier.scala 27:49]
  reg [129:0] REG_2; // @[PipedMultiplier.scala 26:44]
  wire  _T_4 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  reg  REG_3; // @[PipedMultiplier.scala 25:43]
  reg  REG_4; // @[PipedMultiplier.scala 26:44]
  reg  busy; // @[PipedMultiplier.scala 31:21]
  wire  _GEN_0 = io_in_valid & ~busy | busy; // @[PipedMultiplier.scala 32:31 PipedMultiplier.scala 32:38 PipedMultiplier.scala 31:21]
  assign io_in_ready = ~busy; // @[PipedMultiplier.scala 34:49]
  assign io_out_valid = REG_4; // @[PipedMultiplier.scala 29:16]
  assign io_out_bits = REG_2; // @[PipedMultiplier.scala 28:37]
  always @(posedge clock) begin
    if (reset) begin // @[PipedMultiplier.scala 25:43]
      REG <= 65'h0; // @[PipedMultiplier.scala 25:43]
    end else begin
      REG <= io_in_bits_0; // @[PipedMultiplier.scala 25:43]
    end
    if (reset) begin // @[PipedMultiplier.scala 25:43]
      REG_1 <= 65'h0; // @[PipedMultiplier.scala 25:43]
    end else begin
      REG_1 <= io_in_bits_1; // @[PipedMultiplier.scala 25:43]
    end
    if (reset) begin // @[PipedMultiplier.scala 26:44]
      REG_2 <= 130'sh0; // @[PipedMultiplier.scala 26:44]
    end else begin
      REG_2 <= mulRes; // @[PipedMultiplier.scala 26:44]
    end
    if (reset) begin // @[PipedMultiplier.scala 25:43]
      REG_3 <= 1'h0; // @[PipedMultiplier.scala 25:43]
    end else begin
      REG_3 <= _T_4; // @[PipedMultiplier.scala 25:43]
    end
    if (reset) begin // @[PipedMultiplier.scala 26:44]
      REG_4 <= 1'h0; // @[PipedMultiplier.scala 26:44]
    end else begin
      REG_4 <= REG_3; // @[PipedMultiplier.scala 26:44]
    end
    if (reset) begin // @[PipedMultiplier.scala 31:21]
      busy <= 1'h0; // @[PipedMultiplier.scala 31:21]
    end else if (io_out_valid) begin // @[PipedMultiplier.scala 33:23]
      busy <= 1'h0; // @[PipedMultiplier.scala 33:30]
    end else begin
      busy <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  REG = _RAND_0[64:0];
  _RAND_1 = {3{`RANDOM}};
  REG_1 = _RAND_1[64:0];
  _RAND_2 = {5{`RANDOM}};
  REG_2 = _RAND_2[129:0];
  _RAND_3 = {1{`RANDOM}};
  REG_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  busy = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_Radix4Divider(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [63:0]  io_in_bits_0,
  input  [63:0]  io_in_bits_1,
  input          io_sign,
  output         io_out_valid,
  output [127:0] io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [95:0] _RAND_8;
  reg [95:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Radix4Divider.scala 31:22]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  newReq = state == 3'h0 & _T_1; // @[Radix4Divider.scala 32:35]
  wire  _T_2 = state == 3'h2; // @[Radix4Divider.scala 34:48]
  wire  _T_3 = state == 3'h3; // @[Radix4Divider.scala 34:70]
  wire  _T_4 = state == 3'h2 | state == 3'h3; // @[Radix4Divider.scala 34:62]
  reg [5:0] cnt; // @[Reg.scala 27:20]
  reg [5:0] bLeadingZeros; // @[Reg.scala 27:20]
  wire [6:0] _T_280 = {1'h0,bLeadingZeros}; // @[Radix4Divider.scala 96:49]
  reg [5:0] aLeadingZeros; // @[Reg.scala 27:20]
  wire [6:0] _T_282 = {1'h0,aLeadingZeros}; // @[Radix4Divider.scala 96:89]
  wire [6:0] diff = $signed(_T_280) - $signed(_T_282); // @[Radix4Divider.scala 96:52]
  wire  isNegDiff = diff[6]; // @[Radix4Divider.scala 97:23]
  wire [6:0] _T_285 = $signed(_T_280) - $signed(_T_282); // @[Radix4Divider.scala 98:53]
  wire [6:0] quotientBits = isNegDiff ? 7'h0 : _T_285; // @[Radix4Divider.scala 98:25]
  wire [6:0] _T_315 = quotientBits + 7'h3; // @[Radix4Divider.scala 126:55]
  wire [5:0] _T_318 = cnt - 6'h1; // @[Radix4Divider.scala 126:72]
  wire [5:0] cnt_next = _T_2 ? _T_315[6:1] : _T_318; // @[Radix4Divider.scala 126:18]
  wire  rec_enough = cnt_next == 6'h0; // @[Radix4Divider.scala 35:29]
  wire  aSign = io_in_bits_0[63] & io_sign; // @[Radix4Divider.scala 38:24]
  wire [63:0] _T_7 = 64'h0 - io_in_bits_0; // @[Radix4Divider.scala 39:16]
  wire [63:0] aVal = aSign ? _T_7 : io_in_bits_0; // @[Radix4Divider.scala 39:12]
  wire  bSign = io_in_bits_1[63] & io_sign; // @[Radix4Divider.scala 38:24]
  wire [63:0] _T_10 = 64'h0 - io_in_bits_1; // @[Radix4Divider.scala 39:16]
  wire [63:0] bVal = bSign ? _T_10 : io_in_bits_1; // @[Radix4Divider.scala 39:12]
  reg  aSignReg; // @[Reg.scala 27:20]
  wire  _T_11 = aSign ^ bSign; // @[Radix4Divider.scala 45:34]
  reg  qSignReg; // @[Reg.scala 27:20]
  wire  divZero = io_in_bits_1 == 64'h0; // @[Radix4Divider.scala 46:19]
  reg  divZeroReg; // @[Reg.scala 27:20]
  wire  _T_12 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_15 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_17 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_5 = rec_enough ? 3'h4 : state; // @[Radix4Divider.scala 60:23 Radix4Divider.scala 60:31 Radix4Divider.scala 31:22]
  wire  _T_18 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_19 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_6 = io_out_valid ? 3'h0 : state; // @[Radix4Divider.scala 66:26 Radix4Divider.scala 66:34 Radix4Divider.scala 31:22]
  wire [2:0] _GEN_7 = _T_19 ? _GEN_6 : state; // @[Conditional.scala 39:67 Radix4Divider.scala 31:22]
  wire [2:0] _GEN_8 = _T_18 ? 3'h5 : _GEN_7; // @[Conditional.scala 39:67 Radix4Divider.scala 63:13]
  wire [2:0] _GEN_9 = _T_17 ? _GEN_5 : _GEN_8; // @[Conditional.scala 39:67]
  reg [67:0] ws; // @[Radix4Divider.scala 82:23]
  reg [67:0] wc; // @[Radix4Divider.scala 82:23]
  reg [67:0] d; // @[Radix4Divider.scala 84:18]
  wire [5:0] _T_86 = ws[1] ? 6'h3e : 6'h3f; // @[Mux.scala 47:69]
  wire [5:0] _T_87 = ws[2] ? 6'h3d : _T_86; // @[Mux.scala 47:69]
  wire [5:0] _T_88 = ws[3] ? 6'h3c : _T_87; // @[Mux.scala 47:69]
  wire [5:0] _T_89 = ws[4] ? 6'h3b : _T_88; // @[Mux.scala 47:69]
  wire [5:0] _T_90 = ws[5] ? 6'h3a : _T_89; // @[Mux.scala 47:69]
  wire [5:0] _T_91 = ws[6] ? 6'h39 : _T_90; // @[Mux.scala 47:69]
  wire [5:0] _T_92 = ws[7] ? 6'h38 : _T_91; // @[Mux.scala 47:69]
  wire [5:0] _T_93 = ws[8] ? 6'h37 : _T_92; // @[Mux.scala 47:69]
  wire [5:0] _T_94 = ws[9] ? 6'h36 : _T_93; // @[Mux.scala 47:69]
  wire [5:0] _T_95 = ws[10] ? 6'h35 : _T_94; // @[Mux.scala 47:69]
  wire [5:0] _T_96 = ws[11] ? 6'h34 : _T_95; // @[Mux.scala 47:69]
  wire [5:0] _T_97 = ws[12] ? 6'h33 : _T_96; // @[Mux.scala 47:69]
  wire [5:0] _T_98 = ws[13] ? 6'h32 : _T_97; // @[Mux.scala 47:69]
  wire [5:0] _T_99 = ws[14] ? 6'h31 : _T_98; // @[Mux.scala 47:69]
  wire [5:0] _T_100 = ws[15] ? 6'h30 : _T_99; // @[Mux.scala 47:69]
  wire [5:0] _T_101 = ws[16] ? 6'h2f : _T_100; // @[Mux.scala 47:69]
  wire [5:0] _T_102 = ws[17] ? 6'h2e : _T_101; // @[Mux.scala 47:69]
  wire [5:0] _T_103 = ws[18] ? 6'h2d : _T_102; // @[Mux.scala 47:69]
  wire [5:0] _T_104 = ws[19] ? 6'h2c : _T_103; // @[Mux.scala 47:69]
  wire [5:0] _T_105 = ws[20] ? 6'h2b : _T_104; // @[Mux.scala 47:69]
  wire [5:0] _T_106 = ws[21] ? 6'h2a : _T_105; // @[Mux.scala 47:69]
  wire [5:0] _T_107 = ws[22] ? 6'h29 : _T_106; // @[Mux.scala 47:69]
  wire [5:0] _T_108 = ws[23] ? 6'h28 : _T_107; // @[Mux.scala 47:69]
  wire [5:0] _T_109 = ws[24] ? 6'h27 : _T_108; // @[Mux.scala 47:69]
  wire [5:0] _T_110 = ws[25] ? 6'h26 : _T_109; // @[Mux.scala 47:69]
  wire [5:0] _T_111 = ws[26] ? 6'h25 : _T_110; // @[Mux.scala 47:69]
  wire [5:0] _T_112 = ws[27] ? 6'h24 : _T_111; // @[Mux.scala 47:69]
  wire [5:0] _T_113 = ws[28] ? 6'h23 : _T_112; // @[Mux.scala 47:69]
  wire [5:0] _T_114 = ws[29] ? 6'h22 : _T_113; // @[Mux.scala 47:69]
  wire [5:0] _T_115 = ws[30] ? 6'h21 : _T_114; // @[Mux.scala 47:69]
  wire [5:0] _T_116 = ws[31] ? 6'h20 : _T_115; // @[Mux.scala 47:69]
  wire [5:0] _T_117 = ws[32] ? 6'h1f : _T_116; // @[Mux.scala 47:69]
  wire [5:0] _T_118 = ws[33] ? 6'h1e : _T_117; // @[Mux.scala 47:69]
  wire [5:0] _T_119 = ws[34] ? 6'h1d : _T_118; // @[Mux.scala 47:69]
  wire [5:0] _T_120 = ws[35] ? 6'h1c : _T_119; // @[Mux.scala 47:69]
  wire [5:0] _T_121 = ws[36] ? 6'h1b : _T_120; // @[Mux.scala 47:69]
  wire [5:0] _T_122 = ws[37] ? 6'h1a : _T_121; // @[Mux.scala 47:69]
  wire [5:0] _T_123 = ws[38] ? 6'h19 : _T_122; // @[Mux.scala 47:69]
  wire [5:0] _T_124 = ws[39] ? 6'h18 : _T_123; // @[Mux.scala 47:69]
  wire [5:0] _T_125 = ws[40] ? 6'h17 : _T_124; // @[Mux.scala 47:69]
  wire [5:0] _T_126 = ws[41] ? 6'h16 : _T_125; // @[Mux.scala 47:69]
  wire [5:0] _T_127 = ws[42] ? 6'h15 : _T_126; // @[Mux.scala 47:69]
  wire [5:0] _T_128 = ws[43] ? 6'h14 : _T_127; // @[Mux.scala 47:69]
  wire [5:0] _T_129 = ws[44] ? 6'h13 : _T_128; // @[Mux.scala 47:69]
  wire [5:0] _T_130 = ws[45] ? 6'h12 : _T_129; // @[Mux.scala 47:69]
  wire [5:0] _T_131 = ws[46] ? 6'h11 : _T_130; // @[Mux.scala 47:69]
  wire [5:0] _T_132 = ws[47] ? 6'h10 : _T_131; // @[Mux.scala 47:69]
  wire [5:0] _T_133 = ws[48] ? 6'hf : _T_132; // @[Mux.scala 47:69]
  wire [5:0] _T_134 = ws[49] ? 6'he : _T_133; // @[Mux.scala 47:69]
  wire [5:0] _T_135 = ws[50] ? 6'hd : _T_134; // @[Mux.scala 47:69]
  wire [5:0] _T_136 = ws[51] ? 6'hc : _T_135; // @[Mux.scala 47:69]
  wire [5:0] _T_137 = ws[52] ? 6'hb : _T_136; // @[Mux.scala 47:69]
  wire [5:0] _T_138 = ws[53] ? 6'ha : _T_137; // @[Mux.scala 47:69]
  wire [5:0] _T_139 = ws[54] ? 6'h9 : _T_138; // @[Mux.scala 47:69]
  wire [5:0] _T_140 = ws[55] ? 6'h8 : _T_139; // @[Mux.scala 47:69]
  wire [5:0] _T_141 = ws[56] ? 6'h7 : _T_140; // @[Mux.scala 47:69]
  wire [5:0] _T_142 = ws[57] ? 6'h6 : _T_141; // @[Mux.scala 47:69]
  wire [5:0] _T_143 = ws[58] ? 6'h5 : _T_142; // @[Mux.scala 47:69]
  wire [5:0] _T_144 = ws[59] ? 6'h4 : _T_143; // @[Mux.scala 47:69]
  wire [5:0] _T_145 = ws[60] ? 6'h3 : _T_144; // @[Mux.scala 47:69]
  wire [5:0] _T_146 = ws[61] ? 6'h2 : _T_145; // @[Mux.scala 47:69]
  wire  _T_149 = state == 3'h1; // @[Radix4Divider.scala 89:19]
  wire [5:0] _T_215 = d[1] ? 6'h3e : 6'h3f; // @[Mux.scala 47:69]
  wire [5:0] _T_216 = d[2] ? 6'h3d : _T_215; // @[Mux.scala 47:69]
  wire [5:0] _T_217 = d[3] ? 6'h3c : _T_216; // @[Mux.scala 47:69]
  wire [5:0] _T_218 = d[4] ? 6'h3b : _T_217; // @[Mux.scala 47:69]
  wire [5:0] _T_219 = d[5] ? 6'h3a : _T_218; // @[Mux.scala 47:69]
  wire [5:0] _T_220 = d[6] ? 6'h39 : _T_219; // @[Mux.scala 47:69]
  wire [5:0] _T_221 = d[7] ? 6'h38 : _T_220; // @[Mux.scala 47:69]
  wire [5:0] _T_222 = d[8] ? 6'h37 : _T_221; // @[Mux.scala 47:69]
  wire [5:0] _T_223 = d[9] ? 6'h36 : _T_222; // @[Mux.scala 47:69]
  wire [5:0] _T_224 = d[10] ? 6'h35 : _T_223; // @[Mux.scala 47:69]
  wire [5:0] _T_225 = d[11] ? 6'h34 : _T_224; // @[Mux.scala 47:69]
  wire [5:0] _T_226 = d[12] ? 6'h33 : _T_225; // @[Mux.scala 47:69]
  wire [5:0] _T_227 = d[13] ? 6'h32 : _T_226; // @[Mux.scala 47:69]
  wire [5:0] _T_228 = d[14] ? 6'h31 : _T_227; // @[Mux.scala 47:69]
  wire [5:0] _T_229 = d[15] ? 6'h30 : _T_228; // @[Mux.scala 47:69]
  wire [5:0] _T_230 = d[16] ? 6'h2f : _T_229; // @[Mux.scala 47:69]
  wire [5:0] _T_231 = d[17] ? 6'h2e : _T_230; // @[Mux.scala 47:69]
  wire [5:0] _T_232 = d[18] ? 6'h2d : _T_231; // @[Mux.scala 47:69]
  wire [5:0] _T_233 = d[19] ? 6'h2c : _T_232; // @[Mux.scala 47:69]
  wire [5:0] _T_234 = d[20] ? 6'h2b : _T_233; // @[Mux.scala 47:69]
  wire [5:0] _T_235 = d[21] ? 6'h2a : _T_234; // @[Mux.scala 47:69]
  wire [5:0] _T_236 = d[22] ? 6'h29 : _T_235; // @[Mux.scala 47:69]
  wire [5:0] _T_237 = d[23] ? 6'h28 : _T_236; // @[Mux.scala 47:69]
  wire [5:0] _T_238 = d[24] ? 6'h27 : _T_237; // @[Mux.scala 47:69]
  wire [5:0] _T_239 = d[25] ? 6'h26 : _T_238; // @[Mux.scala 47:69]
  wire [5:0] _T_240 = d[26] ? 6'h25 : _T_239; // @[Mux.scala 47:69]
  wire [5:0] _T_241 = d[27] ? 6'h24 : _T_240; // @[Mux.scala 47:69]
  wire [5:0] _T_242 = d[28] ? 6'h23 : _T_241; // @[Mux.scala 47:69]
  wire [5:0] _T_243 = d[29] ? 6'h22 : _T_242; // @[Mux.scala 47:69]
  wire [5:0] _T_244 = d[30] ? 6'h21 : _T_243; // @[Mux.scala 47:69]
  wire [5:0] _T_245 = d[31] ? 6'h20 : _T_244; // @[Mux.scala 47:69]
  wire [5:0] _T_246 = d[32] ? 6'h1f : _T_245; // @[Mux.scala 47:69]
  wire [5:0] _T_247 = d[33] ? 6'h1e : _T_246; // @[Mux.scala 47:69]
  wire [5:0] _T_248 = d[34] ? 6'h1d : _T_247; // @[Mux.scala 47:69]
  wire [5:0] _T_249 = d[35] ? 6'h1c : _T_248; // @[Mux.scala 47:69]
  wire [5:0] _T_250 = d[36] ? 6'h1b : _T_249; // @[Mux.scala 47:69]
  wire [5:0] _T_251 = d[37] ? 6'h1a : _T_250; // @[Mux.scala 47:69]
  wire [5:0] _T_252 = d[38] ? 6'h19 : _T_251; // @[Mux.scala 47:69]
  wire [5:0] _T_253 = d[39] ? 6'h18 : _T_252; // @[Mux.scala 47:69]
  wire [5:0] _T_254 = d[40] ? 6'h17 : _T_253; // @[Mux.scala 47:69]
  wire [5:0] _T_255 = d[41] ? 6'h16 : _T_254; // @[Mux.scala 47:69]
  wire [5:0] _T_256 = d[42] ? 6'h15 : _T_255; // @[Mux.scala 47:69]
  wire [5:0] _T_257 = d[43] ? 6'h14 : _T_256; // @[Mux.scala 47:69]
  wire [5:0] _T_258 = d[44] ? 6'h13 : _T_257; // @[Mux.scala 47:69]
  wire [5:0] _T_259 = d[45] ? 6'h12 : _T_258; // @[Mux.scala 47:69]
  wire [5:0] _T_260 = d[46] ? 6'h11 : _T_259; // @[Mux.scala 47:69]
  wire [5:0] _T_261 = d[47] ? 6'h10 : _T_260; // @[Mux.scala 47:69]
  wire [5:0] _T_262 = d[48] ? 6'hf : _T_261; // @[Mux.scala 47:69]
  wire [5:0] _T_263 = d[49] ? 6'he : _T_262; // @[Mux.scala 47:69]
  wire [5:0] _T_264 = d[50] ? 6'hd : _T_263; // @[Mux.scala 47:69]
  wire [5:0] _T_265 = d[51] ? 6'hc : _T_264; // @[Mux.scala 47:69]
  wire [5:0] _T_266 = d[52] ? 6'hb : _T_265; // @[Mux.scala 47:69]
  wire [5:0] _T_267 = d[53] ? 6'ha : _T_266; // @[Mux.scala 47:69]
  wire [5:0] _T_268 = d[54] ? 6'h9 : _T_267; // @[Mux.scala 47:69]
  wire [5:0] _T_269 = d[55] ? 6'h8 : _T_268; // @[Mux.scala 47:69]
  wire [5:0] _T_270 = d[56] ? 6'h7 : _T_269; // @[Mux.scala 47:69]
  wire [5:0] _T_271 = d[57] ? 6'h6 : _T_270; // @[Mux.scala 47:69]
  wire [5:0] _T_272 = d[58] ? 6'h5 : _T_271; // @[Mux.scala 47:69]
  wire [5:0] _T_273 = d[59] ? 6'h4 : _T_272; // @[Mux.scala 47:69]
  wire [5:0] _T_274 = d[60] ? 6'h3 : _T_273; // @[Mux.scala 47:69]
  wire [5:0] _T_275 = d[61] ? 6'h2 : _T_274; // @[Mux.scala 47:69]
  wire  qBitsIsOdd = quotientBits[0]; // @[Radix4Divider.scala 99:32]
  wire [6:0] _GEN_30 = {{1'd0}, bLeadingZeros}; // @[Radix4Divider.scala 100:39]
  wire [6:0] _T_287 = 7'h40 - _GEN_30; // @[Radix4Divider.scala 100:39]
  reg [6:0] recoveryShift; // @[Reg.scala 27:20]
  wire [126:0] _GEN_31 = {{63'd0}, ws[63:0]}; // @[Radix4Divider.scala 103:18]
  wire [126:0] _T_290 = _GEN_31 << bLeadingZeros; // @[Radix4Divider.scala 103:18]
  wire [126:0] _T_292 = _GEN_31 << aLeadingZeros; // @[Radix4Divider.scala 104:18]
  wire [126:0] _T_293 = isNegDiff ? _T_290 : _T_292; // @[Radix4Divider.scala 102:19]
  wire [126:0] _GEN_33 = {{63'd0}, d[63:0]}; // @[Radix4Divider.scala 106:28]
  wire [126:0] _T_295 = _GEN_33 << bLeadingZeros; // @[Radix4Divider.scala 106:28]
  wire [67:0] rem_temp = ws + wc; // @[Radix4Divider.scala 108:21]
  wire [67:0] _T_299 = rem_temp + d; // @[Radix4Divider.scala 109:50]
  wire [67:0] rem_fixed = rem_temp[67] ? _T_299 : rem_temp; // @[Radix4Divider.scala 109:22]
  wire [194:0] _GEN_34 = {{127'd0}, rem_fixed}; // @[Radix4Divider.scala 110:28]
  wire [194:0] _T_300 = _GEN_34 << recoveryShift; // @[Radix4Divider.scala 110:28]
  wire [63:0] rem_abs = _T_300[128:65]; // @[Radix4Divider.scala 110:45]
  wire [63:0] lo = divZero ? io_in_bits_0 : aVal; // @[Radix4Divider.scala 113:28]
  wire [67:0] _T_301 = {4'h0,lo}; // @[Cat.scala 30:58]
  wire [67:0] _T_302 = {4'h0,bVal}; // @[Cat.scala 30:58]
  wire [63:0] b_shifted = _T_295[63:0]; // @[Radix4Divider.scala 101:34 Radix4Divider.scala 106:13]
  wire [67:0] _T_304 = {3'h0,b_shifted,1'h0}; // @[Cat.scala 30:58]
  wire [63:0] a_shifted = _T_293[63:0]; // @[Radix4Divider.scala 101:34 Radix4Divider.scala 102:13]
  wire [64:0] _T_305 = {a_shifted, 1'h0}; // @[Radix4Divider.scala 118:48]
  wire [64:0] _T_306 = qBitsIsOdd ? {{1'd0}, a_shifted} : _T_305; // @[Radix4Divider.scala 118:14]
  wire [65:0] hi_1 = wc[67:2]; // @[Radix4Divider.scala 183:22]
  wire [2:0] d_truncated = d[63:61]; // @[Radix4Divider.scala 146:22]
  wire [6:0] w_truncated = ws[67:61] + wc[67:61]; // @[Radix4Divider.scala 145:73]
  wire  _T_348 = $signed(w_truncated) >= 7'sh18; // @[Radix4Divider.scala 163:56]
  wire  _T_346 = $signed(w_truncated) >= 7'sh8; // @[Radix4Divider.scala 163:56]
  wire  _T_343 = $signed(w_truncated) >= -7'sh8; // @[Radix4Divider.scala 163:56]
  wire  _T_349 = $signed(w_truncated) >= -7'sh18; // @[Radix4Divider.scala 163:56]
  wire [2:0] _T_378 = _T_349 ? 3'h3 : 3'h4; // @[Mux.scala 98:16]
  wire [2:0] _T_379 = _T_343 ? 3'h0 : _T_378; // @[Mux.scala 98:16]
  wire [2:0] _T_380 = _T_346 ? 3'h1 : _T_379; // @[Mux.scala 98:16]
  wire [2:0] _T_381 = _T_348 ? 3'h2 : _T_380; // @[Mux.scala 98:16]
  wire  _T_345 = $signed(w_truncated) >= 7'sh14; // @[Radix4Divider.scala 163:56]
  wire  _T_347 = $signed(w_truncated) >= -7'sh16; // @[Radix4Divider.scala 163:56]
  wire [2:0] _T_374 = _T_347 ? 3'h3 : 3'h4; // @[Mux.scala 98:16]
  wire [2:0] _T_375 = _T_343 ? 3'h0 : _T_374; // @[Mux.scala 98:16]
  wire [2:0] _T_376 = _T_346 ? 3'h1 : _T_375; // @[Mux.scala 98:16]
  wire [2:0] _T_377 = _T_345 ? 3'h2 : _T_376; // @[Mux.scala 98:16]
  wire  _T_342 = $signed(w_truncated) >= 7'sh6; // @[Radix4Divider.scala 163:56]
  wire  _T_344 = $signed(w_truncated) >= -7'sh14; // @[Radix4Divider.scala 163:56]
  wire [2:0] _T_370 = _T_344 ? 3'h3 : 3'h4; // @[Mux.scala 98:16]
  wire [2:0] _T_371 = _T_343 ? 3'h0 : _T_370; // @[Mux.scala 98:16]
  wire [2:0] _T_372 = _T_342 ? 3'h1 : _T_371; // @[Mux.scala 98:16]
  wire [2:0] _T_373 = _T_345 ? 3'h2 : _T_372; // @[Mux.scala 98:16]
  wire  _T_341 = $signed(w_truncated) >= 7'sh12; // @[Radix4Divider.scala 163:56]
  wire [2:0] _T_369 = _T_341 ? 3'h2 : _T_372; // @[Mux.scala 98:16]
  wire  _T_339 = $signed(w_truncated) >= 7'sh10; // @[Radix4Divider.scala 163:56]
  wire  _T_331 = $signed(w_truncated) >= 7'sh4; // @[Radix4Divider.scala 163:56]
  wire  _T_335 = $signed(w_truncated) >= -7'sh6; // @[Radix4Divider.scala 163:56]
  wire  _T_340 = $signed(w_truncated) >= -7'sh12; // @[Radix4Divider.scala 163:56]
  wire [2:0] _T_362 = _T_340 ? 3'h3 : 3'h4; // @[Mux.scala 98:16]
  wire [2:0] _T_363 = _T_335 ? 3'h0 : _T_362; // @[Mux.scala 98:16]
  wire [2:0] _T_364 = _T_331 ? 3'h1 : _T_363; // @[Mux.scala 98:16]
  wire [2:0] _T_365 = _T_339 ? 3'h2 : _T_364; // @[Mux.scala 98:16]
  wire  _T_337 = $signed(w_truncated) >= 7'shf; // @[Radix4Divider.scala 163:56]
  wire  _T_338 = $signed(w_truncated) >= -7'sh10; // @[Radix4Divider.scala 163:56]
  wire [2:0] _T_358 = _T_338 ? 3'h3 : 3'h4; // @[Mux.scala 98:16]
  wire [2:0] _T_359 = _T_335 ? 3'h0 : _T_358; // @[Mux.scala 98:16]
  wire [2:0] _T_360 = _T_331 ? 3'h1 : _T_359; // @[Mux.scala 98:16]
  wire [2:0] _T_361 = _T_337 ? 3'h2 : _T_360; // @[Mux.scala 98:16]
  wire  _T_334 = $signed(w_truncated) >= 7'she; // @[Radix4Divider.scala 163:56]
  wire  _T_336 = $signed(w_truncated) >= -7'shf; // @[Radix4Divider.scala 163:56]
  wire [2:0] _T_354 = _T_336 ? 3'h3 : 3'h4; // @[Mux.scala 98:16]
  wire [2:0] _T_355 = _T_335 ? 3'h0 : _T_354; // @[Mux.scala 98:16]
  wire [2:0] _T_356 = _T_331 ? 3'h1 : _T_355; // @[Mux.scala 98:16]
  wire [2:0] _T_357 = _T_334 ? 3'h2 : _T_356; // @[Mux.scala 98:16]
  wire  _T_330 = $signed(w_truncated) >= 7'shc; // @[Radix4Divider.scala 163:56]
  wire  _T_332 = $signed(w_truncated) >= -7'sh4; // @[Radix4Divider.scala 163:56]
  wire  _T_333 = $signed(w_truncated) >= -7'shd; // @[Radix4Divider.scala 163:56]
  wire [2:0] _T_350 = _T_333 ? 3'h3 : 3'h4; // @[Mux.scala 98:16]
  wire [2:0] _T_351 = _T_332 ? 3'h0 : _T_350; // @[Mux.scala 98:16]
  wire [2:0] _T_352 = _T_331 ? 3'h1 : _T_351; // @[Mux.scala 98:16]
  wire [2:0] _T_353 = _T_330 ? 3'h2 : _T_352; // @[Mux.scala 98:16]
  wire [2:0] _T_383 = 3'h1 == d_truncated ? _T_357 : _T_353; // @[Mux.scala 80:57]
  wire [2:0] _T_385 = 3'h2 == d_truncated ? _T_361 : _T_383; // @[Mux.scala 80:57]
  wire [2:0] _T_387 = 3'h3 == d_truncated ? _T_365 : _T_385; // @[Mux.scala 80:57]
  wire [2:0] _T_389 = 3'h4 == d_truncated ? _T_369 : _T_387; // @[Mux.scala 80:57]
  wire [2:0] _T_391 = 3'h5 == d_truncated ? _T_373 : _T_389; // @[Mux.scala 80:57]
  wire [2:0] _T_393 = 3'h6 == d_truncated ? _T_377 : _T_391; // @[Mux.scala 80:57]
  wire [2:0] q_sel = 3'h7 == d_truncated ? _T_381 : _T_393; // @[Mux.scala 80:57]
  wire [1:0] _T_324 = 3'h1 == q_sel ? 2'h1 : 2'h0; // @[Mux.scala 80:57]
  wire [1:0] wc_adj = 3'h2 == q_sel ? 2'h2 : _T_324; // @[Mux.scala 80:57]
  wire [67:0] csa_in_1 = {hi_1,wc_adj}; // @[Cat.scala 30:58]
  wire [67:0] _T_405 = ws ^ csa_in_1; // @[CarrySaveAdder.scala 39:21]
  wire [68:0] _T_320 = {d, 1'h0}; // @[Radix4Divider.scala 135:12]
  wire [67:0] dx2 = _T_320[67:0]; // @[Radix4Divider.scala 134:33 Radix4Divider.scala 135:7]
  wire [67:0] neg_d = ~d; // @[Radix4Divider.scala 136:13]
  wire [68:0] _T_322 = {neg_d, 1'h0}; // @[Radix4Divider.scala 137:20]
  wire [67:0] neg_dx2 = _T_322[67:0]; // @[Radix4Divider.scala 134:33 Radix4Divider.scala 137:11]
  wire [67:0] _T_398 = 3'h1 == q_sel ? neg_d : 68'h0; // @[Mux.scala 80:57]
  wire [67:0] _T_400 = 3'h2 == q_sel ? neg_dx2 : _T_398; // @[Mux.scala 80:57]
  wire [67:0] _T_402 = 3'h3 == q_sel ? d : _T_400; // @[Mux.scala 80:57]
  wire [67:0] csa_in_2 = 3'h4 == q_sel ? dx2 : _T_402; // @[Mux.scala 80:57]
  wire [67:0] csa_out_0 = _T_405 ^ csa_in_2; // @[CarrySaveAdder.scala 41:23]
  wire [69:0] _T_308 = {csa_out_0, 2'h0}; // @[Radix4Divider.scala 120:44]
  wire [69:0] _T_309 = rec_enough ? {{2'd0}, csa_out_0} : _T_308; // @[Radix4Divider.scala 120:14]
  wire [67:0] _T_406 = ws & csa_in_1; // @[CarrySaveAdder.scala 40:21]
  wire [67:0] _T_407 = _T_405 & csa_in_2; // @[CarrySaveAdder.scala 42:35]
  wire [67:0] csa_out_1 = _T_406 | _T_407; // @[CarrySaveAdder.scala 42:24]
  wire [68:0] _T_408 = {csa_out_1, 1'h0}; // @[Radix4Divider.scala 192:25]
  wire [67:0] wc_next = _T_408[67:0]; // @[Radix4Divider.scala 83:30 Radix4Divider.scala 192:11]
  wire [69:0] _T_310 = {wc_next, 2'h0}; // @[Radix4Divider.scala 121:44]
  wire [69:0] _T_311 = rec_enough ? {{2'd0}, wc_next} : _T_310; // @[Radix4Divider.scala 121:14]
  wire  _T_312 = state == 3'h4; // @[Radix4Divider.scala 122:20]
  wire [67:0] _GEN_16 = state == 3'h4 ? {{4'd0}, rem_abs} : ws; // @[Radix4Divider.scala 122:35 Radix4Divider.scala 123:8 Radix4Divider.scala 82:23]
  wire [69:0] _GEN_17 = _T_3 ? _T_309 : {{2'd0}, _GEN_16}; // @[Radix4Divider.scala 119:37 Radix4Divider.scala 120:8]
  wire [69:0] _GEN_18 = _T_3 ? _T_311 : {{2'd0}, wc}; // @[Radix4Divider.scala 119:37 Radix4Divider.scala 121:8 Radix4Divider.scala 82:23]
  wire [69:0] _GEN_20 = _T_2 ? {{5'd0}, _T_306} : _GEN_17; // @[Radix4Divider.scala 116:35 Radix4Divider.scala 118:8]
  wire [69:0] _GEN_21 = _T_2 ? {{2'd0}, wc} : _GEN_18; // @[Radix4Divider.scala 116:35 Radix4Divider.scala 82:23]
  wire [69:0] _GEN_22 = newReq ? {{2'd0}, _T_301} : _GEN_20; // @[Radix4Divider.scala 112:15 Radix4Divider.scala 113:8]
  wire [69:0] _GEN_23 = newReq ? 70'h0 : _GEN_21; // @[Radix4Divider.scala 112:15 Radix4Divider.scala 114:8]
  reg [63:0] q; // @[Radix4Divider.scala 195:22]
  reg [63:0] qm; // @[Radix4Divider.scala 195:22]
  wire [61:0] hi_2 = q[61:0]; // @[Radix4Divider.scala 208:40]
  wire [63:0] _T_410 = {hi_2,2'h0}; // @[Cat.scala 30:58]
  wire [63:0] _T_411 = {hi_2,2'h1}; // @[Cat.scala 30:58]
  wire [63:0] _T_412 = {hi_2,2'h2}; // @[Cat.scala 30:58]
  wire [61:0] hi_5 = qm[61:0]; // @[Radix4Divider.scala 208:40]
  wire [63:0] _T_413 = {hi_5,2'h3}; // @[Cat.scala 30:58]
  wire [63:0] _T_414 = {hi_5,2'h2}; // @[Cat.scala 30:58]
  wire [63:0] _T_416 = 3'h0 == q_sel ? _T_410 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _T_418 = 3'h1 == q_sel ? _T_411 : _T_416; // @[Mux.scala 80:57]
  wire [63:0] _T_420 = 3'h2 == q_sel ? _T_412 : _T_418; // @[Mux.scala 80:57]
  wire [63:0] _T_422 = 3'h3 == q_sel ? _T_413 : _T_420; // @[Mux.scala 80:57]
  wire [63:0] _T_429 = {hi_5,2'h1}; // @[Cat.scala 30:58]
  wire [63:0] _T_431 = 3'h0 == q_sel ? _T_413 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _T_433 = 3'h1 == q_sel ? _T_410 : _T_431; // @[Mux.scala 80:57]
  wire [63:0] _T_435 = 3'h2 == q_sel ? _T_411 : _T_433; // @[Mux.scala 80:57]
  wire [63:0] _T_437 = 3'h3 == q_sel ? _T_414 : _T_435; // @[Mux.scala 80:57]
  wire [63:0] _T_442 = rem_temp[67] ? qm : q; // @[Radix4Divider.scala 221:13]
  wire [63:0] _T_445 = 64'h0 - ws[63:0]; // @[Radix4Divider.scala 225:33]
  wire [63:0] remainder = aSignReg ? _T_445 : ws[63:0]; // @[Radix4Divider.scala 225:22]
  wire [63:0] _T_448 = 64'h0 - q; // @[Radix4Divider.scala 226:32]
  wire [63:0] quotient = qSignReg ? _T_448 : q; // @[Radix4Divider.scala 226:21]
  wire [127:0] _T_451 = {ws[63:0],64'hffffffffffffffff}; // @[Cat.scala 30:58]
  wire [127:0] _T_452 = {remainder,quotient}; // @[Cat.scala 30:58]
  assign io_in_ready = state == 3'h0; // @[Radix4Divider.scala 227:23]
  assign io_out_valid = state == 3'h5; // @[Radix4Divider.scala 228:24]
  assign io_out_bits = divZeroReg ? _T_451 : _T_452; // @[Radix4Divider.scala 229:21]
  always @(posedge clock) begin
    if (reset) begin // @[Radix4Divider.scala 31:22]
      state <= 3'h0; // @[Radix4Divider.scala 31:22]
    end else if (_T_12) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Radix4Divider.scala 51:25]
        if (divZero) begin // @[Radix4Divider.scala 51:39]
          state <= 3'h5;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (_T_15) begin // @[Conditional.scala 39:67]
      state <= 3'h2; // @[Radix4Divider.scala 54:13]
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      state <= 3'h3; // @[Radix4Divider.scala 57:13]
    end else begin
      state <= _GEN_9;
    end
    if (reset) begin // @[Reg.scala 27:20]
      cnt <= 6'h0; // @[Reg.scala 27:20]
    end else if (_T_4) begin // @[Reg.scala 28:19]
      if (_T_2) begin // @[Radix4Divider.scala 126:18]
        cnt <= _T_315[6:1];
      end else begin
        cnt <= _T_318;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      bLeadingZeros <= 6'h0; // @[Reg.scala 27:20]
    end else if (_T_149) begin // @[Reg.scala 28:19]
      if (d[63]) begin // @[Mux.scala 47:69]
        bLeadingZeros <= 6'h0;
      end else if (d[62]) begin // @[Mux.scala 47:69]
        bLeadingZeros <= 6'h1;
      end else begin
        bLeadingZeros <= _T_275;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      aLeadingZeros <= 6'h0; // @[Reg.scala 27:20]
    end else if (_T_149) begin // @[Reg.scala 28:19]
      if (ws[63]) begin // @[Mux.scala 47:69]
        aLeadingZeros <= 6'h0;
      end else if (ws[62]) begin // @[Mux.scala 47:69]
        aLeadingZeros <= 6'h1;
      end else begin
        aLeadingZeros <= _T_146;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      aSignReg <= 1'h0; // @[Reg.scala 27:20]
    end else if (newReq) begin // @[Reg.scala 28:19]
      aSignReg <= aSign; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      qSignReg <= 1'h0; // @[Reg.scala 27:20]
    end else if (newReq) begin // @[Reg.scala 28:19]
      qSignReg <= _T_11; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      divZeroReg <= 1'h0; // @[Reg.scala 27:20]
    end else if (newReq) begin // @[Reg.scala 28:19]
      divZeroReg <= divZero; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Radix4Divider.scala 82:23]
      ws <= 68'h0; // @[Radix4Divider.scala 82:23]
    end else begin
      ws <= _GEN_22[67:0];
    end
    if (reset) begin // @[Radix4Divider.scala 82:23]
      wc <= 68'h0; // @[Radix4Divider.scala 82:23]
    end else begin
      wc <= _GEN_23[67:0];
    end
    if (reset) begin // @[Radix4Divider.scala 84:18]
      d <= 68'h0; // @[Radix4Divider.scala 84:18]
    end else if (newReq) begin // @[Radix4Divider.scala 112:15]
      d <= _T_302; // @[Radix4Divider.scala 115:7]
    end else if (_T_2) begin // @[Radix4Divider.scala 116:35]
      d <= _T_304; // @[Radix4Divider.scala 117:7]
    end
    if (reset) begin // @[Reg.scala 27:20]
      recoveryShift <= 7'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      recoveryShift <= _T_287; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Radix4Divider.scala 195:22]
      q <= 64'h0; // @[Radix4Divider.scala 195:22]
    end else if (newReq) begin // @[Radix4Divider.scala 196:15]
      q <= 64'h0; // @[Radix4Divider.scala 197:7]
    end else if (_T_3) begin // @[Radix4Divider.scala 199:37]
      if (3'h4 == q_sel) begin // @[Mux.scala 80:57]
        q <= _T_414;
      end else begin
        q <= _T_422;
      end
    end else if (_T_312) begin // @[Radix4Divider.scala 220:35]
      q <= _T_442; // @[Radix4Divider.scala 221:7]
    end
    if (reset) begin // @[Radix4Divider.scala 195:22]
      qm <= 64'h0; // @[Radix4Divider.scala 195:22]
    end else if (newReq) begin // @[Radix4Divider.scala 196:15]
      qm <= 64'h0; // @[Radix4Divider.scala 198:8]
    end else if (_T_3) begin // @[Radix4Divider.scala 199:37]
      if (3'h4 == q_sel) begin // @[Mux.scala 80:57]
        qm <= _T_429;
      end else begin
        qm <= _T_437;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  cnt = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  bLeadingZeros = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  aLeadingZeros = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  aSignReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  qSignReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  divZeroReg = _RAND_6[0:0];
  _RAND_7 = {3{`RANDOM}};
  ws = _RAND_7[67:0];
  _RAND_8 = {3{`RANDOM}};
  wc = _RAND_8[67:0];
  _RAND_9 = {3{`RANDOM}};
  d = _RAND_9[67:0];
  _RAND_10 = {1{`RANDOM}};
  recoveryShift = _RAND_10[6:0];
  _RAND_11 = {2{`RANDOM}};
  q = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  qm = _RAND_12[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_MDU(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  mul_clock; // @[MDU.scala 81:19]
  wire  mul_reset; // @[MDU.scala 81:19]
  wire  mul_io_in_ready; // @[MDU.scala 81:19]
  wire  mul_io_in_valid; // @[MDU.scala 81:19]
  wire [64:0] mul_io_in_bits_0; // @[MDU.scala 81:19]
  wire [64:0] mul_io_in_bits_1; // @[MDU.scala 81:19]
  wire  mul_io_out_ready; // @[MDU.scala 81:19]
  wire  mul_io_out_valid; // @[MDU.scala 81:19]
  wire [129:0] mul_io_out_bits; // @[MDU.scala 81:19]
  wire  div_clock; // @[MDU.scala 82:19]
  wire  div_reset; // @[MDU.scala 82:19]
  wire  div_io_in_ready; // @[MDU.scala 82:19]
  wire  div_io_in_valid; // @[MDU.scala 82:19]
  wire [63:0] div_io_in_bits_0; // @[MDU.scala 82:19]
  wire [63:0] div_io_in_bits_1; // @[MDU.scala 82:19]
  wire  div_io_sign; // @[MDU.scala 82:19]
  wire  div_io_out_valid; // @[MDU.scala 82:19]
  wire [127:0] div_io_out_bits; // @[MDU.scala 82:19]
  wire  isDiv = io_in_bits_func[2]; // @[MDU.scala 41:27]
  wire  isDivSign = isDiv & ~io_in_bits_func[0]; // @[MDU.scala 42:39]
  wire  isW = io_in_bits_func[3]; // @[MDU.scala 43:25]
  wire [64:0] _T_4 = {1'h0,io_in_bits_src1}; // @[Cat.scala 30:58]
  wire  hi = io_in_bits_src1[63]; // @[BitUtils.scala 39:20]
  wire [64:0] _T_5 = {hi,io_in_bits_src1}; // @[Cat.scala 30:58]
  wire  _T_8 = 2'h0 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_9 = 2'h1 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_10 = 2'h2 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_11 = 2'h3 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire [64:0] _T_12 = _T_8 ? _T_4 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_13 = _T_9 ? _T_5 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_14 = _T_10 ? _T_5 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_15 = _T_11 ? _T_4 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_16 = _T_12 | _T_13; // @[Mux.scala 27:72]
  wire [64:0] _T_17 = _T_16 | _T_14; // @[Mux.scala 27:72]
  wire [64:0] _T_20 = {1'h0,io_in_bits_src2}; // @[Cat.scala 30:58]
  wire  hi_2 = io_in_bits_src2[63]; // @[BitUtils.scala 39:20]
  wire [64:0] _T_21 = {hi_2,io_in_bits_src2}; // @[Cat.scala 30:58]
  wire [64:0] _T_28 = _T_8 ? _T_20 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_29 = _T_9 ? _T_21 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_30 = _T_10 ? _T_20 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_31 = _T_11 ? _T_20 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_32 = _T_28 | _T_29; // @[Mux.scala 27:72]
  wire [64:0] _T_33 = _T_32 | _T_30; // @[Mux.scala 27:72]
  wire [31:0] lo = io_in_bits_src1[31:0]; // @[MDU.scala 99:68]
  wire [31:0] hi_3 = lo[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_37 = {hi_3,lo}; // @[Cat.scala 30:58]
  wire [63:0] _T_38 = {32'h0,lo}; // @[Cat.scala 30:58]
  wire [63:0] _T_39 = isDivSign ? _T_37 : _T_38; // @[MDU.scala 99:47]
  wire [31:0] lo_2 = io_in_bits_src2[31:0]; // @[MDU.scala 99:68]
  wire [31:0] hi_4 = lo_2[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_43 = {hi_4,lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _T_44 = {32'h0,lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _T_45 = isDivSign ? _T_43 : _T_44; // @[MDU.scala 99:47]
  wire [63:0] mulRes = io_in_bits_func[1:0] == 2'h0 ? mul_io_out_bits[63:0] : mul_io_out_bits[127:64]; // @[MDU.scala 106:19]
  wire [63:0] divRes = io_in_bits_func[1] ? div_io_out_bits[127:64] : div_io_out_bits[63:0]; // @[MDU.scala 107:19]
  wire [63:0] res = isDiv ? divRes : mulRes; // @[MDU.scala 108:16]
  wire [31:0] lo_4 = res[31:0]; // @[MDU.scala 109:38]
  wire [31:0] hi_5 = lo_4[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_59 = {hi_5,lo_4}; // @[Cat.scala 30:58]
  wire  _T_61 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[MDU.scala 111:50]
  wire  isDivReg = _T_61 ? isDiv : REG; // @[MDU.scala 111:21]
  wire  _T_64 = mul_io_out_ready & mul_io_out_valid; // @[Decoupled.scala 40:37]
  ysyx_210000_PipedMultiplier mul ( // @[MDU.scala 81:19]
    .clock(mul_clock),
    .reset(mul_reset),
    .io_in_ready(mul_io_in_ready),
    .io_in_valid(mul_io_in_valid),
    .io_in_bits_0(mul_io_in_bits_0),
    .io_in_bits_1(mul_io_in_bits_1),
    .io_out_ready(mul_io_out_ready),
    .io_out_valid(mul_io_out_valid),
    .io_out_bits(mul_io_out_bits)
  );
  ysyx_210000_Radix4Divider div ( // @[MDU.scala 82:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_in_ready(div_io_in_ready),
    .io_in_valid(div_io_in_valid),
    .io_in_bits_0(div_io_in_bits_0),
    .io_in_bits_1(div_io_in_bits_1),
    .io_sign(div_io_sign),
    .io_out_valid(div_io_out_valid),
    .io_out_bits(div_io_out_bits)
  );
  assign io_in_ready = isDiv ? div_io_in_ready : mul_io_in_ready; // @[MDU.scala 112:21]
  assign io_out_valid = isDivReg ? div_io_out_valid : mul_io_out_valid; // @[MDU.scala 113:22]
  assign io_out_bits = isW ? _T_59 : res; // @[MDU.scala 109:21]
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_in_valid = io_in_valid & ~isDiv; // @[MDU.scala 103:34]
  assign mul_io_in_bits_0 = _T_17 | _T_15; // @[Mux.scala 27:72]
  assign mul_io_in_bits_1 = _T_33 | _T_31; // @[Mux.scala 27:72]
  assign mul_io_out_ready = 1'h1; // @[MDU.scala 85:17]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_in_valid = io_in_valid & isDiv; // @[MDU.scala 104:34]
  assign div_io_in_bits_0 = isW ? _T_39 : io_in_bits_src1; // @[MDU.scala 99:38]
  assign div_io_in_bits_1 = isW ? _T_45 : io_in_bits_src2; // @[MDU.scala 99:38]
  assign div_io_sign = isDiv & ~io_in_bits_func[0]; // @[MDU.scala 42:39]
  always @(posedge clock) begin
    if (reset) begin // @[MDU.scala 111:50]
      REG <= 1'h0; // @[MDU.scala 111:50]
    end else begin
      REG <= isDiv; // @[MDU.scala 111:50]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_CSR(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits,
  input  [63:0] io_cfIn_instr,
  input  [38:0] io_cfIn_pc,
  input         io_cfIn_exceptionVec_1,
  input         io_cfIn_exceptionVec_2,
  input         io_cfIn_exceptionVec_4,
  input         io_cfIn_exceptionVec_6,
  input         io_cfIn_exceptionVec_12,
  input         io_cfIn_intrVec_0,
  input         io_cfIn_intrVec_1,
  input         io_cfIn_intrVec_2,
  input         io_cfIn_intrVec_3,
  input         io_cfIn_intrVec_4,
  input         io_cfIn_intrVec_5,
  input         io_cfIn_intrVec_6,
  input         io_cfIn_intrVec_7,
  input         io_cfIn_intrVec_8,
  input         io_cfIn_intrVec_9,
  input         io_cfIn_intrVec_10,
  input         io_cfIn_intrVec_11,
  input         io_cfIn_crossPageIPFFix,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input         io_instrValid,
  input         io_lsuIsLoad,
  input         io_lsuPermitLibLoad,
  input         io_lsuPermitLibStore,
  output [1:0]  io_imemMMU_priviledgeMode,
  output [1:0]  io_dmemMMU_priviledgeMode,
  output        io_dmemMMU_status_sum,
  output        io_dmemMMU_status_mxr,
  input         io_dmemMMU_loadPF,
  input         io_dmemMMU_storePF,
  input  [38:0] io_dmemMMU_addr,
  output        io_wenFix,
  input         set_lr,
  input         is_pulpret,
  output [63:0] satp_0,
  input         perfCntCondMinstret,
  input         mtip_0,
  output        lsuDeny_0,
  input         meip_0,
  input         redirect_valid,
  input  [63:0] isu_addr,
  output        isuPermitLibLoad_0,
  output        isuPermitLibStore_0,
  input  [38:0] redirect_target,
  input  [63:0] LSUEXECADDR,
  output [11:0] intrVec_0,
  input         msip_0,
  input         lsu_is_valid,
  input  [63:0] set_lr_addr,
  input  [63:0] lsu_addr,
  input         perfCntCondMultiCommit,
  input         set_lr_val,
  output [63:0] lrAddr_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtvec; // @[CSR.scala 287:22]
  reg [63:0] mcounteren; // @[CSR.scala 288:27]
  reg [63:0] mcause; // @[CSR.scala 289:23]
  reg [63:0] mtval; // @[CSR.scala 290:22]
  reg [63:0] mepc; // @[CSR.scala 291:21]
  reg [63:0] mie; // @[CSR.scala 293:20]
  reg [63:0] mipReg; // @[CSR.scala 295:24]
  wire [11:0] _T_1 = {meip_0,1'h0,1'h0,1'h0,mtip_0,1'h0,2'h0,msip_0,3'h0}; // @[CSR.scala 297:22]
  wire [63:0] _GEN_195 = {{52'd0}, _T_1}; // @[CSR.scala 297:29]
  wire [63:0] _T_2 = _GEN_195 | mipReg; // @[CSR.scala 297:29]
  wire  mip_s_u = _T_2[0]; // @[CSR.scala 297:47]
  wire  mip_s_s = _T_2[1]; // @[CSR.scala 297:47]
  wire  mip_s_h = _T_2[2]; // @[CSR.scala 297:47]
  wire  mip_s_m = _T_2[3]; // @[CSR.scala 297:47]
  wire  mip_t_u = _T_2[4]; // @[CSR.scala 297:47]
  wire  mip_t_s = _T_2[5]; // @[CSR.scala 297:47]
  wire  mip_t_h = _T_2[6]; // @[CSR.scala 297:47]
  wire  mip_t_m = _T_2[7]; // @[CSR.scala 297:47]
  wire  mip_e_u = _T_2[8]; // @[CSR.scala 297:47]
  wire  mip_e_s = _T_2[9]; // @[CSR.scala 297:47]
  wire  mip_e_h = _T_2[10]; // @[CSR.scala 297:47]
  wire  mip_e_m = _T_2[11]; // @[CSR.scala 297:47]
  reg [63:0] misa; // @[CSR.scala 306:21]
  reg [63:0] mstatus; // @[CSR.scala 314:24]
  wire  mstatusStruct_ie_u = mstatus[0]; // @[CSR.scala 335:39]
  wire  mstatusStruct_ie_s = mstatus[1]; // @[CSR.scala 335:39]
  wire  mstatusStruct_ie_h = mstatus[2]; // @[CSR.scala 335:39]
  wire  mstatusStruct_ie_m = mstatus[3]; // @[CSR.scala 335:39]
  wire  mstatusStruct_pie_u = mstatus[4]; // @[CSR.scala 335:39]
  wire  mstatusStruct_pie_s = mstatus[5]; // @[CSR.scala 335:39]
  wire  mstatusStruct_pie_h = mstatus[6]; // @[CSR.scala 335:39]
  wire  mstatusStruct_pie_m = mstatus[7]; // @[CSR.scala 335:39]
  wire  mstatusStruct_spp = mstatus[8]; // @[CSR.scala 335:39]
  wire [1:0] mstatusStruct_hpp = mstatus[10:9]; // @[CSR.scala 335:39]
  wire [1:0] mstatusStruct_mpp = mstatus[12:11]; // @[CSR.scala 335:39]
  wire [1:0] mstatusStruct_fs = mstatus[14:13]; // @[CSR.scala 335:39]
  wire [1:0] mstatusStruct_xs = mstatus[16:15]; // @[CSR.scala 335:39]
  wire  mstatusStruct_mprv = mstatus[17]; // @[CSR.scala 335:39]
  wire  mstatusStruct_sum = mstatus[18]; // @[CSR.scala 335:39]
  wire  mstatusStruct_mxr = mstatus[19]; // @[CSR.scala 335:39]
  wire  mstatusStruct_tvm = mstatus[20]; // @[CSR.scala 335:39]
  wire  mstatusStruct_tw = mstatus[21]; // @[CSR.scala 335:39]
  wire  mstatusStruct_tsr = mstatus[22]; // @[CSR.scala 335:39]
  wire [8:0] mstatusStruct_pad0 = mstatus[31:23]; // @[CSR.scala 335:39]
  wire [1:0] mstatusStruct_uxl = mstatus[33:32]; // @[CSR.scala 335:39]
  wire [1:0] mstatusStruct_sxl = mstatus[35:34]; // @[CSR.scala 335:39]
  wire [26:0] mstatusStruct_pad1 = mstatus[62:36]; // @[CSR.scala 335:39]
  wire  mstatusStruct_sd = mstatus[63]; // @[CSR.scala 335:39]
  reg [63:0] medeleg; // @[CSR.scala 342:24]
  reg [63:0] mideleg; // @[CSR.scala 343:24]
  reg [63:0] mscratch; // @[CSR.scala 344:25]
  reg [63:0] pmpcfg0; // @[CSR.scala 346:24]
  reg [63:0] pmpcfg1; // @[CSR.scala 347:24]
  reg [63:0] pmpcfg2; // @[CSR.scala 348:24]
  reg [63:0] pmpcfg3; // @[CSR.scala 349:24]
  reg [63:0] pmpaddr0; // @[CSR.scala 350:25]
  reg [63:0] pmpaddr1; // @[CSR.scala 351:25]
  reg [63:0] pmpaddr2; // @[CSR.scala 352:25]
  reg [63:0] pmpaddr3; // @[CSR.scala 353:25]
  reg [63:0] dasicsSMainCfg; // @[CSR.scala 356:35]
  reg [63:0] dasicsSMainBoundHi; // @[CSR.scala 357:35]
  reg [63:0] dasicsSMainBoundLo; // @[CSR.scala 358:35]
  reg [63:0] stvec; // @[CSR.scala 378:22]
  wire [63:0] sieMask = 64'h222 & mideleg; // @[CSR.scala 380:26]
  reg [63:0] satp; // @[CSR.scala 383:21]
  reg [63:0] sepc; // @[CSR.scala 384:21]
  reg [63:0] scause; // @[CSR.scala 385:23]
  reg [63:0] stval; // @[CSR.scala 386:22]
  reg [63:0] sscratch; // @[CSR.scala 387:25]
  reg [63:0] scounteren; // @[CSR.scala 388:27]
  reg [63:0] sedeleg; // @[CSR.scala 390:24]
  reg [63:0] sideleg; // @[CSR.scala 391:24]
  reg [63:0] dasicsUMainCfg; // @[CSR.scala 394:35]
  reg [63:0] dasicsUMainBoundHi; // @[CSR.scala 395:35]
  reg [63:0] dasicsUMainBoundLo; // @[CSR.scala 396:35]
  wire [63:0] uieMask = 64'h111 & sideleg; // @[CSR.scala 411:26]
  reg [63:0] uepc; // @[CSR.scala 413:21]
  reg [63:0] ucause; // @[CSR.scala 414:23]
  reg [63:0] uscratch; // @[CSR.scala 415:25]
  reg [63:0] utvec; // @[CSR.scala 416:22]
  reg [63:0] utval; // @[CSR.scala 417:22]
  reg [63:0] dasicsLibBoundHiList_0; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_1; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_2; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_3; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_4; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_5; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_6; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_7; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_8; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_9; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_10; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_11; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_12; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_13; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_14; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundHiList_15; // @[CSR.scala 420:64]
  reg [63:0] dasicsLibBoundLoList_0; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_1; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_2; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_3; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_4; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_5; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_6; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_7; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_8; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_9; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_10; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_11; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_12; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_13; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_14; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibBoundLoList_15; // @[CSR.scala 421:64]
  reg [63:0] dasicsLibCfg0; // @[CSR.scala 425:31]
  reg [63:0] dasicsLibCfg1; // @[CSR.scala 426:31]
  reg [63:0] dasicsReturnPC; // @[CSR.scala 427:31]
  reg [63:0] dasicsFreeZoneReturnPC; // @[CSR.scala 428:39]
  reg [63:0] dasicsMaincallEntry; // @[CSR.scala 429:39]
  reg  lr; // @[CSR.scala 445:19]
  reg [63:0] lrAddr; // @[CSR.scala 446:23]
  reg [1:0] priviledgeMode; // @[CSR.scala 459:31]
  reg [63:0] perfCnts_0; // @[CSR.scala 464:47]
  reg [63:0] perfCnts_1; // @[CSR.scala 464:47]
  reg [63:0] perfCnts_2; // @[CSR.scala 464:47]
  wire [5:0] lo_2 = {mip_t_s,mip_t_u,mip_s_m,mip_s_h,mip_s_s,mip_s_u}; // @[CSR.scala 480:27]
  wire [11:0] _T_165 = {mip_e_m,mip_e_h,mip_e_s,mip_e_u,mip_t_m,mip_t_h,lo_2}; // @[CSR.scala 480:27]
  wire [11:0] addr = io_in_bits_src2[11:0]; // @[CSR.scala 548:18]
  wire [4:0] lo_5 = io_cfIn_instr[19:15]; // @[CSR.scala 550:35]
  wire [63:0] csri = {59'h0,lo_5}; // @[Cat.scala 30:58]
  wire  _T_397 = 12'h897 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_487 = _T_397 ? dasicsLibBoundHiList_10 : 64'h0; // @[Mux.scala 27:72]
  wire  _T_398 = 12'hbc0 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_488 = _T_398 ? dasicsSMainCfg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_577 = _T_487 | _T_488; // @[Mux.scala 27:72]
  wire  _T_399 = 12'h0 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_309 = mstatus & 64'h11; // @[RegMap.scala 48:84]
  wire [63:0] _T_489 = _T_399 ? _T_309 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_578 = _T_577 | _T_489; // @[Mux.scala 27:72]
  wire  _T_400 = 12'h8a2 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_490 = _T_400 ? dasicsLibBoundLoList_15 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_579 = _T_578 | _T_490; // @[Mux.scala 27:72]
  wire  _T_401 = 12'hf12 == addr; // @[LookupTree.scala 24:34]
  wire  _T_402 = 12'h5 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_492 = _T_402 ? utvec : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_581 = _T_579 | _T_492; // @[Mux.scala 27:72]
  wire  _T_403 = 12'h893 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_493 = _T_403 ? dasicsLibBoundHiList_8 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_582 = _T_581 | _T_493; // @[Mux.scala 27:72]
  wire  _T_404 = 12'h180 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_494 = _T_404 ? satp : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_583 = _T_582 | _T_494; // @[Mux.scala 27:72]
  wire  _T_405 = 12'h888 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_495 = _T_405 ? dasicsLibBoundLoList_2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_584 = _T_583 | _T_495; // @[Mux.scala 27:72]
  wire  _T_406 = 12'h3b1 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_496 = _T_406 ? pmpaddr1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_585 = _T_584 | _T_496; // @[Mux.scala 27:72]
  wire  _T_407 = 12'h3a2 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_497 = _T_407 ? pmpcfg2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_586 = _T_585 | _T_497; // @[Mux.scala 27:72]
  wire  _T_408 = 12'h140 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_498 = _T_408 ? sscratch : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_587 = _T_586 | _T_498; // @[Mux.scala 27:72]
  wire  _T_409 = 12'h889 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_499 = _T_409 ? dasicsLibBoundHiList_3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_588 = _T_587 | _T_499; // @[Mux.scala 27:72]
  wire  _T_410 = 12'h302 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_500 = _T_410 ? medeleg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_589 = _T_588 | _T_500; // @[Mux.scala 27:72]
  wire  _T_411 = 12'h105 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_501 = _T_411 ? stvec : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_590 = _T_589 | _T_501; // @[Mux.scala 27:72]
  wire  _T_412 = 12'h882 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_502 = _T_412 ? dasicsLibCfg1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_591 = _T_590 | _T_502; // @[Mux.scala 27:72]
  wire  _T_413 = 12'h141 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_503 = _T_413 ? sepc : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_592 = _T_591 | _T_503; // @[Mux.scala 27:72]
  wire  _T_414 = 12'h342 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_504 = _T_414 ? mcause : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_593 = _T_592 | _T_504; // @[Mux.scala 27:72]
  wire  _T_415 = 12'h88e == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_505 = _T_415 ? dasicsLibBoundLoList_5 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_594 = _T_593 | _T_505; // @[Mux.scala 27:72]
  wire  _T_416 = 12'h306 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_506 = _T_416 ? mcounteren : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_595 = _T_594 | _T_506; // @[Mux.scala 27:72]
  wire  _T_417 = 12'h89d == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_507 = _T_417 ? dasicsLibBoundHiList_13 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_596 = _T_595 | _T_507; // @[Mux.scala 27:72]
  wire  _T_418 = 12'hf11 == addr; // @[LookupTree.scala 24:34]
  wire  _T_419 = 12'h89c == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_509 = _T_419 ? dasicsLibBoundLoList_12 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_598 = _T_596 | _T_509; // @[Mux.scala 27:72]
  wire  _T_420 = 12'h104 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_330 = mie & sieMask; // @[RegMap.scala 48:84]
  wire [63:0] _T_510 = _T_420 ? _T_330 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_599 = _T_598 | _T_510; // @[Mux.scala 27:72]
  wire  _T_421 = 12'h41 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_511 = _T_421 ? uepc : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_600 = _T_599 | _T_511; // @[Mux.scala 27:72]
  wire  _T_422 = 12'h898 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_512 = _T_422 ? dasicsLibBoundLoList_10 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_601 = _T_600 | _T_512; // @[Mux.scala 27:72]
  wire  _T_423 = 12'h883 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_513 = _T_423 ? dasicsLibBoundHiList_0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_602 = _T_601 | _T_513; // @[Mux.scala 27:72]
  wire  _T_424 = 12'h885 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_514 = _T_424 ? dasicsLibBoundHiList_1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_603 = _T_602 | _T_514; // @[Mux.scala 27:72]
  wire  _T_425 = 12'h8a5 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_515 = _T_425 ? dasicsFreeZoneReturnPC : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_604 = _T_603 | _T_515; // @[Mux.scala 27:72]
  wire  _T_426 = 12'h8a3 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_516 = _T_426 ? dasicsMaincallEntry : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_605 = _T_604 | _T_516; // @[Mux.scala 27:72]
  wire  _T_427 = 12'h144 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _GEN_196 = {{52'd0}, _T_165}; // @[RegMap.scala 48:84]
  wire [63:0] _T_337 = _GEN_196 & sieMask; // @[RegMap.scala 48:84]
  wire [63:0] _T_517 = _T_427 ? _T_337 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_606 = _T_605 | _T_517; // @[Mux.scala 27:72]
  wire  _T_428 = 12'h100 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_338 = mstatus & 64'h80000003000de122; // @[RegMap.scala 48:84]
  wire [63:0] _T_518 = _T_428 ? _T_338 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_607 = _T_606 | _T_518; // @[Mux.scala 27:72]
  wire  _T_429 = 12'hbc2 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_519 = _T_429 ? dasicsSMainBoundLo : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_608 = _T_607 | _T_519; // @[Mux.scala 27:72]
  wire  _T_430 = 12'h894 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_520 = _T_430 ? dasicsLibBoundLoList_8 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_609 = _T_608 | _T_520; // @[Mux.scala 27:72]
  wire  _T_431 = 12'h89b == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_521 = _T_431 ? dasicsLibBoundHiList_12 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_610 = _T_609 | _T_521; // @[Mux.scala 27:72]
  wire  _T_432 = 12'h8a0 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_522 = _T_432 ? dasicsLibBoundLoList_14 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_611 = _T_610 | _T_522; // @[Mux.scala 27:72]
  wire  _T_433 = 12'h88d == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_523 = _T_433 ? dasicsLibBoundHiList_5 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_612 = _T_611 | _T_523; // @[Mux.scala 27:72]
  wire  _T_434 = 12'h305 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_524 = _T_434 ? mtvec : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_613 = _T_612 | _T_524; // @[Mux.scala 27:72]
  wire  _T_435 = 12'h40 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_525 = _T_435 ? uscratch : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_614 = _T_613 | _T_525; // @[Mux.scala 27:72]
  wire  _T_436 = 12'h88c == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_526 = _T_436 ? dasicsLibBoundLoList_4 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_615 = _T_614 | _T_526; // @[Mux.scala 27:72]
  wire  _T_437 = 12'h304 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_527 = _T_437 ? mie : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_616 = _T_615 | _T_527; // @[Mux.scala 27:72]
  wire  _T_438 = 12'hb01 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_528 = _T_438 ? perfCnts_1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_617 = _T_616 | _T_528; // @[Mux.scala 27:72]
  wire  _T_439 = 12'h103 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_529 = _T_439 ? sideleg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_618 = _T_617 | _T_529; // @[Mux.scala 27:72]
  wire  _T_440 = 12'h891 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_530 = _T_440 ? dasicsLibBoundHiList_7 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_619 = _T_618 | _T_530; // @[Mux.scala 27:72]
  wire  _T_441 = 12'h3b3 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_531 = _T_441 ? pmpaddr3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_620 = _T_619 | _T_531; // @[Mux.scala 27:72]
  wire  _T_442 = 12'h895 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_532 = _T_442 ? dasicsLibBoundHiList_9 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_621 = _T_620 | _T_532; // @[Mux.scala 27:72]
  wire  _T_443 = 12'h884 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_533 = _T_443 ? dasicsLibBoundLoList_0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_622 = _T_621 | _T_533; // @[Mux.scala 27:72]
  wire  _T_444 = 12'h886 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_534 = _T_444 ? dasicsLibBoundLoList_1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_623 = _T_622 | _T_534; // @[Mux.scala 27:72]
  wire  _T_445 = 12'h143 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_535 = _T_445 ? stval : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_624 = _T_623 | _T_535; // @[Mux.scala 27:72]
  wire  _T_446 = 12'h42 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_536 = _T_446 ? ucause : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_625 = _T_624 | _T_536; // @[Mux.scala 27:72]
  wire  _T_447 = 12'h301 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_537 = _T_447 ? misa : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_626 = _T_625 | _T_537; // @[Mux.scala 27:72]
  wire  _T_448 = 12'h5c2 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_538 = _T_448 ? dasicsUMainBoundLo : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_627 = _T_626 | _T_538; // @[Mux.scala 27:72]
  wire  _T_449 = 12'h8a4 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_539 = _T_449 ? dasicsReturnPC : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_628 = _T_627 | _T_539; // @[Mux.scala 27:72]
  wire  _T_450 = 12'h300 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_540 = _T_450 ? mstatus : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_629 = _T_628 | _T_540; // @[Mux.scala 27:72]
  wire  _T_451 = 12'h89f == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_541 = _T_451 ? dasicsLibBoundHiList_14 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_630 = _T_629 | _T_541; // @[Mux.scala 27:72]
  wire  _T_452 = 12'hbc1 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_542 = _T_452 ? dasicsSMainBoundHi : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_631 = _T_630 | _T_542; // @[Mux.scala 27:72]
  wire  _T_453 = 12'hb00 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_543 = _T_453 ? perfCnts_0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_632 = _T_631 | _T_543; // @[Mux.scala 27:72]
  wire  _T_454 = 12'h3b0 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_544 = _T_454 ? pmpaddr0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_633 = _T_632 | _T_544; // @[Mux.scala 27:72]
  wire  _T_455 = 12'h89a == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_545 = _T_455 ? dasicsLibBoundLoList_11 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_634 = _T_633 | _T_545; // @[Mux.scala 27:72]
  wire  _T_456 = 12'h5c0 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_546 = _T_456 ? dasicsUMainCfg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_635 = _T_634 | _T_546; // @[Mux.scala 27:72]
  wire  _T_457 = 12'h344 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_547 = _T_457 ? _GEN_196 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_636 = _T_635 | _T_547; // @[Mux.scala 27:72]
  wire  _T_458 = 12'h890 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_548 = _T_458 ? dasicsLibBoundLoList_6 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_637 = _T_636 | _T_548; // @[Mux.scala 27:72]
  wire  _T_459 = 12'h43 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_549 = _T_459 ? utval : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_638 = _T_637 | _T_549; // @[Mux.scala 27:72]
  wire  _T_460 = 12'hb02 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_550 = _T_460 ? perfCnts_2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_639 = _T_638 | _T_550; // @[Mux.scala 27:72]
  wire  _T_461 = 12'h3a3 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_551 = _T_461 ? pmpcfg3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_640 = _T_639 | _T_551; // @[Mux.scala 27:72]
  wire  _T_462 = 12'h892 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_552 = _T_462 ? dasicsLibBoundLoList_7 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_641 = _T_640 | _T_552; // @[Mux.scala 27:72]
  wire  _T_463 = 12'h8a1 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_553 = _T_463 ? dasicsLibBoundHiList_15 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_642 = _T_641 | _T_553; // @[Mux.scala 27:72]
  wire  _T_464 = 12'h88b == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_554 = _T_464 ? dasicsLibBoundHiList_4 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_643 = _T_642 | _T_554; // @[Mux.scala 27:72]
  wire  _T_465 = 12'h303 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_555 = _T_465 ? mideleg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_644 = _T_643 | _T_555; // @[Mux.scala 27:72]
  wire  _T_466 = 12'h3b2 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_556 = _T_466 ? pmpaddr2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_645 = _T_644 | _T_556; // @[Mux.scala 27:72]
  wire  _T_467 = 12'h102 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_557 = _T_467 ? sedeleg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_646 = _T_645 | _T_557; // @[Mux.scala 27:72]
  wire  _T_468 = 12'hf13 == addr; // @[LookupTree.scala 24:34]
  wire  _T_469 = 12'h3a1 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_559 = _T_469 ? pmpcfg1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_648 = _T_646 | _T_559; // @[Mux.scala 27:72]
  wire  _T_470 = 12'h896 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_560 = _T_470 ? dasicsLibBoundLoList_9 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_649 = _T_648 | _T_560; // @[Mux.scala 27:72]
  wire  _T_471 = 12'h887 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_561 = _T_471 ? dasicsLibBoundHiList_2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_650 = _T_649 | _T_561; // @[Mux.scala 27:72]
  wire  _T_472 = 12'h340 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_562 = _T_472 ? mscratch : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_651 = _T_650 | _T_562; // @[Mux.scala 27:72]
  wire  _T_473 = 12'hf14 == addr; // @[LookupTree.scala 24:34]
  wire  _T_474 = 12'h341 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_564 = _T_474 ? mepc : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_653 = _T_651 | _T_564; // @[Mux.scala 27:72]
  wire  _T_475 = 12'h343 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_565 = _T_475 ? mtval : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_654 = _T_653 | _T_565; // @[Mux.scala 27:72]
  wire  _T_476 = 12'h106 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_566 = _T_476 ? scounteren : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_655 = _T_654 | _T_566; // @[Mux.scala 27:72]
  wire  _T_477 = 12'h4 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_387 = mie & uieMask; // @[RegMap.scala 48:84]
  wire [63:0] _T_567 = _T_477 ? _T_387 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_656 = _T_655 | _T_567; // @[Mux.scala 27:72]
  wire  _T_478 = 12'h899 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_568 = _T_478 ? dasicsLibBoundHiList_11 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_657 = _T_656 | _T_568; // @[Mux.scala 27:72]
  wire  _T_479 = 12'h88a == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_569 = _T_479 ? dasicsLibBoundLoList_3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_658 = _T_657 | _T_569; // @[Mux.scala 27:72]
  wire  _T_480 = 12'h5c1 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_570 = _T_480 ? dasicsUMainBoundHi : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_659 = _T_658 | _T_570; // @[Mux.scala 27:72]
  wire  _T_481 = 12'h3a0 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_571 = _T_481 ? pmpcfg0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_660 = _T_659 | _T_571; // @[Mux.scala 27:72]
  wire  _T_482 = 12'h44 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_392 = _GEN_196 & uieMask; // @[RegMap.scala 48:84]
  wire [63:0] _T_572 = _T_482 ? _T_392 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_661 = _T_660 | _T_572; // @[Mux.scala 27:72]
  wire  _T_483 = 12'h142 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_573 = _T_483 ? scause : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_662 = _T_661 | _T_573; // @[Mux.scala 27:72]
  wire  _T_484 = 12'h89e == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_574 = _T_484 ? dasicsLibBoundLoList_13 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_663 = _T_662 | _T_574; // @[Mux.scala 27:72]
  wire  _T_485 = 12'h88f == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_575 = _T_485 ? dasicsLibBoundHiList_6 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_664 = _T_663 | _T_575; // @[Mux.scala 27:72]
  wire  _T_486 = 12'h881 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_576 = _T_486 ? dasicsLibCfg0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] rdata = _T_664 | _T_576; // @[Mux.scala 27:72]
  wire [63:0] _T_226 = rdata | io_in_bits_src1; // @[CSR.scala 553:30]
  wire [63:0] _T_227 = ~io_in_bits_src1; // @[CSR.scala 554:32]
  wire [63:0] _T_228 = rdata & _T_227; // @[CSR.scala 554:30]
  wire [63:0] _T_229 = rdata | csri; // @[CSR.scala 556:30]
  wire [63:0] _T_230 = ~csri; // @[CSR.scala 557:32]
  wire [63:0] _T_231 = rdata & _T_230; // @[CSR.scala 557:30]
  wire  _T_232 = 7'h1 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_233 = 7'h2 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_234 = 7'h3 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_235 = 7'h5 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_236 = 7'h6 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_237 = 7'h7 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire [63:0] _T_238 = _T_232 ? io_in_bits_src1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_239 = _T_233 ? _T_226 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_240 = _T_234 ? _T_228 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_241 = _T_235 ? csri : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_242 = _T_236 ? _T_229 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_243 = _T_237 ? _T_231 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_244 = _T_238 | _T_239; // @[Mux.scala 27:72]
  wire [63:0] _T_245 = _T_244 | _T_240; // @[Mux.scala 27:72]
  wire [63:0] _T_246 = _T_245 | _T_241; // @[Mux.scala 27:72]
  wire [63:0] _T_247 = _T_246 | _T_242; // @[Mux.scala 27:72]
  wire [63:0] wdata = _T_247 | _T_243; // @[Mux.scala 27:72]
  wire  satpLegalMode = wdata[63:60] == 4'h0 | wdata[63:60] == 4'h8; // @[CSR.scala 561:69]
  wire  isDasicsActive = dasicsSMainCfg[2]; // @[CSR.scala 566:38]
  wire  _T_258 = isDasicsActive & dasicsSMainCfg[1]; // @[CSR.scala 567:104]
  wire  isSMainEnable = _T_258 & dasicsSMainBoundLo <= dasicsSMainBoundHi; // @[CSR.scala 565:88]
  wire  _T_263 = isDasicsActive & dasicsUMainCfg[1]; // @[CSR.scala 568:104]
  wire  isUMainEnable = _T_263 & dasicsUMainBoundLo <= dasicsUMainBoundHi; // @[CSR.scala 565:88]
  wire  _T_267 = priviledgeMode == 2'h1; // @[CSR.scala 571:97]
  wire  _T_268 = priviledgeMode == 2'h1 & isSMainEnable; // @[CSR.scala 571:107]
  wire [63:0] _GEN_198 = {{25'd0}, io_cfIn_pc}; // @[CSR.scala 565:82]
  wire  _T_272 = _T_268 & _GEN_198 >= dasicsSMainBoundLo & _GEN_198 <= dasicsSMainBoundHi; // @[CSR.scala 565:88]
  wire  _T_273 = priviledgeMode == 2'h0; // @[CSR.scala 572:97]
  wire  _T_274 = priviledgeMode == 2'h0 & isUMainEnable; // @[CSR.scala 572:107]
  wire  _T_278 = _T_274 & _GEN_198 >= dasicsUMainBoundLo & _GEN_198 <= dasicsUMainBoundHi; // @[CSR.scala 565:88]
  wire  _T_282 = _T_272 | _T_267 & ~isSMainEnable; // @[CSR.scala 574:38]
  wire  _T_286 = _T_278 | _T_273 & ~isUMainEnable; // @[CSR.scala 575:38]
  wire  inTrustedZone = priviledgeMode > 2'h1 | _T_282 | _T_286; // @[CSR.scala 577:46]
  wire  wen = io_in_valid & io_in_bits_func != 7'h0 & (addr != 12'h180 | satpLegalMode); // @[CSR.scala 582:47]
  wire  isIllegalMode = priviledgeMode < addr[9:8] & inTrustedZone; // @[CSR.scala 583:51]
  wire  justRead = (io_in_bits_func == 7'h2 | io_in_bits_func == 7'h6) & io_in_bits_src1 == 64'h0; // @[CSR.scala 584:70]
  wire  isIllegalWrite = wen & addr[11:10] == 2'h3 & ~justRead; // @[CSR.scala 585:58]
  wire  isIllegalAccess = isIllegalMode | isIllegalWrite; // @[CSR.scala 586:39]
  wire  _T_306 = wen & ~isIllegalAccess; // @[CSR.scala 588:51]
  wire [63:0] _GEN_3 = _T_306 & addr == 12'hbc0 ? wdata : dasicsSMainCfg; // @[RegMap.scala 50:72 RegMap.scala 50:76 CSR.scala 356:35]
  wire  _T_678 = addr == 12'h0; // @[RegMap.scala 50:65]
  wire [63:0] _T_680 = wdata & 64'h11; // @[BitUtils.scala 32:13]
  wire [63:0] _T_682 = mstatus & 64'he; // @[BitUtils.scala 32:36]
  wire [63:0] _T_683 = _T_680 | _T_682; // @[BitUtils.scala 32:25]
  wire  hi_5 = _T_683[14:13] == 2'h3; // @[CSR.scala 338:40]
  wire [62:0] lo_6 = _T_683[62:0]; // @[CSR.scala 338:60]
  wire [63:0] _T_708 = {hi_5,lo_6}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_4 = _T_306 & addr == 12'h0 ? _T_708 : mstatus; // @[RegMap.scala 50:72 RegMap.scala 50:76 CSR.scala 314:24]
  wire  _T_727 = addr == 12'h180; // @[RegMap.scala 50:65]
  wire  _T_763 = addr == 12'h302; // @[RegMap.scala 50:65]
  wire [63:0] _T_765 = wdata & 64'h3fbbff; // @[BitUtils.scala 32:13]
  wire [63:0] _T_767 = medeleg & 64'h4400; // @[BitUtils.scala 32:36]
  wire [63:0] _T_768 = _T_765 | _T_767; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_17 = _T_306 & addr == 12'h141 ? wdata : sepc; // @[RegMap.scala 50:72 RegMap.scala 50:76 CSR.scala 384:21]
  wire [63:0] _GEN_18 = _T_306 & addr == 12'h342 ? wdata : mcause; // @[RegMap.scala 50:72 RegMap.scala 50:76 CSR.scala 289:23]
  wire [63:0] _T_819 = wdata & sieMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_820 = ~sieMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_821 = mie & _T_820; // @[BitUtils.scala 32:36]
  wire [63:0] _T_822 = _T_819 | _T_821; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_24 = _T_306 & addr == 12'h41 ? wdata : uepc; // @[RegMap.scala 50:72 RegMap.scala 50:76 CSR.scala 413:21]
  wire [63:0] _T_861 = wdata & 64'hc6122; // @[BitUtils.scala 32:13]
  wire [63:0] _T_863 = mstatus & 64'h39edd; // @[BitUtils.scala 32:36]
  wire [63:0] _T_864 = _T_861 | _T_863; // @[BitUtils.scala 32:25]
  wire  hi_6 = _T_864[14:13] == 2'h3; // @[CSR.scala 338:40]
  wire [62:0] lo_7 = _T_864[62:0]; // @[CSR.scala 338:60]
  wire [63:0] _T_889 = {hi_6,lo_7}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_30 = _T_306 & addr == 12'h100 ? _T_889 : _GEN_4; // @[RegMap.scala 50:72 RegMap.scala 50:76]
  wire [63:0] _GEN_47 = _T_306 & addr == 12'h143 ? wdata : stval; // @[RegMap.scala 50:72 RegMap.scala 50:76 CSR.scala 386:22]
  wire [63:0] _GEN_48 = _T_306 & addr == 12'h42 ? wdata : ucause; // @[RegMap.scala 50:72 RegMap.scala 50:76 CSR.scala 414:23]
  wire [63:0] _GEN_50 = _T_306 & addr == 12'h5c2 ? wdata : dasicsUMainBoundLo; // @[RegMap.scala 50:72 RegMap.scala 50:76 CSR.scala 396:35]
  wire  hi_7 = wdata[14:13] == 2'h3; // @[CSR.scala 338:40]
  wire [62:0] lo_8 = wdata[62:0]; // @[CSR.scala 338:60]
  wire [63:0] _T_1046 = {hi_7,lo_8}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_52 = _T_306 & addr == 12'h300 ? _T_1046 : _GEN_30; // @[RegMap.scala 50:72 RegMap.scala 50:76]
  wire [63:0] _GEN_60 = _T_306 & addr == 12'h43 ? wdata : utval; // @[RegMap.scala 50:72 RegMap.scala 50:76 CSR.scala 417:22]
  wire [63:0] _T_1127 = wdata & 64'h222; // @[BitUtils.scala 32:13]
  wire [63:0] _T_1129 = mideleg & 64'h1dd; // @[BitUtils.scala 32:36]
  wire [63:0] _T_1130 = _T_1127 | _T_1129; // @[BitUtils.scala 32:25]
  wire  _T_1137 = addr == 12'h102; // @[RegMap.scala 50:65]
  wire [63:0] _GEN_73 = _T_306 & addr == 12'h341 ? wdata : mepc; // @[RegMap.scala 50:72 RegMap.scala 50:76 CSR.scala 291:21]
  wire [63:0] _GEN_74 = _T_306 & addr == 12'h343 ? wdata : mtval; // @[RegMap.scala 50:72 RegMap.scala 50:76 CSR.scala 290:22]
  wire [63:0] _GEN_78 = _T_306 & addr == 12'h5c1 ? wdata : dasicsUMainBoundHi; // @[RegMap.scala 50:72 RegMap.scala 50:76 CSR.scala 395:35]
  wire [63:0] _GEN_80 = _T_306 & addr == 12'h142 ? wdata : scause; // @[RegMap.scala 50:72 RegMap.scala 50:76 CSR.scala 385:23]
  wire  _T_1234 = _T_397 ? 1'h0 : 1'h1; // @[Mux.scala 80:57]
  wire  _T_1236 = _T_398 ? 1'h0 : _T_1234; // @[Mux.scala 80:57]
  wire  _T_1238 = _T_399 ? 1'h0 : _T_1236; // @[Mux.scala 80:57]
  wire  _T_1240 = _T_400 ? 1'h0 : _T_1238; // @[Mux.scala 80:57]
  wire  _T_1242 = _T_401 ? 1'h0 : _T_1240; // @[Mux.scala 80:57]
  wire  _T_1244 = _T_402 ? 1'h0 : _T_1242; // @[Mux.scala 80:57]
  wire  _T_1246 = _T_403 ? 1'h0 : _T_1244; // @[Mux.scala 80:57]
  wire  _T_1248 = _T_404 ? 1'h0 : _T_1246; // @[Mux.scala 80:57]
  wire  _T_1250 = _T_405 ? 1'h0 : _T_1248; // @[Mux.scala 80:57]
  wire  _T_1252 = _T_406 ? 1'h0 : _T_1250; // @[Mux.scala 80:57]
  wire  _T_1254 = _T_407 ? 1'h0 : _T_1252; // @[Mux.scala 80:57]
  wire  _T_1256 = _T_408 ? 1'h0 : _T_1254; // @[Mux.scala 80:57]
  wire  _T_1258 = _T_409 ? 1'h0 : _T_1256; // @[Mux.scala 80:57]
  wire  _T_1260 = _T_410 ? 1'h0 : _T_1258; // @[Mux.scala 80:57]
  wire  _T_1262 = _T_411 ? 1'h0 : _T_1260; // @[Mux.scala 80:57]
  wire  _T_1264 = _T_412 ? 1'h0 : _T_1262; // @[Mux.scala 80:57]
  wire  _T_1266 = _T_413 ? 1'h0 : _T_1264; // @[Mux.scala 80:57]
  wire  _T_1268 = _T_414 ? 1'h0 : _T_1266; // @[Mux.scala 80:57]
  wire  _T_1270 = _T_415 ? 1'h0 : _T_1268; // @[Mux.scala 80:57]
  wire  _T_1272 = _T_416 ? 1'h0 : _T_1270; // @[Mux.scala 80:57]
  wire  _T_1274 = _T_417 ? 1'h0 : _T_1272; // @[Mux.scala 80:57]
  wire  _T_1276 = _T_418 ? 1'h0 : _T_1274; // @[Mux.scala 80:57]
  wire  _T_1278 = _T_419 ? 1'h0 : _T_1276; // @[Mux.scala 80:57]
  wire  _T_1280 = _T_420 ? 1'h0 : _T_1278; // @[Mux.scala 80:57]
  wire  _T_1282 = _T_421 ? 1'h0 : _T_1280; // @[Mux.scala 80:57]
  wire  _T_1284 = _T_422 ? 1'h0 : _T_1282; // @[Mux.scala 80:57]
  wire  _T_1286 = _T_423 ? 1'h0 : _T_1284; // @[Mux.scala 80:57]
  wire  _T_1288 = _T_424 ? 1'h0 : _T_1286; // @[Mux.scala 80:57]
  wire  _T_1290 = _T_425 ? 1'h0 : _T_1288; // @[Mux.scala 80:57]
  wire  _T_1292 = _T_426 ? 1'h0 : _T_1290; // @[Mux.scala 80:57]
  wire  _T_1294 = _T_427 ? 1'h0 : _T_1292; // @[Mux.scala 80:57]
  wire  _T_1296 = _T_428 ? 1'h0 : _T_1294; // @[Mux.scala 80:57]
  wire  _T_1298 = _T_429 ? 1'h0 : _T_1296; // @[Mux.scala 80:57]
  wire  _T_1300 = _T_430 ? 1'h0 : _T_1298; // @[Mux.scala 80:57]
  wire  _T_1302 = _T_431 ? 1'h0 : _T_1300; // @[Mux.scala 80:57]
  wire  _T_1304 = _T_432 ? 1'h0 : _T_1302; // @[Mux.scala 80:57]
  wire  _T_1306 = _T_433 ? 1'h0 : _T_1304; // @[Mux.scala 80:57]
  wire  _T_1308 = _T_434 ? 1'h0 : _T_1306; // @[Mux.scala 80:57]
  wire  _T_1310 = _T_435 ? 1'h0 : _T_1308; // @[Mux.scala 80:57]
  wire  _T_1312 = _T_436 ? 1'h0 : _T_1310; // @[Mux.scala 80:57]
  wire  _T_1314 = _T_437 ? 1'h0 : _T_1312; // @[Mux.scala 80:57]
  wire  _T_1316 = _T_438 ? 1'h0 : _T_1314; // @[Mux.scala 80:57]
  wire  _T_1318 = _T_439 ? 1'h0 : _T_1316; // @[Mux.scala 80:57]
  wire  _T_1320 = _T_440 ? 1'h0 : _T_1318; // @[Mux.scala 80:57]
  wire  _T_1322 = _T_441 ? 1'h0 : _T_1320; // @[Mux.scala 80:57]
  wire  _T_1324 = _T_442 ? 1'h0 : _T_1322; // @[Mux.scala 80:57]
  wire  _T_1326 = _T_443 ? 1'h0 : _T_1324; // @[Mux.scala 80:57]
  wire  _T_1328 = _T_444 ? 1'h0 : _T_1326; // @[Mux.scala 80:57]
  wire  _T_1330 = _T_445 ? 1'h0 : _T_1328; // @[Mux.scala 80:57]
  wire  _T_1332 = _T_446 ? 1'h0 : _T_1330; // @[Mux.scala 80:57]
  wire  _T_1334 = _T_447 ? 1'h0 : _T_1332; // @[Mux.scala 80:57]
  wire  _T_1336 = _T_448 ? 1'h0 : _T_1334; // @[Mux.scala 80:57]
  wire  _T_1338 = _T_449 ? 1'h0 : _T_1336; // @[Mux.scala 80:57]
  wire  _T_1340 = _T_450 ? 1'h0 : _T_1338; // @[Mux.scala 80:57]
  wire  _T_1342 = _T_451 ? 1'h0 : _T_1340; // @[Mux.scala 80:57]
  wire  _T_1344 = _T_452 ? 1'h0 : _T_1342; // @[Mux.scala 80:57]
  wire  _T_1346 = _T_453 ? 1'h0 : _T_1344; // @[Mux.scala 80:57]
  wire  _T_1348 = _T_454 ? 1'h0 : _T_1346; // @[Mux.scala 80:57]
  wire  _T_1350 = _T_455 ? 1'h0 : _T_1348; // @[Mux.scala 80:57]
  wire  _T_1352 = _T_456 ? 1'h0 : _T_1350; // @[Mux.scala 80:57]
  wire  _T_1354 = _T_457 ? 1'h0 : _T_1352; // @[Mux.scala 80:57]
  wire  _T_1356 = _T_458 ? 1'h0 : _T_1354; // @[Mux.scala 80:57]
  wire  _T_1358 = _T_459 ? 1'h0 : _T_1356; // @[Mux.scala 80:57]
  wire  _T_1360 = _T_460 ? 1'h0 : _T_1358; // @[Mux.scala 80:57]
  wire  _T_1362 = _T_461 ? 1'h0 : _T_1360; // @[Mux.scala 80:57]
  wire  _T_1364 = _T_462 ? 1'h0 : _T_1362; // @[Mux.scala 80:57]
  wire  _T_1366 = _T_463 ? 1'h0 : _T_1364; // @[Mux.scala 80:57]
  wire  _T_1368 = _T_464 ? 1'h0 : _T_1366; // @[Mux.scala 80:57]
  wire  _T_1370 = _T_465 ? 1'h0 : _T_1368; // @[Mux.scala 80:57]
  wire  _T_1372 = _T_466 ? 1'h0 : _T_1370; // @[Mux.scala 80:57]
  wire  _T_1374 = _T_467 ? 1'h0 : _T_1372; // @[Mux.scala 80:57]
  wire  _T_1376 = _T_468 ? 1'h0 : _T_1374; // @[Mux.scala 80:57]
  wire  _T_1378 = _T_469 ? 1'h0 : _T_1376; // @[Mux.scala 80:57]
  wire  _T_1380 = _T_470 ? 1'h0 : _T_1378; // @[Mux.scala 80:57]
  wire  _T_1382 = _T_471 ? 1'h0 : _T_1380; // @[Mux.scala 80:57]
  wire  _T_1384 = _T_472 ? 1'h0 : _T_1382; // @[Mux.scala 80:57]
  wire  _T_1386 = _T_473 ? 1'h0 : _T_1384; // @[Mux.scala 80:57]
  wire  _T_1388 = _T_474 ? 1'h0 : _T_1386; // @[Mux.scala 80:57]
  wire  _T_1390 = _T_475 ? 1'h0 : _T_1388; // @[Mux.scala 80:57]
  wire  _T_1392 = _T_476 ? 1'h0 : _T_1390; // @[Mux.scala 80:57]
  wire  _T_1394 = _T_477 ? 1'h0 : _T_1392; // @[Mux.scala 80:57]
  wire  _T_1396 = _T_478 ? 1'h0 : _T_1394; // @[Mux.scala 80:57]
  wire  _T_1398 = _T_479 ? 1'h0 : _T_1396; // @[Mux.scala 80:57]
  wire  _T_1400 = _T_480 ? 1'h0 : _T_1398; // @[Mux.scala 80:57]
  wire  _T_1402 = _T_481 ? 1'h0 : _T_1400; // @[Mux.scala 80:57]
  wire  _T_1404 = _T_482 ? 1'h0 : _T_1402; // @[Mux.scala 80:57]
  wire  _T_1406 = _T_483 ? 1'h0 : _T_1404; // @[Mux.scala 80:57]
  wire  _T_1408 = _T_484 ? 1'h0 : _T_1406; // @[Mux.scala 80:57]
  wire  _T_1410 = _T_485 ? 1'h0 : _T_1408; // @[Mux.scala 80:57]
  wire  isIllegalAddr = _T_486 ? 1'h0 : _T_1410; // @[Mux.scala 80:57]
  wire  resetSatp = _T_727 & wen; // @[CSR.scala 590:35]
  wire [63:0] _T_1444 = _T_457 ? mipReg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1441 = mipReg & sieMask; // @[RegMap.scala 48:84]
  wire [63:0] _T_1445 = _T_427 ? _T_1441 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] rdataFix = _T_1444 | _T_1445; // @[Mux.scala 27:72]
  wire [63:0] _T_1415 = rdataFix | io_in_bits_src1; // @[CSR.scala 601:33]
  wire [63:0] _T_1417 = rdataFix & _T_227; // @[CSR.scala 602:33]
  wire [63:0] _T_1418 = rdataFix | csri; // @[CSR.scala 604:33]
  wire [63:0] _T_1420 = rdataFix & _T_230; // @[CSR.scala 605:33]
  wire [63:0] _T_1428 = _T_233 ? _T_1415 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1429 = _T_234 ? _T_1417 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1431 = _T_236 ? _T_1418 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1432 = _T_237 ? _T_1420 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1433 = _T_238 | _T_1428; // @[Mux.scala 27:72]
  wire [63:0] _T_1434 = _T_1433 | _T_1429; // @[Mux.scala 27:72]
  wire [63:0] _T_1435 = _T_1434 | _T_241; // @[Mux.scala 27:72]
  wire [63:0] _T_1436 = _T_1435 | _T_1431; // @[Mux.scala 27:72]
  wire [63:0] wdataFix = _T_1436 | _T_1432; // @[Mux.scala 27:72]
  wire [63:0] _T_1449 = wdataFix & 64'h77f; // @[BitUtils.scala 32:13]
  wire [63:0] _T_1451 = mipReg & 64'h80; // @[BitUtils.scala 32:36]
  wire [63:0] _T_1452 = _T_1449 | _T_1451; // @[BitUtils.scala 32:25]
  wire [63:0] _T_1455 = wdataFix & sieMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_1457 = mipReg & _T_820; // @[BitUtils.scala 32:36]
  wire [63:0] _T_1458 = _T_1455 | _T_1457; // @[BitUtils.scala 32:25]
  wire  _T_1461 = dasicsSMainCfg[0] | dasicsUMainCfg[0]; // @[CSR.scala 610:34]
  wire [62:0] hi_8 = dasicsSMainCfg[63:1]; // @[CSR.scala 617:43]
  wire [63:0] _T_1463 = {hi_8,1'h0}; // @[Cat.scala 30:58]
  wire [62:0] hi_9 = dasicsUMainCfg[63:1]; // @[CSR.scala 625:41]
  wire [63:0] _T_1464 = {hi_9,1'h0}; // @[Cat.scala 30:58]
  wire  _T_1483 = dasicsLibCfg0[3] & dasicsLibCfg0[1]; // @[CSR.scala 647:123]
  wire  _T_1487 = _T_1483 & isu_addr >= dasicsLibBoundLoList_0 & isu_addr <= dasicsLibBoundHiList_0; // @[CSR.scala 565:88]
  wire  _T_1490 = dasicsLibCfg0[11] & dasicsLibCfg0[9]; // @[CSR.scala 647:123]
  wire  _T_1494 = _T_1490 & isu_addr >= dasicsLibBoundLoList_1 & isu_addr <= dasicsLibBoundHiList_1; // @[CSR.scala 565:88]
  wire  _T_1497 = dasicsLibCfg0[19] & dasicsLibCfg0[17]; // @[CSR.scala 647:123]
  wire  _T_1501 = _T_1497 & isu_addr >= dasicsLibBoundLoList_2 & isu_addr <= dasicsLibBoundHiList_2; // @[CSR.scala 565:88]
  wire  _T_1504 = dasicsLibCfg0[27] & dasicsLibCfg0[25]; // @[CSR.scala 647:123]
  wire  _T_1508 = _T_1504 & isu_addr >= dasicsLibBoundLoList_3 & isu_addr <= dasicsLibBoundHiList_3; // @[CSR.scala 565:88]
  wire  _T_1511 = dasicsLibCfg0[35] & dasicsLibCfg0[33]; // @[CSR.scala 647:123]
  wire  _T_1515 = _T_1511 & isu_addr >= dasicsLibBoundLoList_4 & isu_addr <= dasicsLibBoundHiList_4; // @[CSR.scala 565:88]
  wire  _T_1518 = dasicsLibCfg0[43] & dasicsLibCfg0[41]; // @[CSR.scala 647:123]
  wire  _T_1522 = _T_1518 & isu_addr >= dasicsLibBoundLoList_5 & isu_addr <= dasicsLibBoundHiList_5; // @[CSR.scala 565:88]
  wire  _T_1525 = dasicsLibCfg0[51] & dasicsLibCfg0[49]; // @[CSR.scala 647:123]
  wire  _T_1529 = _T_1525 & isu_addr >= dasicsLibBoundLoList_6 & isu_addr <= dasicsLibBoundHiList_6; // @[CSR.scala 565:88]
  wire  _T_1532 = dasicsLibCfg0[59] & dasicsLibCfg0[57]; // @[CSR.scala 647:123]
  wire  _T_1536 = _T_1532 & isu_addr >= dasicsLibBoundLoList_7 & isu_addr <= dasicsLibBoundHiList_7; // @[CSR.scala 565:88]
  wire  _T_1539 = dasicsLibCfg1[3] & dasicsLibCfg1[1]; // @[CSR.scala 647:123]
  wire  _T_1543 = _T_1539 & isu_addr >= dasicsLibBoundLoList_8 & isu_addr <= dasicsLibBoundHiList_8; // @[CSR.scala 565:88]
  wire  _T_1546 = dasicsLibCfg1[11] & dasicsLibCfg1[9]; // @[CSR.scala 647:123]
  wire  _T_1550 = _T_1546 & isu_addr >= dasicsLibBoundLoList_9 & isu_addr <= dasicsLibBoundHiList_9; // @[CSR.scala 565:88]
  wire  _T_1553 = dasicsLibCfg1[19] & dasicsLibCfg1[17]; // @[CSR.scala 647:123]
  wire  _T_1557 = _T_1553 & isu_addr >= dasicsLibBoundLoList_10 & isu_addr <= dasicsLibBoundHiList_10; // @[CSR.scala 565:88]
  wire  _T_1560 = dasicsLibCfg1[27] & dasicsLibCfg1[25]; // @[CSR.scala 647:123]
  wire  _T_1564 = _T_1560 & isu_addr >= dasicsLibBoundLoList_11 & isu_addr <= dasicsLibBoundHiList_11; // @[CSR.scala 565:88]
  wire  _T_1567 = dasicsLibCfg1[35] & dasicsLibCfg1[33]; // @[CSR.scala 647:123]
  wire  _T_1571 = _T_1567 & isu_addr >= dasicsLibBoundLoList_12 & isu_addr <= dasicsLibBoundHiList_12; // @[CSR.scala 565:88]
  wire  _T_1574 = dasicsLibCfg1[43] & dasicsLibCfg1[41]; // @[CSR.scala 647:123]
  wire  _T_1578 = _T_1574 & isu_addr >= dasicsLibBoundLoList_13 & isu_addr <= dasicsLibBoundHiList_13; // @[CSR.scala 565:88]
  wire  _T_1581 = dasicsLibCfg1[51] & dasicsLibCfg1[49]; // @[CSR.scala 647:123]
  wire  _T_1585 = _T_1581 & isu_addr >= dasicsLibBoundLoList_14 & isu_addr <= dasicsLibBoundHiList_14; // @[CSR.scala 565:88]
  wire  _T_1588 = dasicsLibCfg1[59] & dasicsLibCfg1[57]; // @[CSR.scala 647:123]
  wire  _T_1592 = _T_1588 & isu_addr >= dasicsLibBoundLoList_15 & isu_addr <= dasicsLibBoundHiList_15; // @[CSR.scala 565:88]
  wire  isuPermitLibLoad = inTrustedZone | (_T_1487 | (_T_1494 | (_T_1501 | (_T_1508 | (_T_1515 | (_T_1522 | (_T_1529 |
    (_T_1536 | (_T_1543 | (_T_1550 | (_T_1557 | (_T_1564 | (_T_1571 | (_T_1578 | (_T_1585 | _T_1592))))))))))))))); // @[CSR.scala 647:41]
  wire  _T_1611 = dasicsLibCfg0[3] & dasicsLibCfg0[0]; // @[CSR.scala 648:123]
  wire  _T_1615 = _T_1611 & isu_addr >= dasicsLibBoundLoList_0 & isu_addr <= dasicsLibBoundHiList_0; // @[CSR.scala 565:88]
  wire  _T_1618 = dasicsLibCfg0[11] & dasicsLibCfg0[8]; // @[CSR.scala 648:123]
  wire  _T_1622 = _T_1618 & isu_addr >= dasicsLibBoundLoList_1 & isu_addr <= dasicsLibBoundHiList_1; // @[CSR.scala 565:88]
  wire  _T_1625 = dasicsLibCfg0[19] & dasicsLibCfg0[16]; // @[CSR.scala 648:123]
  wire  _T_1629 = _T_1625 & isu_addr >= dasicsLibBoundLoList_2 & isu_addr <= dasicsLibBoundHiList_2; // @[CSR.scala 565:88]
  wire  _T_1632 = dasicsLibCfg0[27] & dasicsLibCfg0[24]; // @[CSR.scala 648:123]
  wire  _T_1636 = _T_1632 & isu_addr >= dasicsLibBoundLoList_3 & isu_addr <= dasicsLibBoundHiList_3; // @[CSR.scala 565:88]
  wire  _T_1639 = dasicsLibCfg0[35] & dasicsLibCfg0[32]; // @[CSR.scala 648:123]
  wire  _T_1643 = _T_1639 & isu_addr >= dasicsLibBoundLoList_4 & isu_addr <= dasicsLibBoundHiList_4; // @[CSR.scala 565:88]
  wire  _T_1646 = dasicsLibCfg0[43] & dasicsLibCfg0[40]; // @[CSR.scala 648:123]
  wire  _T_1650 = _T_1646 & isu_addr >= dasicsLibBoundLoList_5 & isu_addr <= dasicsLibBoundHiList_5; // @[CSR.scala 565:88]
  wire  _T_1653 = dasicsLibCfg0[51] & dasicsLibCfg0[48]; // @[CSR.scala 648:123]
  wire  _T_1657 = _T_1653 & isu_addr >= dasicsLibBoundLoList_6 & isu_addr <= dasicsLibBoundHiList_6; // @[CSR.scala 565:88]
  wire  _T_1660 = dasicsLibCfg0[59] & dasicsLibCfg0[56]; // @[CSR.scala 648:123]
  wire  _T_1664 = _T_1660 & isu_addr >= dasicsLibBoundLoList_7 & isu_addr <= dasicsLibBoundHiList_7; // @[CSR.scala 565:88]
  wire  _T_1667 = dasicsLibCfg1[3] & dasicsLibCfg1[0]; // @[CSR.scala 648:123]
  wire  _T_1671 = _T_1667 & isu_addr >= dasicsLibBoundLoList_8 & isu_addr <= dasicsLibBoundHiList_8; // @[CSR.scala 565:88]
  wire  _T_1674 = dasicsLibCfg1[11] & dasicsLibCfg1[8]; // @[CSR.scala 648:123]
  wire  _T_1678 = _T_1674 & isu_addr >= dasicsLibBoundLoList_9 & isu_addr <= dasicsLibBoundHiList_9; // @[CSR.scala 565:88]
  wire  _T_1681 = dasicsLibCfg1[19] & dasicsLibCfg1[16]; // @[CSR.scala 648:123]
  wire  _T_1685 = _T_1681 & isu_addr >= dasicsLibBoundLoList_10 & isu_addr <= dasicsLibBoundHiList_10; // @[CSR.scala 565:88]
  wire  _T_1688 = dasicsLibCfg1[27] & dasicsLibCfg1[24]; // @[CSR.scala 648:123]
  wire  _T_1692 = _T_1688 & isu_addr >= dasicsLibBoundLoList_11 & isu_addr <= dasicsLibBoundHiList_11; // @[CSR.scala 565:88]
  wire  _T_1695 = dasicsLibCfg1[35] & dasicsLibCfg1[32]; // @[CSR.scala 648:123]
  wire  _T_1699 = _T_1695 & isu_addr >= dasicsLibBoundLoList_12 & isu_addr <= dasicsLibBoundHiList_12; // @[CSR.scala 565:88]
  wire  _T_1702 = dasicsLibCfg1[43] & dasicsLibCfg1[40]; // @[CSR.scala 648:123]
  wire  _T_1706 = _T_1702 & isu_addr >= dasicsLibBoundLoList_13 & isu_addr <= dasicsLibBoundHiList_13; // @[CSR.scala 565:88]
  wire  _T_1709 = dasicsLibCfg1[51] & dasicsLibCfg1[48]; // @[CSR.scala 648:123]
  wire  _T_1713 = _T_1709 & isu_addr >= dasicsLibBoundLoList_14 & isu_addr <= dasicsLibBoundHiList_14; // @[CSR.scala 565:88]
  wire  _T_1716 = dasicsLibCfg1[59] & dasicsLibCfg1[56]; // @[CSR.scala 648:123]
  wire  _T_1720 = _T_1716 & isu_addr >= dasicsLibBoundLoList_15 & isu_addr <= dasicsLibBoundHiList_15; // @[CSR.scala 565:88]
  wire  isuPermitLibStore = inTrustedZone | (_T_1615 | (_T_1622 | (_T_1629 | (_T_1636 | (_T_1643 | (_T_1650 | (_T_1657
     | (_T_1664 | (_T_1671 | (_T_1678 | (_T_1685 | (_T_1692 | (_T_1699 | (_T_1706 | (_T_1713 | _T_1720))))))))))))))); // @[CSR.scala 648:41]
  wire  _T_1739 = ~io_lsuPermitLibLoad; // @[CSR.scala 656:74]
  wire  lsuSLibLoadDeny = io_lsuIsLoad & _T_267 & ~io_lsuPermitLibLoad; // @[CSR.scala 656:71]
  wire  lsuULibLoadDeny = io_lsuIsLoad & _T_273 & _T_1739; // @[CSR.scala 657:71]
  wire  _T_1743 = ~io_lsuIsLoad; // @[CSR.scala 658:32]
  wire  _T_1746 = ~io_lsuPermitLibStore; // @[CSR.scala 658:74]
  wire  lsuSLibStoreDeny = ~io_lsuIsLoad & _T_267 & ~io_lsuPermitLibStore; // @[CSR.scala 658:71]
  wire  lsuULibStoreDeny = _T_1743 & _T_273 & _T_1746; // @[CSR.scala 659:71]
  wire  lsuDeny = lsuSLibLoadDeny | lsuULibLoadDeny | lsuSLibStoreDeny | lsuULibStoreDeny; // @[CSR.scala 660:78]
  wire  lsuSLibLoadFault = lsu_is_valid & lsuSLibLoadDeny; // @[CSR.scala 663:38]
  wire  lsuULibLoadFault = lsu_is_valid & lsuULibLoadDeny; // @[CSR.scala 664:38]
  wire  lsuSLibStoreFault = lsu_is_valid & lsuSLibStoreDeny; // @[CSR.scala 665:38]
  wire  lsuULibStoreFault = lsu_is_valid & lsuULibStoreDeny; // @[CSR.scala 666:38]
  wire  _T_1753 = ~inTrustedZone; // @[CSR.scala 702:67]
  wire  _T_1756 = dasicsLibCfg0[3] & dasicsLibCfg0[2]; // @[CSR.scala 702:159]
  wire  _T_1760 = _T_1756 & _GEN_198 >= dasicsLibBoundLoList_0 & _GEN_198 <= dasicsLibBoundHiList_0; // @[CSR.scala 565:88]
  wire  _T_1763 = dasicsLibCfg0[11] & dasicsLibCfg0[10]; // @[CSR.scala 702:159]
  wire  _T_1767 = _T_1763 & _GEN_198 >= dasicsLibBoundLoList_1 & _GEN_198 <= dasicsLibBoundHiList_1; // @[CSR.scala 565:88]
  wire  _T_1770 = dasicsLibCfg0[19] & dasicsLibCfg0[18]; // @[CSR.scala 702:159]
  wire  _T_1774 = _T_1770 & _GEN_198 >= dasicsLibBoundLoList_2 & _GEN_198 <= dasicsLibBoundHiList_2; // @[CSR.scala 565:88]
  wire  _T_1777 = dasicsLibCfg0[27] & dasicsLibCfg0[26]; // @[CSR.scala 702:159]
  wire  _T_1781 = _T_1777 & _GEN_198 >= dasicsLibBoundLoList_3 & _GEN_198 <= dasicsLibBoundHiList_3; // @[CSR.scala 565:88]
  wire  _T_1784 = dasicsLibCfg0[35] & dasicsLibCfg0[34]; // @[CSR.scala 702:159]
  wire  _T_1788 = _T_1784 & _GEN_198 >= dasicsLibBoundLoList_4 & _GEN_198 <= dasicsLibBoundHiList_4; // @[CSR.scala 565:88]
  wire  _T_1791 = dasicsLibCfg0[43] & dasicsLibCfg0[42]; // @[CSR.scala 702:159]
  wire  _T_1795 = _T_1791 & _GEN_198 >= dasicsLibBoundLoList_5 & _GEN_198 <= dasicsLibBoundHiList_5; // @[CSR.scala 565:88]
  wire  _T_1798 = dasicsLibCfg0[51] & dasicsLibCfg0[50]; // @[CSR.scala 702:159]
  wire  _T_1802 = _T_1798 & _GEN_198 >= dasicsLibBoundLoList_6 & _GEN_198 <= dasicsLibBoundHiList_6; // @[CSR.scala 565:88]
  wire  _T_1805 = dasicsLibCfg0[59] & dasicsLibCfg0[58]; // @[CSR.scala 702:159]
  wire  _T_1809 = _T_1805 & _GEN_198 >= dasicsLibBoundLoList_7 & _GEN_198 <= dasicsLibBoundHiList_7; // @[CSR.scala 565:88]
  wire  _T_1812 = dasicsLibCfg1[3] & dasicsLibCfg1[2]; // @[CSR.scala 702:159]
  wire  _T_1816 = _T_1812 & _GEN_198 >= dasicsLibBoundLoList_8 & _GEN_198 <= dasicsLibBoundHiList_8; // @[CSR.scala 565:88]
  wire  _T_1819 = dasicsLibCfg1[11] & dasicsLibCfg1[10]; // @[CSR.scala 702:159]
  wire  _T_1823 = _T_1819 & _GEN_198 >= dasicsLibBoundLoList_9 & _GEN_198 <= dasicsLibBoundHiList_9; // @[CSR.scala 565:88]
  wire  _T_1826 = dasicsLibCfg1[19] & dasicsLibCfg1[18]; // @[CSR.scala 702:159]
  wire  _T_1830 = _T_1826 & _GEN_198 >= dasicsLibBoundLoList_10 & _GEN_198 <= dasicsLibBoundHiList_10; // @[CSR.scala 565:88]
  wire  _T_1833 = dasicsLibCfg1[27] & dasicsLibCfg1[26]; // @[CSR.scala 702:159]
  wire  _T_1837 = _T_1833 & _GEN_198 >= dasicsLibBoundLoList_11 & _GEN_198 <= dasicsLibBoundHiList_11; // @[CSR.scala 565:88]
  wire  _T_1840 = dasicsLibCfg1[35] & dasicsLibCfg1[34]; // @[CSR.scala 702:159]
  wire  _T_1844 = _T_1840 & _GEN_198 >= dasicsLibBoundLoList_12 & _GEN_198 <= dasicsLibBoundHiList_12; // @[CSR.scala 565:88]
  wire  _T_1847 = dasicsLibCfg1[43] & dasicsLibCfg1[42]; // @[CSR.scala 702:159]
  wire  _T_1851 = _T_1847 & _GEN_198 >= dasicsLibBoundLoList_13 & _GEN_198 <= dasicsLibBoundHiList_13; // @[CSR.scala 565:88]
  wire  _T_1854 = dasicsLibCfg1[51] & dasicsLibCfg1[50]; // @[CSR.scala 702:159]
  wire  _T_1858 = _T_1854 & _GEN_198 >= dasicsLibBoundLoList_14 & _GEN_198 <= dasicsLibBoundHiList_14; // @[CSR.scala 565:88]
  wire  _T_1861 = dasicsLibCfg1[59] & dasicsLibCfg1[58]; // @[CSR.scala 702:159]
  wire  _T_1865 = _T_1861 & _GEN_198 >= dasicsLibBoundLoList_15 & _GEN_198 <= dasicsLibBoundHiList_15; // @[CSR.scala 565:88]
  wire  inLibFreeZone = ~inTrustedZone & (_T_1760 | (_T_1767 | (_T_1774 | (_T_1781 | (_T_1788 | (_T_1795 | (_T_1802 | (
    _T_1809 | (_T_1816 | (_T_1823 | (_T_1830 | (_T_1837 | (_T_1844 | (_T_1851 | (_T_1858 | _T_1865))))))))))))))); // @[CSR.scala 702:80]
  wire [63:0] aluRedirectTarget = {{25'd0}, redirect_target};
  wire  _T_1887 = _T_268 & aluRedirectTarget >= dasicsSMainBoundLo & aluRedirectTarget <= dasicsSMainBoundHi; // @[CSR.scala 565:88]
  wire  _T_1893 = _T_274 & aluRedirectTarget >= dasicsUMainBoundLo & aluRedirectTarget <= dasicsUMainBoundHi; // @[CSR.scala 565:88]
  wire  _T_1897 = _T_1887 | _T_267 & ~isSMainEnable; // @[CSR.scala 574:38]
  wire  _T_1901 = _T_1893 | _T_273 & ~isUMainEnable; // @[CSR.scala 575:38]
  wire  targetInTrustedZone = priviledgeMode > 2'h1 | _T_1897 | _T_1901; // @[CSR.scala 577:46]
  wire  _T_1904 = ~targetInTrustedZone; // @[CSR.scala 702:67]
  wire  _T_1911 = _T_1756 & aluRedirectTarget >= dasicsLibBoundLoList_0 & aluRedirectTarget <= dasicsLibBoundHiList_0; // @[CSR.scala 565:88]
  wire  _T_1918 = _T_1763 & aluRedirectTarget >= dasicsLibBoundLoList_1 & aluRedirectTarget <= dasicsLibBoundHiList_1; // @[CSR.scala 565:88]
  wire  _T_1925 = _T_1770 & aluRedirectTarget >= dasicsLibBoundLoList_2 & aluRedirectTarget <= dasicsLibBoundHiList_2; // @[CSR.scala 565:88]
  wire  _T_1932 = _T_1777 & aluRedirectTarget >= dasicsLibBoundLoList_3 & aluRedirectTarget <= dasicsLibBoundHiList_3; // @[CSR.scala 565:88]
  wire  _T_1939 = _T_1784 & aluRedirectTarget >= dasicsLibBoundLoList_4 & aluRedirectTarget <= dasicsLibBoundHiList_4; // @[CSR.scala 565:88]
  wire  _T_1946 = _T_1791 & aluRedirectTarget >= dasicsLibBoundLoList_5 & aluRedirectTarget <= dasicsLibBoundHiList_5; // @[CSR.scala 565:88]
  wire  _T_1953 = _T_1798 & aluRedirectTarget >= dasicsLibBoundLoList_6 & aluRedirectTarget <= dasicsLibBoundHiList_6; // @[CSR.scala 565:88]
  wire  _T_1960 = _T_1805 & aluRedirectTarget >= dasicsLibBoundLoList_7 & aluRedirectTarget <= dasicsLibBoundHiList_7; // @[CSR.scala 565:88]
  wire  _T_1967 = _T_1812 & aluRedirectTarget >= dasicsLibBoundLoList_8 & aluRedirectTarget <= dasicsLibBoundHiList_8; // @[CSR.scala 565:88]
  wire  _T_1974 = _T_1819 & aluRedirectTarget >= dasicsLibBoundLoList_9 & aluRedirectTarget <= dasicsLibBoundHiList_9; // @[CSR.scala 565:88]
  wire  _T_1981 = _T_1826 & aluRedirectTarget >= dasicsLibBoundLoList_10 & aluRedirectTarget <= dasicsLibBoundHiList_10; // @[CSR.scala 565:88]
  wire  _T_1988 = _T_1833 & aluRedirectTarget >= dasicsLibBoundLoList_11 & aluRedirectTarget <= dasicsLibBoundHiList_11; // @[CSR.scala 565:88]
  wire  _T_1995 = _T_1840 & aluRedirectTarget >= dasicsLibBoundLoList_12 & aluRedirectTarget <= dasicsLibBoundHiList_12; // @[CSR.scala 565:88]
  wire  _T_2002 = _T_1847 & aluRedirectTarget >= dasicsLibBoundLoList_13 & aluRedirectTarget <= dasicsLibBoundHiList_13; // @[CSR.scala 565:88]
  wire  _T_2009 = _T_1854 & aluRedirectTarget >= dasicsLibBoundLoList_14 & aluRedirectTarget <= dasicsLibBoundHiList_14; // @[CSR.scala 565:88]
  wire  _T_2016 = _T_1861 & aluRedirectTarget >= dasicsLibBoundLoList_15 & aluRedirectTarget <= dasicsLibBoundHiList_15; // @[CSR.scala 565:88]
  wire  targetInLibFreeZone = ~targetInTrustedZone & (_T_1911 | (_T_1918 | (_T_1925 | (_T_1932 | (_T_1939 | (_T_1946 | (
    _T_1953 | (_T_1960 | (_T_1967 | (_T_1974 | (_T_1981 | (_T_1988 | (_T_1995 | (_T_2002 | (_T_2009 | _T_2016)))))))))))
    )))); // @[CSR.scala 702:80]
  wire  _T_2037 = redirect_valid & inTrustedZone & _T_1904 & ~is_pulpret; // @[CSR.scala 707:67]
  wire [38:0] _T_2039 = io_cfIn_pc + 39'h4; // @[CSR.scala 709:34]
  wire  _T_2044 = redirect_valid & _T_1753 & ~inLibFreeZone & targetInLibFreeZone; // @[CSR.scala 712:62]
  wire  _T_2054 = inTrustedZone | _T_1753 & targetInTrustedZone & (aluRedirectTarget == dasicsReturnPC |
    aluRedirectTarget == dasicsMaincallEntry) | targetInLibFreeZone; // @[CSR.scala 717:178]
  wire  aluPermitRedirect = _T_2054 | inLibFreeZone & _T_1904 & ~targetInLibFreeZone & aluRedirectTarget ==
    dasicsFreeZoneReturnPC; // @[CSR.scala 718:47]
  wire  _T_2064 = ~aluPermitRedirect; // @[CSR.scala 720:92]
  wire  aluSLibInstrFault = isSMainEnable & _T_267 & redirect_valid & ~aluPermitRedirect; // @[CSR.scala 720:89]
  wire  aluULibInstrFault = isUMainEnable & _T_273 & redirect_valid & _T_2064; // @[CSR.scala 721:89]
  wire  _T_2070 = io_in_bits_func == 7'h0; // @[CSR.scala 734:46]
  wire  isEbreak = addr == 12'h1 & io_in_bits_func == 7'h0; // @[CSR.scala 734:38]
  wire  isEcall = _T_678 & _T_2070; // @[CSR.scala 735:36]
  wire  isMret = _T_763 & _T_2070; // @[CSR.scala 736:36]
  wire  isSret = _T_1137 & _T_2070; // @[CSR.scala 737:36]
  wire  isUret = addr == 12'h2 & _T_2070; // @[CSR.scala 738:36]
  wire  hasInstrPageFault = io_cfIn_exceptionVec_12 & io_in_valid; // @[CSR.scala 795:63]
  wire  _T_2104 = aluSLibInstrFault | lsuSLibLoadFault | lsuSLibStoreFault; // @[CSR.scala 804:46]
  wire [63:0] _T_2109 = aluSLibInstrFault ? aluRedirectTarget : lsu_addr; // @[CSR.scala 806:17]
  wire [63:0] _GEN_129 = _T_2104 ? _T_2109 : _GEN_74; // @[CSR.scala 805:3 CSR.scala 806:11]
  wire  _T_2111 = hasInstrPageFault | io_dmemMMU_loadPF | io_dmemMMU_storePF; // @[CSR.scala 809:46]
  wire [38:0] lo_9 = io_cfIn_pc + 39'h2; // @[CSR.scala 810:88]
  wire [24:0] hi_10 = lo_9[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2116 = {hi_10,lo_9}; // @[Cat.scala 30:58]
  wire [24:0] hi_11 = io_cfIn_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2119 = {hi_11,io_cfIn_pc}; // @[Cat.scala 30:58]
  wire [63:0] _T_2120 = io_cfIn_crossPageIPFFix ? _T_2116 : _T_2119; // @[CSR.scala 810:42]
  wire [24:0] hi_12 = io_dmemMMU_addr[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2123 = {hi_12,io_dmemMMU_addr}; // @[Cat.scala 30:58]
  wire [63:0] _T_2124 = hasInstrPageFault ? _T_2120 : _T_2123; // @[CSR.scala 810:19]
  wire  _T_2125 = priviledgeMode == 2'h3; // @[CSR.scala 811:25]
  wire [63:0] _GEN_130 = priviledgeMode == 2'h3 ? _T_2124 : _GEN_129; // @[CSR.scala 811:35 CSR.scala 812:13]
  wire [63:0] _GEN_131 = priviledgeMode == 2'h3 ? _GEN_47 : _T_2124; // @[CSR.scala 811:35 CSR.scala 814:13]
  wire [63:0] _GEN_132 = hasInstrPageFault | io_dmemMMU_loadPF | io_dmemMMU_storePF ? _GEN_130 : _GEN_129; // @[CSR.scala 809:67]
  wire [63:0] _GEN_133 = hasInstrPageFault | io_dmemMMU_loadPF | io_dmemMMU_storePF ? _GEN_131 : _GEN_47; // @[CSR.scala 809:67]
  wire  _T_2134 = io_cfIn_exceptionVec_4 | io_cfIn_exceptionVec_6; // @[CSR.scala 819:30]
  wire [38:0] dmemAddrMisalignedAddr = LSUEXECADDR[38:0]; // @[CSR.scala 783:36 CSR.scala 801:28]
  wire [24:0] hi_14 = dmemAddrMisalignedAddr[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_2137 = {hi_14,dmemAddrMisalignedAddr}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_134 = _T_2134 ? _T_2137 : _GEN_132; // @[CSR.scala 820:3 CSR.scala 821:11]
  wire  _T_2147 = aluULibInstrFault | lsuULibLoadFault | lsuULibStoreFault; // @[CSR.scala 825:46]
  wire [63:0] _T_2152 = aluULibInstrFault ? aluRedirectTarget : lsu_addr; // @[CSR.scala 827:17]
  wire [63:0] _GEN_135 = _T_2147 ? _T_2152 : _GEN_60; // @[CSR.scala 826:3 CSR.scala 827:11]
  wire  mipRaiseIntr_e_s = mip_e_s | meip_0; // @[CSR.scala 849:31]
  wire [11:0] _T_2154 = {mip_e_m,mip_e_h,mipRaiseIntr_e_s,mip_e_u,mip_t_m,mip_t_h,lo_2}; // @[CSR.scala 851:41]
  wire [63:0] _GEN_234 = {{52'd0}, _T_2154}; // @[CSR.scala 851:26]
  wire [63:0] ideleg = mideleg & _GEN_234; // @[CSR.scala 851:26]
  wire  _T_2221 = priviledgeMode < 2'h1; // @[CSR.scala 852:125]
  wire  _T_2225 = priviledgeMode < 2'h3; // @[CSR.scala 853:106]
  wire  _T_2226 = _T_2125 & mstatusStruct_ie_m | priviledgeMode < 2'h3; // @[CSR.scala 853:87]
  wire  intrVecEnable_0 = ideleg[0] ? _T_267 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_2226; // @[CSR.scala 852:51]
  wire  intrVecEnable_1 = ideleg[1] ? _T_267 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_2226; // @[CSR.scala 852:51]
  wire  intrVecEnable_2 = ideleg[2] ? _T_267 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_2226; // @[CSR.scala 852:51]
  wire  intrVecEnable_3 = ideleg[3] ? _T_267 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_2226; // @[CSR.scala 852:51]
  wire  intrVecEnable_4 = ideleg[4] ? _T_267 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_2226; // @[CSR.scala 852:51]
  wire  intrVecEnable_5 = ideleg[5] ? _T_267 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_2226; // @[CSR.scala 852:51]
  wire  intrVecEnable_6 = ideleg[6] ? _T_267 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_2226; // @[CSR.scala 852:51]
  wire  intrVecEnable_7 = ideleg[7] ? _T_267 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_2226; // @[CSR.scala 852:51]
  wire  intrVecEnable_8 = ideleg[8] ? _T_267 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_2226; // @[CSR.scala 852:51]
  wire  intrVecEnable_9 = ideleg[9] ? _T_267 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_2226; // @[CSR.scala 852:51]
  wire  intrVecEnable_10 = ideleg[10] ? _T_267 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_2226; // @[CSR.scala 852:51]
  wire  intrVecEnable_11 = ideleg[11] ? _T_267 & mstatusStruct_ie_s | priviledgeMode < 2'h1 : _T_2226; // @[CSR.scala 852:51]
  wire [11:0] _T_2329 = mie[11:0] & _T_2154; // @[CSR.scala 857:27]
  wire [5:0] lo_13 = {intrVecEnable_5,intrVecEnable_4,intrVecEnable_3,intrVecEnable_2,intrVecEnable_1,intrVecEnable_0}; // @[CSR.scala 857:65]
  wire [11:0] _T_2330 = {intrVecEnable_11,intrVecEnable_10,intrVecEnable_9,intrVecEnable_8,intrVecEnable_7,
    intrVecEnable_6,lo_13}; // @[CSR.scala 857:65]
  wire [11:0] intrVec = _T_2329 & _T_2330; // @[CSR.scala 857:49]
  wire [2:0] _T_2331 = io_cfIn_intrVec_4 ? 3'h4 : 3'h0; // @[CSR.scala 861:69]
  wire [3:0] _T_2332 = io_cfIn_intrVec_8 ? 4'h8 : {{1'd0}, _T_2331}; // @[CSR.scala 861:69]
  wire [3:0] _T_2333 = io_cfIn_intrVec_0 ? 4'h0 : _T_2332; // @[CSR.scala 861:69]
  wire [3:0] _T_2334 = io_cfIn_intrVec_5 ? 4'h5 : _T_2333; // @[CSR.scala 861:69]
  wire [3:0] _T_2335 = io_cfIn_intrVec_9 ? 4'h9 : _T_2334; // @[CSR.scala 861:69]
  wire [3:0] _T_2336 = io_cfIn_intrVec_1 ? 4'h1 : _T_2335; // @[CSR.scala 861:69]
  wire [3:0] _T_2337 = io_cfIn_intrVec_7 ? 4'h7 : _T_2336; // @[CSR.scala 861:69]
  wire [3:0] _T_2338 = io_cfIn_intrVec_11 ? 4'hb : _T_2337; // @[CSR.scala 861:69]
  wire [3:0] intrNO = io_cfIn_intrVec_3 ? 4'h3 : _T_2338; // @[CSR.scala 861:69]
  wire [5:0] lo_14 = {io_cfIn_intrVec_5,io_cfIn_intrVec_4,io_cfIn_intrVec_3,io_cfIn_intrVec_2,io_cfIn_intrVec_1,
    io_cfIn_intrVec_0}; // @[CSR.scala 863:35]
  wire [11:0] _T_2339 = {io_cfIn_intrVec_11,io_cfIn_intrVec_10,io_cfIn_intrVec_9,io_cfIn_intrVec_8,io_cfIn_intrVec_7,
    io_cfIn_intrVec_6,lo_14}; // @[CSR.scala 863:35]
  wire  raiseIntr = |_T_2339; // @[CSR.scala 863:42]
  wire  csrExceptionVec_3 = io_in_valid & isEbreak; // @[CSR.scala 870:46]
  wire  csrExceptionVec_11 = _T_2125 & io_in_valid & isEcall; // @[CSR.scala 871:70]
  wire  csrExceptionVec_9 = _T_267 & io_in_valid & isEcall; // @[CSR.scala 872:70]
  wire  csrExceptionVec_8 = _T_273 & io_in_valid & isEcall; // @[CSR.scala 873:70]
  wire  csrExceptionVec_2 = (isIllegalAddr | isIllegalAccess) & wen; // @[CSR.scala 874:71]
  wire [10:0] lo_15 = {1'h0,csrExceptionVec_9,csrExceptionVec_8,3'h0,1'h0,csrExceptionVec_3,csrExceptionVec_2,2'h0}; // @[CSR.scala 884:49]
  wire [4:0] hi_lo_9 = {io_dmemMMU_storePF,1'h0,io_dmemMMU_loadPF,1'h0,csrExceptionVec_11}; // @[CSR.scala 884:49]
  wire [21:0] _T_2354 = {lsuSLibStoreFault,lsuULibStoreFault,lsuSLibLoadFault,lsuULibLoadFault,aluSLibInstrFault,
    aluULibInstrFault,hi_lo_9,lo_15}; // @[CSR.scala 884:49]
  wire [10:0] lo_16 = {3'h0,1'h0,io_cfIn_exceptionVec_6,1'h0,io_cfIn_exceptionVec_4,1'h0,io_cfIn_exceptionVec_2,
    io_cfIn_exceptionVec_1,1'h0}; // @[CSR.scala 884:76]
  wire [21:0] _T_2355 = {6'h0,3'h0,io_cfIn_exceptionVec_12,1'h0,lo_16}; // @[CSR.scala 884:76]
  wire [21:0] raiseExceptionVec = _T_2354 | _T_2355; // @[CSR.scala 884:52]
  wire  raiseException = |raiseExceptionVec; // @[CSR.scala 885:42]
  wire [4:0] _T_2357 = raiseExceptionVec[20] ? 5'h14 : 5'h0; // @[CSR.scala 886:74]
  wire [4:0] _T_2359 = raiseExceptionVec[18] ? 5'h12 : _T_2357; // @[CSR.scala 886:74]
  wire [4:0] _T_2361 = raiseExceptionVec[16] ? 5'h10 : _T_2359; // @[CSR.scala 886:74]
  wire [4:0] _T_2363 = raiseExceptionVec[21] ? 5'h15 : _T_2361; // @[CSR.scala 886:74]
  wire [4:0] _T_2365 = raiseExceptionVec[19] ? 5'h13 : _T_2363; // @[CSR.scala 886:74]
  wire [4:0] _T_2367 = raiseExceptionVec[17] ? 5'h11 : _T_2365; // @[CSR.scala 886:74]
  wire [4:0] _T_2369 = raiseExceptionVec[5] ? 5'h5 : _T_2367; // @[CSR.scala 886:74]
  wire [4:0] _T_2371 = raiseExceptionVec[7] ? 5'h7 : _T_2369; // @[CSR.scala 886:74]
  wire [4:0] _T_2373 = raiseExceptionVec[13] ? 5'hd : _T_2371; // @[CSR.scala 886:74]
  wire [4:0] _T_2375 = raiseExceptionVec[15] ? 5'hf : _T_2373; // @[CSR.scala 886:74]
  wire [4:0] _T_2377 = raiseExceptionVec[4] ? 5'h4 : _T_2375; // @[CSR.scala 886:74]
  wire [4:0] _T_2379 = raiseExceptionVec[6] ? 5'h6 : _T_2377; // @[CSR.scala 886:74]
  wire [4:0] _T_2381 = raiseExceptionVec[8] ? 5'h8 : _T_2379; // @[CSR.scala 886:74]
  wire [4:0] _T_2383 = raiseExceptionVec[9] ? 5'h9 : _T_2381; // @[CSR.scala 886:74]
  wire [4:0] _T_2385 = raiseExceptionVec[11] ? 5'hb : _T_2383; // @[CSR.scala 886:74]
  wire [4:0] _T_2387 = raiseExceptionVec[0] ? 5'h0 : _T_2385; // @[CSR.scala 886:74]
  wire [4:0] _T_2389 = raiseExceptionVec[2] ? 5'h2 : _T_2387; // @[CSR.scala 886:74]
  wire [4:0] _T_2391 = raiseExceptionVec[1] ? 5'h1 : _T_2389; // @[CSR.scala 886:74]
  wire [4:0] _T_2393 = raiseExceptionVec[12] ? 5'hc : _T_2391; // @[CSR.scala 886:74]
  wire [4:0] exceptionNO = raiseExceptionVec[3] ? 5'h3 : _T_2393; // @[CSR.scala 886:74]
  wire [63:0] _T_2395 = {raiseIntr, 63'h0}; // @[CSR.scala 889:28]
  wire [4:0] _T_2396 = raiseIntr ? {{1'd0}, intrNO} : exceptionNO; // @[CSR.scala 889:46]
  wire [63:0] _GEN_235 = {{59'd0}, _T_2396}; // @[CSR.scala 889:41]
  wire [63:0] causeNO = _T_2395 | _GEN_235; // @[CSR.scala 889:41]
  wire  raiseExceptionIntr = (raiseException | raiseIntr) & io_instrValid; // @[CSR.scala 892:58]
  wire [63:0] delegVecM = raiseIntr ? mideleg : medeleg; // @[CSR.scala 907:22]
  wire [63:0] _T_2428 = delegVecM >> causeNO[4:0]; // @[CSR.scala 910:26]
  wire  delegS = _T_2428[0] & _T_2225; // @[CSR.scala 910:42]
  wire [63:0] delegVecS = raiseIntr ? sideleg : sedeleg; // @[CSR.scala 908:22]
  wire [63:0] _T_2432 = delegVecS >> causeNO[4:0]; // @[CSR.scala 911:26]
  wire  delegU = _T_2432[0] & _T_2221; // @[CSR.scala 911:42]
  wire [63:0] _T_2448 = delegU ? utvec : stvec; // @[CSR.scala 917:32]
  wire [63:0] _T_2449 = delegS ? _T_2448 : mtvec; // @[CSR.scala 917:20]
  wire [38:0] trapTarget = _T_2449[38:0]; // @[CSR.scala 917:62]
  wire [38:0] _GEN_143 = io_in_valid & isSret ? sepc[38:0] : mepc[38:0]; // @[CSR.scala 942:26 CSR.scala 952:15]
  wire [38:0] retTarget = io_in_valid & isUret ? uepc[38:0] : _GEN_143; // @[CSR.scala 955:26 CSR.scala 963:15]
  wire [38:0] _T_2405 = raiseExceptionIntr ? trapTarget : retTarget; // @[CSR.scala 897:61]
  wire  _T_2439 = _T_2111 | io_cfIn_exceptionVec_4 | io_cfIn_exceptionVec_6 | aluULibInstrFault; // @[CSR.scala 912:129]
  wire  _T_2442 = _T_2439 | lsuULibLoadFault | lsuULibStoreFault | aluSLibInstrFault; // @[CSR.scala 913:78]
  wire  _T_2444 = _T_2442 | lsuSLibLoadFault | lsuSLibStoreFault; // @[CSR.scala 914:57]
  wire  _T_2445 = ~_T_2444; // @[CSR.scala 912:17]
  wire  tvalWen = _T_2445 | raiseIntr; // @[CSR.scala 914:79]
  wire [5:0] lo_lo_14 = {mstatusStruct_pie_s,mstatusStruct_pie_u,mstatusStruct_pie_m,mstatusStruct_ie_h,
    mstatusStruct_ie_s,mstatusStruct_ie_u}; // @[CSR.scala 937:27]
  wire [14:0] lo_20 = {mstatusStruct_fs,2'h0,mstatusStruct_hpp,mstatusStruct_spp,1'h1,mstatusStruct_pie_h,lo_lo_14}; // @[CSR.scala 937:27]
  wire [6:0] hi_lo_14 = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,mstatusStruct_mprv,
    mstatusStruct_xs}; // @[CSR.scala 937:27]
  wire [63:0] _T_2500 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,
    mstatusStruct_tsr,hi_lo_14,lo_20}; // @[CSR.scala 937:27]
  wire [1:0] _GEN_136 = io_in_valid & isMret ? mstatusStruct_mpp : priviledgeMode; // @[CSR.scala 929:26 CSR.scala 934:20 CSR.scala 459:31]
  wire [63:0] _GEN_137 = io_in_valid & isMret ? _T_2500 : _GEN_52; // @[CSR.scala 929:26 CSR.scala 937:13]
  wire [1:0] _T_2551 = {1'h0,mstatusStruct_spp}; // @[Cat.scala 30:58]
  wire [5:0] lo_lo_15 = {1'h1,mstatusStruct_pie_u,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_pie_s,
    mstatusStruct_ie_u}; // @[CSR.scala 950:27]
  wire [14:0] lo_21 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,1'h0,mstatusStruct_pie_m,mstatusStruct_pie_h
    ,lo_lo_15}; // @[CSR.scala 950:27]
  wire [63:0] _T_2552 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,
    mstatusStruct_tsr,hi_lo_14,lo_21}; // @[CSR.scala 950:27]
  wire [5:0] lo_lo_16 = {mstatusStruct_pie_s,1'h1,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_ie_s,
    mstatusStruct_pie_u}; // @[CSR.scala 962:27]
  wire [14:0] lo_22 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,mstatusStruct_spp,mstatusStruct_pie_m,
    mstatusStruct_pie_h,lo_lo_16}; // @[CSR.scala 962:27]
  wire [63:0] _T_2603 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,
    mstatusStruct_tsr,hi_lo_14,lo_22}; // @[CSR.scala 962:27]
  wire [63:0] _GEN_148 = tvalWen ? 64'h0 : _GEN_135; // @[CSR.scala 986:20 CSR.scala 986:27]
  wire [63:0] _GEN_149 = tvalWen ? 64'h0 : _GEN_134; // @[CSR.scala 994:20 CSR.scala 994:27]
  wire  _GEN_152 = delegS & delegU ? mstatusStruct_ie_u : mstatusStruct_pie_u; // @[CSR.scala 980:35 CSR.scala 983:24]
  wire  _GEN_153 = delegS & delegU ? 1'h0 : mstatusStruct_ie_u; // @[CSR.scala 980:35 CSR.scala 984:23]
  wire [1:0] _GEN_158 = delegS & delegU ? mstatusStruct_mpp : priviledgeMode; // @[CSR.scala 980:35 CSR.scala 990:22]
  wire  _GEN_159 = delegS & delegU ? mstatusStruct_pie_m : mstatusStruct_ie_m; // @[CSR.scala 980:35 CSR.scala 991:24]
  wire  _GEN_160 = delegS & delegU & mstatusStruct_ie_m; // @[CSR.scala 980:35 CSR.scala 992:23]
  wire [1:0] _GEN_164 = delegS & ~delegU ? priviledgeMode : {{1'd0}, mstatusStruct_spp}; // @[CSR.scala 970:30 CSR.scala 973:22]
  wire  _GEN_165 = delegS & ~delegU ? mstatusStruct_ie_s : mstatusStruct_pie_s; // @[CSR.scala 970:30 CSR.scala 974:24]
  wire  _GEN_166 = delegS & ~delegU ? 1'h0 : mstatusStruct_ie_s; // @[CSR.scala 970:30 CSR.scala 975:23]
  wire  _GEN_171 = delegS & ~delegU ? mstatusStruct_pie_u : _GEN_152; // @[CSR.scala 970:30]
  wire  _GEN_172 = delegS & ~delegU ? mstatusStruct_ie_u : _GEN_153; // @[CSR.scala 970:30]
  wire [1:0] _GEN_176 = delegS & ~delegU ? mstatusStruct_mpp : _GEN_158; // @[CSR.scala 970:30]
  wire  _GEN_177 = delegS & ~delegU ? mstatusStruct_pie_m : _GEN_159; // @[CSR.scala 970:30]
  wire  _GEN_178 = delegS & ~delegU ? mstatusStruct_ie_m : _GEN_160; // @[CSR.scala 970:30]
  wire [5:0] lo_lo_17 = {_GEN_165,_GEN_171,_GEN_178,mstatusStruct_ie_h,_GEN_166,_GEN_172}; // @[CSR.scala 1004:27]
  wire [14:0] lo_23 = {mstatusStruct_fs,_GEN_176,mstatusStruct_hpp,_GEN_164[0],_GEN_177,mstatusStruct_pie_h,lo_lo_17}; // @[CSR.scala 1004:27]
  wire [63:0] _T_2665 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,
    mstatusStruct_tsr,hi_lo_14,lo_23}; // @[CSR.scala 1004:27]
  wire [63:0] _T_2667 = perfCnts_0 + 64'h1; // @[CSR.scala 1113:71]
  wire  _WIRE_52 = 1'h1;
  wire [63:0] _T_2671 = perfCnts_2 + 64'h1; // @[CSR.scala 1113:71]
  wire [63:0] _T_2673 = perfCnts_2 + 64'h2; // @[CSR.scala 1121:86]
  assign io_out_valid = io_in_valid; // @[CSR.scala 1008:16]
  assign io_out_bits = _T_664 | _T_576; // @[Mux.scala 27:72]
  assign io_redirect_target = resetSatp ? _T_2039 : _T_2405; // @[CSR.scala 897:28]
  assign io_redirect_valid = io_in_valid & _T_2070 | raiseExceptionIntr | resetSatp; // @[CSR.scala 895:80]
  assign io_imemMMU_priviledgeMode = priviledgeMode; // @[CSR.scala 769:29]
  assign io_dmemMMU_priviledgeMode = mstatusStruct_mprv ? mstatusStruct_mpp : priviledgeMode; // @[CSR.scala 770:35]
  assign io_dmemMMU_status_sum = mstatus[18]; // @[CSR.scala 335:39]
  assign io_dmemMMU_status_mxr = mstatus[19]; // @[CSR.scala 335:39]
  assign io_wenFix = |raiseExceptionVec; // @[CSR.scala 885:42]
  assign satp_0 = satp;
  assign lsuDeny_0 = lsuDeny;
  assign isuPermitLibLoad_0 = isuPermitLibLoad;
  assign isuPermitLibStore_0 = isuPermitLibStore;
  assign intrVec_0 = intrVec;
  assign lrAddr_0 = lrAddr;
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 287:22]
      mtvec <= 64'h0; // @[CSR.scala 287:22]
    end else if (_T_306 & addr == 12'h305) begin // @[RegMap.scala 50:72]
      mtvec <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 288:27]
      mcounteren <= 64'h0; // @[CSR.scala 288:27]
    end else if (_T_306 & addr == 12'h306) begin // @[RegMap.scala 50:72]
      mcounteren <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 289:23]
      mcause <= 64'h0; // @[CSR.scala 289:23]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 966:29]
      if (delegS & ~delegU) begin // @[CSR.scala 970:30]
        mcause <= _GEN_18;
      end else if (delegS & delegU) begin // @[CSR.scala 980:35]
        mcause <= _GEN_18;
      end else begin
        mcause <= causeNO; // @[CSR.scala 988:14]
      end
    end else begin
      mcause <= _GEN_18;
    end
    if (reset) begin // @[CSR.scala 290:22]
      mtval <= 64'h0; // @[CSR.scala 290:22]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 966:29]
      if (delegS & ~delegU) begin // @[CSR.scala 970:30]
        mtval <= _GEN_134;
      end else if (delegS & delegU) begin // @[CSR.scala 980:35]
        mtval <= _GEN_134;
      end else begin
        mtval <= _GEN_149;
      end
    end else begin
      mtval <= _GEN_134;
    end
    if (reset) begin // @[CSR.scala 291:21]
      mepc <= 64'h0; // @[CSR.scala 291:21]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 966:29]
      if (delegS & ~delegU) begin // @[CSR.scala 970:30]
        mepc <= _GEN_73;
      end else if (delegS & delegU) begin // @[CSR.scala 980:35]
        mepc <= _GEN_73;
      end else begin
        mepc <= _T_2119; // @[CSR.scala 989:12]
      end
    end else begin
      mepc <= _GEN_73;
    end
    if (reset) begin // @[CSR.scala 293:20]
      mie <= 64'h0; // @[CSR.scala 293:20]
    end else if (_T_306 & addr == 12'h304) begin // @[RegMap.scala 50:72]
      mie <= wdata; // @[RegMap.scala 50:76]
    end else if (_T_306 & addr == 12'h104) begin // @[RegMap.scala 50:72]
      mie <= _T_822; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 295:24]
      mipReg <= 64'h0; // @[CSR.scala 295:24]
    end else if (_T_306 & addr == 12'h144) begin // @[RegMap.scala 50:72]
      mipReg <= _T_1458; // @[RegMap.scala 50:76]
    end else if (_T_306 & addr == 12'h344) begin // @[RegMap.scala 50:72]
      mipReg <= _T_1452; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 306:21]
      misa <= 64'h8000000000143105; // @[CSR.scala 306:21]
    end else if (_T_306 & addr == 12'h301) begin // @[RegMap.scala 50:72]
      misa <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 314:24]
      mstatus <= 64'h1800; // @[CSR.scala 314:24]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 966:29]
      mstatus <= _T_2665; // @[CSR.scala 1004:13]
    end else if (io_in_valid & isUret) begin // @[CSR.scala 955:26]
      mstatus <= _T_2603; // @[CSR.scala 962:13]
    end else if (io_in_valid & isSret) begin // @[CSR.scala 942:26]
      mstatus <= _T_2552; // @[CSR.scala 950:13]
    end else begin
      mstatus <= _GEN_137;
    end
    if (reset) begin // @[CSR.scala 342:24]
      medeleg <= 64'h0; // @[CSR.scala 342:24]
    end else if (_T_306 & addr == 12'h302) begin // @[RegMap.scala 50:72]
      medeleg <= _T_768; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 343:24]
      mideleg <= 64'h0; // @[CSR.scala 343:24]
    end else if (_T_306 & addr == 12'h303) begin // @[RegMap.scala 50:72]
      mideleg <= _T_1130; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 344:25]
      mscratch <= 64'h0; // @[CSR.scala 344:25]
    end else if (_T_306 & addr == 12'h340) begin // @[RegMap.scala 50:72]
      mscratch <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 346:24]
      pmpcfg0 <= 64'h0; // @[CSR.scala 346:24]
    end else if (_T_306 & addr == 12'h3a0) begin // @[RegMap.scala 50:72]
      pmpcfg0 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 347:24]
      pmpcfg1 <= 64'h0; // @[CSR.scala 347:24]
    end else if (_T_306 & addr == 12'h3a1) begin // @[RegMap.scala 50:72]
      pmpcfg1 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 348:24]
      pmpcfg2 <= 64'h0; // @[CSR.scala 348:24]
    end else if (_T_306 & addr == 12'h3a2) begin // @[RegMap.scala 50:72]
      pmpcfg2 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 349:24]
      pmpcfg3 <= 64'h0; // @[CSR.scala 349:24]
    end else if (_T_306 & addr == 12'h3a3) begin // @[RegMap.scala 50:72]
      pmpcfg3 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 350:25]
      pmpaddr0 <= 64'h0; // @[CSR.scala 350:25]
    end else if (_T_306 & addr == 12'h3b0) begin // @[RegMap.scala 50:72]
      pmpaddr0 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 351:25]
      pmpaddr1 <= 64'h0; // @[CSR.scala 351:25]
    end else if (_T_306 & addr == 12'h3b1) begin // @[RegMap.scala 50:72]
      pmpaddr1 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 352:25]
      pmpaddr2 <= 64'h0; // @[CSR.scala 352:25]
    end else if (_T_306 & addr == 12'h3b2) begin // @[RegMap.scala 50:72]
      pmpaddr2 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 353:25]
      pmpaddr3 <= 64'h0; // @[CSR.scala 353:25]
    end else if (_T_306 & addr == 12'h3b3) begin // @[RegMap.scala 50:72]
      pmpaddr3 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 356:35]
      dasicsSMainCfg <= 64'h0; // @[CSR.scala 356:35]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      if (dasicsSMainCfg[0]) begin // @[CSR.scala 613:5]
        dasicsSMainCfg <= _T_1463; // @[CSR.scala 617:22]
      end else begin
        dasicsSMainCfg <= _GEN_3;
      end
    end else begin
      dasicsSMainCfg <= _GEN_3;
    end
    if (reset) begin // @[CSR.scala 357:35]
      dasicsSMainBoundHi <= 64'h0; // @[CSR.scala 357:35]
    end else if (_T_306 & addr == 12'hbc1) begin // @[RegMap.scala 50:72]
      dasicsSMainBoundHi <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 358:35]
      dasicsSMainBoundLo <= 64'h0; // @[CSR.scala 358:35]
    end else if (_T_306 & addr == 12'hbc2) begin // @[RegMap.scala 50:72]
      dasicsSMainBoundLo <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 378:22]
      stvec <= 64'h0; // @[CSR.scala 378:22]
    end else if (_T_306 & addr == 12'h105) begin // @[RegMap.scala 50:72]
      stvec <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 383:21]
      satp <= 64'h0; // @[CSR.scala 383:21]
    end else if (_T_306 & addr == 12'h180) begin // @[RegMap.scala 50:72]
      satp <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 384:21]
      sepc <= 64'h0; // @[CSR.scala 384:21]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 966:29]
      if (delegS & ~delegU) begin // @[CSR.scala 970:30]
        sepc <= _T_2119; // @[CSR.scala 972:12]
      end else begin
        sepc <= _GEN_17;
      end
    end else begin
      sepc <= _GEN_17;
    end
    if (reset) begin // @[CSR.scala 385:23]
      scause <= 64'h0; // @[CSR.scala 385:23]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 966:29]
      if (delegS & ~delegU) begin // @[CSR.scala 970:30]
        scause <= causeNO; // @[CSR.scala 971:14]
      end else begin
        scause <= _GEN_80;
      end
    end else begin
      scause <= _GEN_80;
    end
    if (reset) begin // @[CSR.scala 386:22]
      stval <= 64'h0; // @[CSR.scala 386:22]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 966:29]
      if (delegS & ~delegU) begin // @[CSR.scala 970:30]
        if (tvalWen) begin // @[CSR.scala 977:20]
          stval <= 64'h0; // @[CSR.scala 977:27]
        end else begin
          stval <= _GEN_133;
        end
      end else begin
        stval <= _GEN_133;
      end
    end else begin
      stval <= _GEN_133;
    end
    if (reset) begin // @[CSR.scala 387:25]
      sscratch <= 64'h0; // @[CSR.scala 387:25]
    end else if (_T_306 & addr == 12'h140) begin // @[RegMap.scala 50:72]
      sscratch <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 388:27]
      scounteren <= 64'h0; // @[CSR.scala 388:27]
    end else if (_T_306 & addr == 12'h106) begin // @[RegMap.scala 50:72]
      scounteren <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 390:24]
      sedeleg <= 64'h0; // @[CSR.scala 390:24]
    end else if (_T_306 & addr == 12'h102) begin // @[RegMap.scala 50:72]
      sedeleg <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 391:24]
      sideleg <= 64'h0; // @[CSR.scala 391:24]
    end else if (_T_306 & addr == 12'h103) begin // @[RegMap.scala 50:72]
      sideleg <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 394:35]
      dasicsUMainCfg <= 64'h0; // @[CSR.scala 394:35]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsUMainCfg <= _T_1464; // @[CSR.scala 625:20]
    end else if (_T_306 & addr == 12'h5c0) begin // @[RegMap.scala 50:72]
      dasicsUMainCfg <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 395:35]
      dasicsUMainBoundHi <= 64'h0; // @[CSR.scala 395:35]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      if (dasicsSMainCfg[0]) begin // @[CSR.scala 613:5]
        dasicsUMainBoundHi <= 64'h0; // @[CSR.scala 614:26]
      end else begin
        dasicsUMainBoundHi <= _GEN_78;
      end
    end else begin
      dasicsUMainBoundHi <= _GEN_78;
    end
    if (reset) begin // @[CSR.scala 396:35]
      dasicsUMainBoundLo <= 64'h0; // @[CSR.scala 396:35]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      if (dasicsSMainCfg[0]) begin // @[CSR.scala 613:5]
        dasicsUMainBoundLo <= 64'h0; // @[CSR.scala 615:26]
      end else begin
        dasicsUMainBoundLo <= _GEN_50;
      end
    end else begin
      dasicsUMainBoundLo <= _GEN_50;
    end
    if (reset) begin // @[CSR.scala 413:21]
      uepc <= 64'h0; // @[CSR.scala 413:21]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 966:29]
      if (delegS & ~delegU) begin // @[CSR.scala 970:30]
        uepc <= _GEN_24;
      end else if (delegS & delegU) begin // @[CSR.scala 980:35]
        uepc <= _T_2119; // @[CSR.scala 982:12]
      end else begin
        uepc <= _GEN_24;
      end
    end else begin
      uepc <= _GEN_24;
    end
    if (reset) begin // @[CSR.scala 414:23]
      ucause <= 64'h0; // @[CSR.scala 414:23]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 966:29]
      if (delegS & ~delegU) begin // @[CSR.scala 970:30]
        ucause <= _GEN_48;
      end else if (delegS & delegU) begin // @[CSR.scala 980:35]
        ucause <= causeNO; // @[CSR.scala 981:14]
      end else begin
        ucause <= _GEN_48;
      end
    end else begin
      ucause <= _GEN_48;
    end
    if (reset) begin // @[CSR.scala 415:25]
      uscratch <= 64'h0; // @[CSR.scala 415:25]
    end else if (_T_306 & addr == 12'h40) begin // @[RegMap.scala 50:72]
      uscratch <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 416:22]
      utvec <= 64'h0; // @[CSR.scala 416:22]
    end else if (_T_306 & addr == 12'h5) begin // @[RegMap.scala 50:72]
      utvec <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 417:22]
      utval <= 64'h0; // @[CSR.scala 417:22]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 966:29]
      if (delegS & ~delegU) begin // @[CSR.scala 970:30]
        utval <= _GEN_135;
      end else if (delegS & delegU) begin // @[CSR.scala 980:35]
        utval <= _GEN_148;
      end else begin
        utval <= _GEN_135;
      end
    end else begin
      utval <= _GEN_135;
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_0 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_0 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h883) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_0 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_1 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_1 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h885) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_1 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_2 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_2 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h887) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_2 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_3 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_3 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h889) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_3 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_4 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_4 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h88b) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_4 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_5 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_5 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h88d) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_5 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_6 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_6 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h88f) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_6 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_7 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_7 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h891) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_7 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_8 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_8 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h893) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_8 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_9 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_9 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h895) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_9 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_10 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_10 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h897) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_10 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_11 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_11 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h899) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_11 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_12 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_12 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h89b) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_12 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_13 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_13 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h89d) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_13 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_14 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_14 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h89f) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_14 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 420:64]
      dasicsLibBoundHiList_15 <= 64'h0; // @[CSR.scala 420:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundHiList_15 <= 64'h0; // @[CSR.scala 620:45]
    end else if (_T_306 & addr == 12'h8a1) begin // @[RegMap.scala 50:72]
      dasicsLibBoundHiList_15 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_0 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_0 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h884) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_0 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_1 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_1 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h886) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_1 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_2 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_2 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h888) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_2 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_3 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_3 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h88a) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_3 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_4 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_4 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h88c) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_4 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_5 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_5 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h88e) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_5 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_6 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_6 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h890) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_6 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_7 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_7 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h892) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_7 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_8 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_8 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h894) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_8 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_9 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_9 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h896) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_9 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_10 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_10 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h898) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_10 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_11 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_11 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h89a) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_11 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_12 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_12 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h89c) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_12 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_13 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_13 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h89e) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_13 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_14 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_14 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h8a0) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_14 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 421:64]
      dasicsLibBoundLoList_15 <= 64'h0; // @[CSR.scala 421:64]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibBoundLoList_15 <= 64'h0; // @[CSR.scala 621:45]
    end else if (_T_306 & addr == 12'h8a2) begin // @[RegMap.scala 50:72]
      dasicsLibBoundLoList_15 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 425:31]
      dasicsLibCfg0 <= 64'h0; // @[CSR.scala 425:31]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibCfg0 <= 64'h0; // @[CSR.scala 622:19]
    end else if (_T_306 & addr == 12'h881) begin // @[RegMap.scala 50:72]
      dasicsLibCfg0 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 426:31]
      dasicsLibCfg1 <= 64'h0; // @[CSR.scala 426:31]
    end else if (_T_1461) begin // @[CSR.scala 611:3]
      dasicsLibCfg1 <= 64'h0; // @[CSR.scala 623:19]
    end else if (_T_306 & addr == 12'h882) begin // @[RegMap.scala 50:72]
      dasicsLibCfg1 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 427:31]
      dasicsReturnPC <= 64'h0; // @[CSR.scala 427:31]
    end else if (_T_2037) begin // @[CSR.scala 708:3]
      dasicsReturnPC <= {{25'd0}, _T_2039}; // @[CSR.scala 709:20]
    end else if (_T_306 & addr == 12'h8a4) begin // @[RegMap.scala 50:72]
      dasicsReturnPC <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 428:39]
      dasicsFreeZoneReturnPC <= 64'h0; // @[CSR.scala 428:39]
    end else if (_T_2044) begin // @[CSR.scala 713:3]
      dasicsFreeZoneReturnPC <= {{25'd0}, _T_2039}; // @[CSR.scala 714:28]
    end else if (_T_306 & addr == 12'h8a5) begin // @[RegMap.scala 50:72]
      dasicsFreeZoneReturnPC <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 429:39]
      dasicsMaincallEntry <= 64'h0; // @[CSR.scala 429:39]
    end else if (_T_306 & addr == 12'h8a3) begin // @[RegMap.scala 50:72]
      dasicsMaincallEntry <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 445:19]
      lr <= 1'h0; // @[CSR.scala 445:19]
    end else if (io_in_valid & isSret) begin // @[CSR.scala 942:26]
      lr <= 1'h0; // @[CSR.scala 951:8]
    end else if (io_in_valid & isMret) begin // @[CSR.scala 929:26]
      lr <= 1'h0; // @[CSR.scala 938:8]
    end else if (set_lr) begin // @[CSR.scala 453:14]
      lr <= set_lr_val; // @[CSR.scala 454:8]
    end
    if (reset) begin // @[CSR.scala 446:23]
      lrAddr <= 64'h0; // @[CSR.scala 446:23]
    end else if (set_lr) begin // @[CSR.scala 453:14]
      lrAddr <= set_lr_addr; // @[CSR.scala 455:12]
    end
    if (reset) begin // @[CSR.scala 459:31]
      priviledgeMode <= 2'h3; // @[CSR.scala 459:31]
    end else if (raiseExceptionIntr) begin // @[CSR.scala 966:29]
      if (delegS & ~delegU) begin // @[CSR.scala 970:30]
        priviledgeMode <= 2'h1; // @[CSR.scala 976:22]
      end else if (delegS & delegU) begin // @[CSR.scala 980:35]
        priviledgeMode <= 2'h0; // @[CSR.scala 985:22]
      end else begin
        priviledgeMode <= 2'h3; // @[CSR.scala 993:22]
      end
    end else if (io_in_valid & isUret) begin // @[CSR.scala 955:26]
      priviledgeMode <= 2'h0; // @[CSR.scala 960:20]
    end else if (io_in_valid & isSret) begin // @[CSR.scala 942:26]
      priviledgeMode <= _T_2551; // @[CSR.scala 947:20]
    end else begin
      priviledgeMode <= _GEN_136;
    end
    if (reset) begin // @[CSR.scala 464:47]
      perfCnts_0 <= 64'h0; // @[CSR.scala 464:47]
    end else begin
      perfCnts_0 <= _T_2667;
    end
    if (reset) begin // @[CSR.scala 464:47]
      perfCnts_1 <= 64'h0; // @[CSR.scala 464:47]
    end else if (_T_306 & addr == 12'hb01) begin // @[RegMap.scala 50:72]
      perfCnts_1 <= wdata; // @[RegMap.scala 50:76]
    end
    if (reset) begin // @[CSR.scala 464:47]
      perfCnts_2 <= 64'h0; // @[CSR.scala 464:47]
    end else if (perfCntCondMultiCommit) begin // @[CSR.scala 1121:35]
      perfCnts_2 <= _T_2673; // @[CSR.scala 1121:60]
    end else if (perfCntCondMinstret) begin // @[CSR.scala 1113:62]
      perfCnts_2 <= _T_2671; // @[CSR.scala 1113:66]
    end else if (_T_306 & addr == 12'hb02) begin // @[RegMap.scala 50:72]
      perfCnts_2 <= wdata; // @[RegMap.scala 50:76]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtvec = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mcounteren = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mcause = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mtval = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mepc = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mie = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mipReg = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  misa = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mstatus = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  medeleg = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  mideleg = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mscratch = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  pmpcfg0 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  pmpcfg1 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  pmpcfg2 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  pmpcfg3 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  pmpaddr0 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  pmpaddr1 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  pmpaddr2 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  pmpaddr3 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  dasicsSMainCfg = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  dasicsSMainBoundHi = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  dasicsSMainBoundLo = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  stvec = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  satp = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  sepc = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  scause = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  stval = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  sscratch = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  scounteren = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  sedeleg = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  sideleg = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  dasicsUMainCfg = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  dasicsUMainBoundHi = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  dasicsUMainBoundLo = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  uepc = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  ucause = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  uscratch = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  utvec = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  utval = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  dasicsLibBoundHiList_0 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  dasicsLibBoundHiList_1 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  dasicsLibBoundHiList_2 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  dasicsLibBoundHiList_3 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  dasicsLibBoundHiList_4 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  dasicsLibBoundHiList_5 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  dasicsLibBoundHiList_6 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  dasicsLibBoundHiList_7 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  dasicsLibBoundHiList_8 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  dasicsLibBoundHiList_9 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  dasicsLibBoundHiList_10 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  dasicsLibBoundHiList_11 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  dasicsLibBoundHiList_12 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  dasicsLibBoundHiList_13 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  dasicsLibBoundHiList_14 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  dasicsLibBoundHiList_15 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  dasicsLibBoundLoList_0 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  dasicsLibBoundLoList_1 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  dasicsLibBoundLoList_2 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  dasicsLibBoundLoList_3 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  dasicsLibBoundLoList_4 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  dasicsLibBoundLoList_5 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  dasicsLibBoundLoList_6 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  dasicsLibBoundLoList_7 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  dasicsLibBoundLoList_8 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  dasicsLibBoundLoList_9 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  dasicsLibBoundLoList_10 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  dasicsLibBoundLoList_11 = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  dasicsLibBoundLoList_12 = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  dasicsLibBoundLoList_13 = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  dasicsLibBoundLoList_14 = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  dasicsLibBoundLoList_15 = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  dasicsLibCfg0 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  dasicsLibCfg1 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  dasicsReturnPC = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  dasicsFreeZoneReturnPC = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  dasicsMaincallEntry = _RAND_76[63:0];
  _RAND_77 = {1{`RANDOM}};
  lr = _RAND_77[0:0];
  _RAND_78 = {2{`RANDOM}};
  lrAddr = _RAND_78[63:0];
  _RAND_79 = {1{`RANDOM}};
  priviledgeMode = _RAND_79[1:0];
  _RAND_80 = {2{`RANDOM}};
  perfCnts_0 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  perfCnts_1 = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  perfCnts_2 = _RAND_82[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_MOU(
  input         io_in_valid,
  input  [6:0]  io_in_bits_func,
  input  [38:0] io_cfIn_pc,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  output        flushICache_0,
  output        flushTLB_0
);
  wire  flushICache = io_in_valid & io_in_bits_func == 7'h1; // @[MOU.scala 52:27]
  wire  flushTLB = io_in_valid & io_in_bits_func == 7'h2; // @[MOU.scala 56:24]
  assign io_redirect_target = io_cfIn_pc + 39'h4; // @[MOU.scala 49:36]
  assign io_redirect_valid = io_in_valid; // @[MOU.scala 50:21]
  assign flushICache_0 = flushICache;
  assign flushTLB_0 = flushTLB;
endmodule
module ysyx_210000_EXU(
  input         clock,
  input         reset,
  output        io__in_ready,
  input         io__in_valid,
  input  [63:0] io__in_bits_cf_instr,
  input  [38:0] io__in_bits_cf_pc,
  input  [38:0] io__in_bits_cf_pnpc,
  input         io__in_bits_cf_exceptionVec_1,
  input         io__in_bits_cf_exceptionVec_2,
  input         io__in_bits_cf_exceptionVec_12,
  input         io__in_bits_cf_intrVec_0,
  input         io__in_bits_cf_intrVec_1,
  input         io__in_bits_cf_intrVec_2,
  input         io__in_bits_cf_intrVec_3,
  input         io__in_bits_cf_intrVec_4,
  input         io__in_bits_cf_intrVec_5,
  input         io__in_bits_cf_intrVec_6,
  input         io__in_bits_cf_intrVec_7,
  input         io__in_bits_cf_intrVec_8,
  input         io__in_bits_cf_intrVec_9,
  input         io__in_bits_cf_intrVec_10,
  input         io__in_bits_cf_intrVec_11,
  input  [3:0]  io__in_bits_cf_brIdx,
  input         io__in_bits_cf_crossPageIPFFix,
  input  [2:0]  io__in_bits_ctrl_fuType,
  input  [6:0]  io__in_bits_ctrl_fuOpType,
  input         io__in_bits_ctrl_rfWen,
  input  [4:0]  io__in_bits_ctrl_rfDest,
  input         io__in_bits_ctrl_permitLibLoad,
  input         io__in_bits_ctrl_permitLibStore,
  input         io__in_bits_ctrl_lsuIsLoad,
  input  [63:0] io__in_bits_data_src1,
  input  [63:0] io__in_bits_data_src2,
  input  [63:0] io__in_bits_data_imm,
  input  [63:0] io__in_bits_data_addr,
  input         io__out_ready,
  output        io__out_valid,
  output [38:0] io__out_bits_decode_cf_pc,
  output [38:0] io__out_bits_decode_cf_redirect_target,
  output        io__out_bits_decode_cf_redirect_valid,
  output [2:0]  io__out_bits_decode_ctrl_fuType,
  output        io__out_bits_decode_ctrl_rfWen,
  output [4:0]  io__out_bits_decode_ctrl_rfDest,
  output [63:0] io__out_bits_commits_0,
  output [63:0] io__out_bits_commits_1,
  output [63:0] io__out_bits_commits_2,
  output [63:0] io__out_bits_commits_3,
  input         io__flush,
  input         io__dmem_req_ready,
  output        io__dmem_req_valid,
  output [38:0] io__dmem_req_bits_addr,
  output [2:0]  io__dmem_req_bits_size,
  output [3:0]  io__dmem_req_bits_cmd,
  output [7:0]  io__dmem_req_bits_wmask,
  output [63:0] io__dmem_req_bits_wdata,
  input         io__dmem_resp_valid,
  input  [63:0] io__dmem_resp_bits_rdata,
  output        io__forward_valid,
  output        io__forward_wb_rfWen,
  output [4:0]  io__forward_wb_rfDest,
  output [63:0] io__forward_wb_rfData,
  output [2:0]  io__forward_fuType,
  output [1:0]  io__memMMU_imem_priviledgeMode,
  output [1:0]  io__memMMU_dmem_priviledgeMode,
  output        io__memMMU_dmem_status_sum,
  output        io__memMMU_dmem_status_mxr,
  input         io__memMMU_dmem_loadPF,
  input         io__memMMU_dmem_storePF,
  input  [38:0] io__memMMU_dmem_addr,
  input         _T_28_0,
  output        flushICache,
  output [63:0] satp,
  output        REG_6_valid,
  output [38:0] REG_6_pc,
  output        REG_6_isMissPredict,
  output [38:0] REG_6_actualTarget,
  output        REG_6_actualTaken,
  output [6:0]  REG_6_fuOpType,
  output [1:0]  REG_6_btbType,
  output        REG_6_isRVC,
  input         io_in_valid,
  input         io_extra_mtip,
  output        amoReq,
  input         io_extra_meip_0,
  input         vmEnable,
  input  [63:0] isuAddr,
  output        isuPermitLibLoad,
  output        isuPermitLibStore,
  output [11:0] intrVec,
  input         _T_27_0,
  input         io_extra_msip,
  output        flushTLB,
  input         falseWire
);
  wire  alu_clock; // @[EXU.scala 45:19]
  wire  alu_reset; // @[EXU.scala 45:19]
  wire  alu_io__in_valid; // @[EXU.scala 45:19]
  wire [63:0] alu_io__in_bits_src1; // @[EXU.scala 45:19]
  wire [63:0] alu_io__in_bits_src2; // @[EXU.scala 45:19]
  wire [6:0] alu_io__in_bits_func; // @[EXU.scala 45:19]
  wire  alu_io__out_ready; // @[EXU.scala 45:19]
  wire  alu_io__out_valid; // @[EXU.scala 45:19]
  wire [63:0] alu_io__out_bits; // @[EXU.scala 45:19]
  wire [63:0] alu_io__cfIn_instr; // @[EXU.scala 45:19]
  wire [38:0] alu_io__cfIn_pc; // @[EXU.scala 45:19]
  wire [38:0] alu_io__cfIn_pnpc; // @[EXU.scala 45:19]
  wire [3:0] alu_io__cfIn_brIdx; // @[EXU.scala 45:19]
  wire [38:0] alu_io__redirect_target; // @[EXU.scala 45:19]
  wire  alu_io__redirect_valid; // @[EXU.scala 45:19]
  wire [63:0] alu_io__offset; // @[EXU.scala 45:19]
  wire  alu__T_113_0; // @[EXU.scala 45:19]
  wire  alu_REG_6_0_valid; // @[EXU.scala 45:19]
  wire [38:0] alu_REG_6_0_pc; // @[EXU.scala 45:19]
  wire  alu_REG_6_0_isMissPredict; // @[EXU.scala 45:19]
  wire [38:0] alu_REG_6_0_actualTarget; // @[EXU.scala 45:19]
  wire  alu_REG_6_0_actualTaken; // @[EXU.scala 45:19]
  wire [6:0] alu_REG_6_0_fuOpType; // @[EXU.scala 45:19]
  wire [1:0] alu_REG_6_0_btbType; // @[EXU.scala 45:19]
  wire  alu_REG_6_0_isRVC; // @[EXU.scala 45:19]
  wire  alu_io_redirect_valid; // @[EXU.scala 45:19]
  wire [38:0] alu_io_redirect_target; // @[EXU.scala 45:19]
  wire  lsu_clock; // @[EXU.scala 53:19]
  wire  lsu_reset; // @[EXU.scala 53:19]
  wire  lsu_io__in_valid; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__in_bits_src1; // @[EXU.scala 53:19]
  wire [6:0] lsu_io__in_bits_func; // @[EXU.scala 53:19]
  wire  lsu_io__out_ready; // @[EXU.scala 53:19]
  wire  lsu_io__out_valid; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__out_bits; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__srcSum; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__wdata; // @[EXU.scala 53:19]
  wire [31:0] lsu_io__instr; // @[EXU.scala 53:19]
  wire  lsu_io__dmem_req_ready; // @[EXU.scala 53:19]
  wire  lsu_io__dmem_req_valid; // @[EXU.scala 53:19]
  wire [38:0] lsu_io__dmem_req_bits_addr; // @[EXU.scala 53:19]
  wire [2:0] lsu_io__dmem_req_bits_size; // @[EXU.scala 53:19]
  wire [3:0] lsu_io__dmem_req_bits_cmd; // @[EXU.scala 53:19]
  wire [7:0] lsu_io__dmem_req_bits_wmask; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__dmem_req_bits_wdata; // @[EXU.scala 53:19]
  wire  lsu_io__dmem_resp_valid; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__dmem_resp_bits_rdata; // @[EXU.scala 53:19]
  wire  lsu_io__dtlbPF; // @[EXU.scala 53:19]
  wire  lsu_io__loadAddrMisaligned; // @[EXU.scala 53:19]
  wire  lsu_io__storeAddrMisaligned; // @[EXU.scala 53:19]
  wire  lsu_setLr_0; // @[EXU.scala 53:19]
  wire  lsu_DTLBPF; // @[EXU.scala 53:19]
  wire  lsu_amoReq_0; // @[EXU.scala 53:19]
  wire  lsu_cannot_access_memory; // @[EXU.scala 53:19]
  wire  lsu_DTLBENABLE; // @[EXU.scala 53:19]
  wire [63:0] lsu_io_in_bits_src1; // @[EXU.scala 53:19]
  wire  lsu_DTLBFINISH; // @[EXU.scala 53:19]
  wire  lsu__T_20_0; // @[EXU.scala 53:19]
  wire [63:0] lsu_setLrAddr_0; // @[EXU.scala 53:19]
  wire [63:0] lsu__T_28_0; // @[EXU.scala 53:19]
  wire  lsu_setLrVal_0; // @[EXU.scala 53:19]
  wire [63:0] lsu_lr_addr; // @[EXU.scala 53:19]
  wire  mdu_clock; // @[EXU.scala 63:19]
  wire  mdu_reset; // @[EXU.scala 63:19]
  wire  mdu_io_in_ready; // @[EXU.scala 63:19]
  wire  mdu_io_in_valid; // @[EXU.scala 63:19]
  wire [63:0] mdu_io_in_bits_src1; // @[EXU.scala 63:19]
  wire [63:0] mdu_io_in_bits_src2; // @[EXU.scala 63:19]
  wire [6:0] mdu_io_in_bits_func; // @[EXU.scala 63:19]
  wire  mdu_io_out_ready; // @[EXU.scala 63:19]
  wire  mdu_io_out_valid; // @[EXU.scala 63:19]
  wire [63:0] mdu_io_out_bits; // @[EXU.scala 63:19]
  wire  csr_clock; // @[EXU.scala 68:19]
  wire  csr_reset; // @[EXU.scala 68:19]
  wire  csr_io_in_valid; // @[EXU.scala 68:19]
  wire [63:0] csr_io_in_bits_src1; // @[EXU.scala 68:19]
  wire [63:0] csr_io_in_bits_src2; // @[EXU.scala 68:19]
  wire [6:0] csr_io_in_bits_func; // @[EXU.scala 68:19]
  wire  csr_io_out_ready; // @[EXU.scala 68:19]
  wire  csr_io_out_valid; // @[EXU.scala 68:19]
  wire [63:0] csr_io_out_bits; // @[EXU.scala 68:19]
  wire [63:0] csr_io_cfIn_instr; // @[EXU.scala 68:19]
  wire [38:0] csr_io_cfIn_pc; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_exceptionVec_1; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_exceptionVec_2; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_exceptionVec_4; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_exceptionVec_6; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_exceptionVec_12; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_0; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_1; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_2; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_3; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_4; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_5; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_6; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_7; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_8; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_9; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_10; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_intrVec_11; // @[EXU.scala 68:19]
  wire  csr_io_cfIn_crossPageIPFFix; // @[EXU.scala 68:19]
  wire [38:0] csr_io_redirect_target; // @[EXU.scala 68:19]
  wire  csr_io_redirect_valid; // @[EXU.scala 68:19]
  wire  csr_io_instrValid; // @[EXU.scala 68:19]
  wire  csr_io_lsuIsLoad; // @[EXU.scala 68:19]
  wire  csr_io_lsuPermitLibLoad; // @[EXU.scala 68:19]
  wire  csr_io_lsuPermitLibStore; // @[EXU.scala 68:19]
  wire [1:0] csr_io_imemMMU_priviledgeMode; // @[EXU.scala 68:19]
  wire [1:0] csr_io_dmemMMU_priviledgeMode; // @[EXU.scala 68:19]
  wire  csr_io_dmemMMU_status_sum; // @[EXU.scala 68:19]
  wire  csr_io_dmemMMU_status_mxr; // @[EXU.scala 68:19]
  wire  csr_io_dmemMMU_loadPF; // @[EXU.scala 68:19]
  wire  csr_io_dmemMMU_storePF; // @[EXU.scala 68:19]
  wire [38:0] csr_io_dmemMMU_addr; // @[EXU.scala 68:19]
  wire  csr_io_wenFix; // @[EXU.scala 68:19]
  wire  csr_set_lr; // @[EXU.scala 68:19]
  wire  csr_is_pulpret; // @[EXU.scala 68:19]
  wire [63:0] csr_satp_0; // @[EXU.scala 68:19]
  wire  csr_perfCntCondMinstret; // @[EXU.scala 68:19]
  wire  csr_mtip_0; // @[EXU.scala 68:19]
  wire  csr_lsuDeny_0; // @[EXU.scala 68:19]
  wire  csr_meip_0; // @[EXU.scala 68:19]
  wire  csr_redirect_valid; // @[EXU.scala 68:19]
  wire [63:0] csr_isu_addr; // @[EXU.scala 68:19]
  wire  csr_isuPermitLibLoad_0; // @[EXU.scala 68:19]
  wire  csr_isuPermitLibStore_0; // @[EXU.scala 68:19]
  wire [38:0] csr_redirect_target; // @[EXU.scala 68:19]
  wire [63:0] csr_LSUEXECADDR; // @[EXU.scala 68:19]
  wire [11:0] csr_intrVec_0; // @[EXU.scala 68:19]
  wire  csr_msip_0; // @[EXU.scala 68:19]
  wire  csr_lsu_is_valid; // @[EXU.scala 68:19]
  wire [63:0] csr_set_lr_addr; // @[EXU.scala 68:19]
  wire [63:0] csr_lsu_addr; // @[EXU.scala 68:19]
  wire  csr_perfCntCondMultiCommit; // @[EXU.scala 68:19]
  wire  csr_set_lr_val; // @[EXU.scala 68:19]
  wire [63:0] csr_lrAddr_0; // @[EXU.scala 68:19]
  wire  mou_io_in_valid; // @[EXU.scala 85:19]
  wire [6:0] mou_io_in_bits_func; // @[EXU.scala 85:19]
  wire [38:0] mou_io_cfIn_pc; // @[EXU.scala 85:19]
  wire [38:0] mou_io_redirect_target; // @[EXU.scala 85:19]
  wire  mou_io_redirect_valid; // @[EXU.scala 85:19]
  wire  mou_flushICache_0; // @[EXU.scala 85:19]
  wire  mou_flushTLB_0; // @[EXU.scala 85:19]
  wire  _T_2 = ~io__flush; // @[EXU.scala 43:84]
  wire  fuValids_1 = io__in_bits_ctrl_fuType == 3'h1 & io__in_valid & ~io__flush; // @[EXU.scala 43:81]
  wire  fuValids_3 = io__in_bits_ctrl_fuType == 3'h3 & io__in_valid & ~io__flush; // @[EXU.scala 43:81]
  wire  lsuTlbPF = lsu_io__dtlbPF;
  wire [38:0] _T_42_target = csr_io_redirect_valid ? csr_io_redirect_target : alu_io__redirect_target; // @[EXU.scala 101:10]
  wire  _T_42_valid = csr_io_redirect_valid ? csr_io_redirect_valid : alu_io__redirect_valid; // @[EXU.scala 101:10]
  wire  _T_55 = 3'h1 == io__in_bits_ctrl_fuType ? lsu_io__out_valid : 1'h1; // @[Mux.scala 80:57]
  wire  _T_57 = 3'h2 == io__in_bits_ctrl_fuType ? mdu_io_out_valid : _T_55; // @[Mux.scala 80:57]
  wire  _T_62 = alu_io__out_ready & alu_io__out_valid; // @[Decoupled.scala 40:37]
  wire  isBru = io__in_bits_ctrl_fuOpType[4]; // @[ALU.scala 64:31]
  wire  _T_66 = _T_62 & ~isBru; // @[EXU.scala 127:43]
  wire  _T_68 = _T_62 & isBru; // @[EXU.scala 128:43]
  wire  _T_69 = lsu_io__out_ready & lsu_io__out_valid; // @[Decoupled.scala 40:37]
  wire  _T_70 = mdu_io_out_ready & mdu_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_71 = csr_io_out_ready & csr_io_out_valid; // @[Decoupled.scala 40:37]
  ysyx_210000_ALU alu ( // @[EXU.scala 45:19]
    .clock(alu_clock),
    .reset(alu_reset),
    .io__in_valid(alu_io__in_valid),
    .io__in_bits_src1(alu_io__in_bits_src1),
    .io__in_bits_src2(alu_io__in_bits_src2),
    .io__in_bits_func(alu_io__in_bits_func),
    .io__out_ready(alu_io__out_ready),
    .io__out_valid(alu_io__out_valid),
    .io__out_bits(alu_io__out_bits),
    .io__cfIn_instr(alu_io__cfIn_instr),
    .io__cfIn_pc(alu_io__cfIn_pc),
    .io__cfIn_pnpc(alu_io__cfIn_pnpc),
    .io__cfIn_brIdx(alu_io__cfIn_brIdx),
    .io__redirect_target(alu_io__redirect_target),
    .io__redirect_valid(alu_io__redirect_valid),
    .io__offset(alu_io__offset),
    ._T_113_0(alu__T_113_0),
    .REG_6_0_valid(alu_REG_6_0_valid),
    .REG_6_0_pc(alu_REG_6_0_pc),
    .REG_6_0_isMissPredict(alu_REG_6_0_isMissPredict),
    .REG_6_0_actualTarget(alu_REG_6_0_actualTarget),
    .REG_6_0_actualTaken(alu_REG_6_0_actualTaken),
    .REG_6_0_fuOpType(alu_REG_6_0_fuOpType),
    .REG_6_0_btbType(alu_REG_6_0_btbType),
    .REG_6_0_isRVC(alu_REG_6_0_isRVC),
    .io_redirect_valid(alu_io_redirect_valid),
    .io_redirect_target(alu_io_redirect_target)
  );
  ysyx_210000_UnpipelinedLSU lsu ( // @[EXU.scala 53:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io__in_valid(lsu_io__in_valid),
    .io__in_bits_src1(lsu_io__in_bits_src1),
    .io__in_bits_func(lsu_io__in_bits_func),
    .io__out_ready(lsu_io__out_ready),
    .io__out_valid(lsu_io__out_valid),
    .io__out_bits(lsu_io__out_bits),
    .io__srcSum(lsu_io__srcSum),
    .io__wdata(lsu_io__wdata),
    .io__instr(lsu_io__instr),
    .io__dmem_req_ready(lsu_io__dmem_req_ready),
    .io__dmem_req_valid(lsu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(lsu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsu_io__dmem_resp_bits_rdata),
    .io__dtlbPF(lsu_io__dtlbPF),
    .io__loadAddrMisaligned(lsu_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsu_io__storeAddrMisaligned),
    .setLr_0(lsu_setLr_0),
    .DTLBPF(lsu_DTLBPF),
    .amoReq_0(lsu_amoReq_0),
    .cannot_access_memory(lsu_cannot_access_memory),
    .DTLBENABLE(lsu_DTLBENABLE),
    .io_in_bits_src1(lsu_io_in_bits_src1),
    .DTLBFINISH(lsu_DTLBFINISH),
    ._T_20_0(lsu__T_20_0),
    .setLrAddr_0(lsu_setLrAddr_0),
    ._T_28_0(lsu__T_28_0),
    .setLrVal_0(lsu_setLrVal_0),
    .lr_addr(lsu_lr_addr)
  );
  ysyx_210000_MDU mdu ( // @[EXU.scala 63:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_in_ready(mdu_io_in_ready),
    .io_in_valid(mdu_io_in_valid),
    .io_in_bits_src1(mdu_io_in_bits_src1),
    .io_in_bits_src2(mdu_io_in_bits_src2),
    .io_in_bits_func(mdu_io_in_bits_func),
    .io_out_ready(mdu_io_out_ready),
    .io_out_valid(mdu_io_out_valid),
    .io_out_bits(mdu_io_out_bits)
  );
  ysyx_210000_CSR csr ( // @[EXU.scala 68:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_in_valid(csr_io_in_valid),
    .io_in_bits_src1(csr_io_in_bits_src1),
    .io_in_bits_src2(csr_io_in_bits_src2),
    .io_in_bits_func(csr_io_in_bits_func),
    .io_out_ready(csr_io_out_ready),
    .io_out_valid(csr_io_out_valid),
    .io_out_bits(csr_io_out_bits),
    .io_cfIn_instr(csr_io_cfIn_instr),
    .io_cfIn_pc(csr_io_cfIn_pc),
    .io_cfIn_exceptionVec_1(csr_io_cfIn_exceptionVec_1),
    .io_cfIn_exceptionVec_2(csr_io_cfIn_exceptionVec_2),
    .io_cfIn_exceptionVec_4(csr_io_cfIn_exceptionVec_4),
    .io_cfIn_exceptionVec_6(csr_io_cfIn_exceptionVec_6),
    .io_cfIn_exceptionVec_12(csr_io_cfIn_exceptionVec_12),
    .io_cfIn_intrVec_0(csr_io_cfIn_intrVec_0),
    .io_cfIn_intrVec_1(csr_io_cfIn_intrVec_1),
    .io_cfIn_intrVec_2(csr_io_cfIn_intrVec_2),
    .io_cfIn_intrVec_3(csr_io_cfIn_intrVec_3),
    .io_cfIn_intrVec_4(csr_io_cfIn_intrVec_4),
    .io_cfIn_intrVec_5(csr_io_cfIn_intrVec_5),
    .io_cfIn_intrVec_6(csr_io_cfIn_intrVec_6),
    .io_cfIn_intrVec_7(csr_io_cfIn_intrVec_7),
    .io_cfIn_intrVec_8(csr_io_cfIn_intrVec_8),
    .io_cfIn_intrVec_9(csr_io_cfIn_intrVec_9),
    .io_cfIn_intrVec_10(csr_io_cfIn_intrVec_10),
    .io_cfIn_intrVec_11(csr_io_cfIn_intrVec_11),
    .io_cfIn_crossPageIPFFix(csr_io_cfIn_crossPageIPFFix),
    .io_redirect_target(csr_io_redirect_target),
    .io_redirect_valid(csr_io_redirect_valid),
    .io_instrValid(csr_io_instrValid),
    .io_lsuIsLoad(csr_io_lsuIsLoad),
    .io_lsuPermitLibLoad(csr_io_lsuPermitLibLoad),
    .io_lsuPermitLibStore(csr_io_lsuPermitLibStore),
    .io_imemMMU_priviledgeMode(csr_io_imemMMU_priviledgeMode),
    .io_dmemMMU_priviledgeMode(csr_io_dmemMMU_priviledgeMode),
    .io_dmemMMU_status_sum(csr_io_dmemMMU_status_sum),
    .io_dmemMMU_status_mxr(csr_io_dmemMMU_status_mxr),
    .io_dmemMMU_loadPF(csr_io_dmemMMU_loadPF),
    .io_dmemMMU_storePF(csr_io_dmemMMU_storePF),
    .io_dmemMMU_addr(csr_io_dmemMMU_addr),
    .io_wenFix(csr_io_wenFix),
    .set_lr(csr_set_lr),
    .is_pulpret(csr_is_pulpret),
    .satp_0(csr_satp_0),
    .perfCntCondMinstret(csr_perfCntCondMinstret),
    .mtip_0(csr_mtip_0),
    .lsuDeny_0(csr_lsuDeny_0),
    .meip_0(csr_meip_0),
    .redirect_valid(csr_redirect_valid),
    .isu_addr(csr_isu_addr),
    .isuPermitLibLoad_0(csr_isuPermitLibLoad_0),
    .isuPermitLibStore_0(csr_isuPermitLibStore_0),
    .redirect_target(csr_redirect_target),
    .LSUEXECADDR(csr_LSUEXECADDR),
    .intrVec_0(csr_intrVec_0),
    .msip_0(csr_msip_0),
    .lsu_is_valid(csr_lsu_is_valid),
    .set_lr_addr(csr_set_lr_addr),
    .lsu_addr(csr_lsu_addr),
    .perfCntCondMultiCommit(csr_perfCntCondMultiCommit),
    .set_lr_val(csr_set_lr_val),
    .lrAddr_0(csr_lrAddr_0)
  );
  ysyx_210000_MOU mou ( // @[EXU.scala 85:19]
    .io_in_valid(mou_io_in_valid),
    .io_in_bits_func(mou_io_in_bits_func),
    .io_cfIn_pc(mou_io_cfIn_pc),
    .io_redirect_target(mou_io_redirect_target),
    .io_redirect_valid(mou_io_redirect_valid),
    .flushICache_0(mou_flushICache_0),
    .flushTLB_0(mou_flushTLB_0)
  );
  assign io__in_ready = ~io__in_valid | io__out_valid; // @[EXU.scala 118:31]
  assign io__out_valid = io__in_valid & _T_57; // @[EXU.scala 107:31]
  assign io__out_bits_decode_cf_pc = io__in_bits_cf_pc; // @[EXU.scala 97:28]
  assign io__out_bits_decode_cf_redirect_target = mou_io_redirect_valid ? mou_io_redirect_target : _T_42_target; // @[EXU.scala 100:8]
  assign io__out_bits_decode_cf_redirect_valid = mou_io_redirect_valid ? mou_io_redirect_valid : _T_42_valid; // @[EXU.scala 100:8]
  assign io__out_bits_decode_ctrl_fuType = io__in_bits_ctrl_fuType; // @[EXU.scala 95:14]
  assign io__out_bits_decode_ctrl_rfWen = io__in_bits_ctrl_rfWen & (~lsuTlbPF & ~lsu_io__loadAddrMisaligned & ~
    lsu_io__storeAddrMisaligned | ~fuValids_1) & ~(csr_io_wenFix & fuValids_3); // @[EXU.scala 93:125]
  assign io__out_bits_decode_ctrl_rfDest = io__in_bits_ctrl_rfDest; // @[EXU.scala 94:14]
  assign io__out_bits_commits_0 = alu_io__out_bits; // @[EXU.scala 112:35]
  assign io__out_bits_commits_1 = lsu_io__out_bits; // @[EXU.scala 113:35]
  assign io__out_bits_commits_2 = mdu_io_out_bits; // @[EXU.scala 115:35]
  assign io__out_bits_commits_3 = csr_io_out_bits; // @[EXU.scala 114:35]
  assign io__dmem_req_valid = lsu_io__dmem_req_valid; // @[EXU.scala 60:11]
  assign io__dmem_req_bits_addr = lsu_io__dmem_req_bits_addr; // @[EXU.scala 60:11]
  assign io__dmem_req_bits_size = lsu_io__dmem_req_bits_size; // @[EXU.scala 60:11]
  assign io__dmem_req_bits_cmd = lsu_io__dmem_req_bits_cmd; // @[EXU.scala 60:11]
  assign io__dmem_req_bits_wmask = lsu_io__dmem_req_bits_wmask; // @[EXU.scala 60:11]
  assign io__dmem_req_bits_wdata = lsu_io__dmem_req_bits_wdata; // @[EXU.scala 60:11]
  assign io__forward_valid = io__in_valid; // @[EXU.scala 120:20]
  assign io__forward_wb_rfWen = io__in_bits_ctrl_rfWen; // @[EXU.scala 121:23]
  assign io__forward_wb_rfDest = io__in_bits_ctrl_rfDest; // @[EXU.scala 122:24]
  assign io__forward_wb_rfData = _T_62 ? alu_io__out_bits : lsu_io__out_bits; // @[EXU.scala 123:30]
  assign io__forward_fuType = io__in_bits_ctrl_fuType; // @[EXU.scala 124:21]
  assign io__memMMU_imem_priviledgeMode = csr_io_imemMMU_priviledgeMode; // @[EXU.scala 82:18]
  assign io__memMMU_dmem_priviledgeMode = csr_io_dmemMMU_priviledgeMode; // @[EXU.scala 83:18]
  assign io__memMMU_dmem_status_sum = csr_io_dmemMMU_status_sum; // @[EXU.scala 83:18]
  assign io__memMMU_dmem_status_mxr = csr_io_dmemMMU_status_mxr; // @[EXU.scala 83:18]
  assign flushICache = mou_flushICache_0;
  assign satp = csr_satp_0;
  assign REG_6_valid = alu_REG_6_0_valid;
  assign REG_6_pc = alu_REG_6_0_pc;
  assign REG_6_isMissPredict = alu_REG_6_0_isMissPredict;
  assign REG_6_actualTarget = alu_REG_6_0_actualTarget;
  assign REG_6_actualTaken = alu_REG_6_0_actualTaken;
  assign REG_6_fuOpType = alu_REG_6_0_fuOpType;
  assign REG_6_btbType = alu_REG_6_0_btbType;
  assign REG_6_isRVC = alu_REG_6_0_isRVC;
  assign amoReq = lsu_amoReq_0;
  assign isuPermitLibLoad = csr_isuPermitLibLoad_0;
  assign isuPermitLibStore = csr_isuPermitLibStore_0;
  assign intrVec = csr_intrVec_0;
  assign flushTLB = mou_flushTLB_0;
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io__in_valid = io__in_bits_ctrl_fuType == 3'h0 & io__in_valid & ~io__flush; // @[EXU.scala 43:81]
  assign alu_io__in_bits_src1 = io__in_bits_data_src1; // @[EXU.scala 37:34]
  assign alu_io__in_bits_src2 = io__in_bits_data_src2; // @[EXU.scala 38:34]
  assign alu_io__in_bits_func = io__in_bits_ctrl_fuOpType; // @[ALU.scala 85:15]
  assign alu_io__out_ready = 1'h1; // @[EXU.scala 49:20]
  assign alu_io__cfIn_instr = io__in_bits_cf_instr; // @[EXU.scala 47:15]
  assign alu_io__cfIn_pc = io__in_bits_cf_pc; // @[EXU.scala 47:15]
  assign alu_io__cfIn_pnpc = io__in_bits_cf_pnpc; // @[EXU.scala 47:15]
  assign alu_io__cfIn_brIdx = io__in_bits_cf_brIdx; // @[EXU.scala 47:15]
  assign alu_io__offset = io__in_bits_data_imm; // @[EXU.scala 48:17]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io__in_valid = io__in_bits_ctrl_fuType == 3'h1 & io__in_valid & ~io__flush; // @[EXU.scala 43:81]
  assign lsu_io__in_bits_src1 = io__in_bits_data_src1; // @[EXU.scala 37:34]
  assign lsu_io__in_bits_func = io__in_bits_ctrl_fuOpType; // @[UnpipelinedLSU.scala 44:15]
  assign lsu_io__out_ready = 1'h1; // @[EXU.scala 61:20]
  assign lsu_io__srcSum = io__in_bits_data_addr; // @[EXU.scala 56:17]
  assign lsu_io__wdata = io__in_bits_data_src2; // @[EXU.scala 38:34]
  assign lsu_io__instr = io__in_bits_cf_instr[31:0]; // @[EXU.scala 58:16]
  assign lsu_io__dmem_req_ready = io__dmem_req_ready; // @[EXU.scala 60:11]
  assign lsu_io__dmem_resp_valid = io__dmem_resp_valid; // @[EXU.scala 60:11]
  assign lsu_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[EXU.scala 60:11]
  assign lsu_DTLBPF = _T_28_0;
  assign lsu_cannot_access_memory = csr_lsuDeny_0;
  assign lsu_DTLBENABLE = vmEnable;
  assign lsu_DTLBFINISH = _T_27_0;
  assign lsu_lr_addr = csr_lrAddr_0;
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_in_valid = io__in_bits_ctrl_fuType == 3'h2 & io__in_valid & ~io__flush; // @[EXU.scala 43:81]
  assign mdu_io_in_bits_src1 = io__in_bits_data_src1; // @[EXU.scala 37:34]
  assign mdu_io_in_bits_src2 = io__in_bits_data_src2; // @[EXU.scala 38:34]
  assign mdu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[MDU.scala 73:15]
  assign mdu_io_out_ready = 1'h1; // @[EXU.scala 65:20]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_in_valid = io__in_bits_ctrl_fuType == 3'h3 & io__in_valid & ~io__flush; // @[EXU.scala 43:81]
  assign csr_io_in_bits_src1 = io__in_bits_data_src1; // @[EXU.scala 37:34]
  assign csr_io_in_bits_src2 = io__in_bits_data_src2; // @[EXU.scala 38:34]
  assign csr_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[CSR.scala 235:15]
  assign csr_io_out_ready = 1'h1; // @[EXU.scala 80:20]
  assign csr_io_cfIn_instr = io__in_bits_cf_instr; // @[EXU.scala 70:15]
  assign csr_io_cfIn_pc = io__in_bits_cf_pc; // @[EXU.scala 70:15]
  assign csr_io_cfIn_exceptionVec_1 = io__in_bits_cf_exceptionVec_1; // @[EXU.scala 70:15]
  assign csr_io_cfIn_exceptionVec_2 = io__in_bits_cf_exceptionVec_2; // @[EXU.scala 70:15]
  assign csr_io_cfIn_exceptionVec_4 = lsu_io__loadAddrMisaligned; // @[EXU.scala 71:48]
  assign csr_io_cfIn_exceptionVec_6 = lsu_io__storeAddrMisaligned; // @[EXU.scala 72:49]
  assign csr_io_cfIn_exceptionVec_12 = io__in_bits_cf_exceptionVec_12; // @[EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_0 = io__in_bits_cf_intrVec_0; // @[EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_1 = io__in_bits_cf_intrVec_1; // @[EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_2 = io__in_bits_cf_intrVec_2; // @[EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_3 = io__in_bits_cf_intrVec_3; // @[EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_4 = io__in_bits_cf_intrVec_4; // @[EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_5 = io__in_bits_cf_intrVec_5; // @[EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_6 = io__in_bits_cf_intrVec_6; // @[EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_7 = io__in_bits_cf_intrVec_7; // @[EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_8 = io__in_bits_cf_intrVec_8; // @[EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_9 = io__in_bits_cf_intrVec_9; // @[EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_10 = io__in_bits_cf_intrVec_10; // @[EXU.scala 70:15]
  assign csr_io_cfIn_intrVec_11 = io__in_bits_cf_intrVec_11; // @[EXU.scala 70:15]
  assign csr_io_cfIn_crossPageIPFFix = io__in_bits_cf_crossPageIPFFix; // @[EXU.scala 70:15]
  assign csr_io_instrValid = io__in_valid & _T_2; // @[EXU.scala 73:36]
  assign csr_io_lsuIsLoad = io__in_bits_ctrl_lsuIsLoad; // @[EXU.scala 75:20]
  assign csr_io_lsuPermitLibLoad = io__in_bits_ctrl_permitLibLoad; // @[EXU.scala 76:27]
  assign csr_io_lsuPermitLibStore = io__in_bits_ctrl_permitLibStore; // @[EXU.scala 77:28]
  assign csr_io_dmemMMU_loadPF = io__memMMU_dmem_loadPF; // @[EXU.scala 83:18]
  assign csr_io_dmemMMU_storePF = io__memMMU_dmem_storePF; // @[EXU.scala 83:18]
  assign csr_io_dmemMMU_addr = io__memMMU_dmem_addr; // @[EXU.scala 83:18]
  assign csr_set_lr = lsu_setLr_0;
  assign csr_is_pulpret = alu__T_113_0;
  assign csr_perfCntCondMinstret = io_in_valid;
  assign csr_mtip_0 = io_extra_mtip;
  assign csr_meip_0 = io_extra_meip_0;
  assign csr_redirect_valid = alu_io_redirect_valid;
  assign csr_isu_addr = isuAddr;
  assign csr_redirect_target = alu_io_redirect_target;
  assign csr_LSUEXECADDR = lsu_io_in_bits_src1;
  assign csr_msip_0 = io_extra_msip;
  assign csr_lsu_is_valid = lsu__T_20_0;
  assign csr_set_lr_addr = lsu_setLrAddr_0;
  assign csr_lsu_addr = lsu__T_28_0;
  assign csr_perfCntCondMultiCommit = falseWire;
  assign csr_set_lr_val = lsu_setLrVal_0;
  assign mou_io_in_valid = io__in_bits_ctrl_fuType == 3'h4 & io__in_valid & ~io__flush; // @[EXU.scala 43:81]
  assign mou_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[MOU.scala 45:15]
  assign mou_io_cfIn_pc = io__in_bits_cf_pc; // @[EXU.scala 88:15]
endmodule
module ysyx_210000_WBU(
  input         io__in_valid,
  input  [38:0] io__in_bits_decode_cf_pc,
  input  [38:0] io__in_bits_decode_cf_redirect_target,
  input         io__in_bits_decode_cf_redirect_valid,
  input  [2:0]  io__in_bits_decode_ctrl_fuType,
  input         io__in_bits_decode_ctrl_rfWen,
  input  [4:0]  io__in_bits_decode_ctrl_rfDest,
  input  [63:0] io__in_bits_commits_0,
  input  [63:0] io__in_bits_commits_1,
  input  [63:0] io__in_bits_commits_2,
  input  [63:0] io__in_bits_commits_3,
  output        io__wb_rfWen,
  output [4:0]  io__wb_rfDest,
  output [63:0] io__wb_rfData,
  output [38:0] io__redirect_target,
  output        io__redirect_valid,
  output        io_in_valid,
  output        falseWire_0
);
  wire [63:0] _GEN_1 = 3'h1 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_1 : io__in_bits_commits_0; // @[WBU.scala 33:16 WBU.scala 33:16]
  wire [63:0] _GEN_2 = 3'h2 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_2 : _GEN_1; // @[WBU.scala 33:16 WBU.scala 33:16]
  wire [63:0] _GEN_3 = 3'h3 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_3 : _GEN_2; // @[WBU.scala 33:16 WBU.scala 33:16]
  wire  falseWire = 1'h0;
  assign io__wb_rfWen = io__in_bits_decode_ctrl_rfWen & io__in_valid; // @[WBU.scala 31:47]
  assign io__wb_rfDest = io__in_bits_decode_ctrl_rfDest; // @[WBU.scala 32:16]
  assign io__wb_rfData = 3'h4 == io__in_bits_decode_ctrl_fuType ? 64'h0 : _GEN_3; // @[WBU.scala 33:16 WBU.scala 33:16]
  assign io__redirect_target = io__in_bits_decode_cf_redirect_target; // @[WBU.scala 37:15]
  assign io__redirect_valid = io__in_bits_decode_cf_redirect_valid & io__in_valid; // @[WBU.scala 38:60]
  assign io_in_valid = io__in_valid;
  assign falseWire_0 = 1'h0;
endmodule
module ysyx_210000_Backend_inorder(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_cf_instr,
  input  [38:0] io_in_0_bits_cf_pc,
  input  [38:0] io_in_0_bits_cf_pnpc,
  input         io_in_0_bits_cf_exceptionVec_1,
  input         io_in_0_bits_cf_exceptionVec_2,
  input         io_in_0_bits_cf_exceptionVec_12,
  input         io_in_0_bits_cf_intrVec_0,
  input         io_in_0_bits_cf_intrVec_1,
  input         io_in_0_bits_cf_intrVec_2,
  input         io_in_0_bits_cf_intrVec_3,
  input         io_in_0_bits_cf_intrVec_4,
  input         io_in_0_bits_cf_intrVec_5,
  input         io_in_0_bits_cf_intrVec_6,
  input         io_in_0_bits_cf_intrVec_7,
  input         io_in_0_bits_cf_intrVec_8,
  input         io_in_0_bits_cf_intrVec_9,
  input         io_in_0_bits_cf_intrVec_10,
  input         io_in_0_bits_cf_intrVec_11,
  input  [3:0]  io_in_0_bits_cf_brIdx,
  input         io_in_0_bits_cf_crossPageIPFFix,
  input         io_in_0_bits_ctrl_src1Type,
  input         io_in_0_bits_ctrl_src2Type,
  input  [2:0]  io_in_0_bits_ctrl_fuType,
  input  [6:0]  io_in_0_bits_ctrl_fuOpType,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2,
  input         io_in_0_bits_ctrl_rfWen,
  input  [4:0]  io_in_0_bits_ctrl_rfDest,
  input  [63:0] io_in_0_bits_data_imm,
  input  [1:0]  io_flush,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [38:0] io_dmem_req_bits_addr,
  output [2:0]  io_dmem_req_bits_size,
  output [3:0]  io_dmem_req_bits_cmd,
  output [7:0]  io_dmem_req_bits_wmask,
  output [63:0] io_dmem_req_bits_wdata,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  output [1:0]  io_memMMU_imem_priviledgeMode,
  output [1:0]  io_memMMU_dmem_priviledgeMode,
  output        io_memMMU_dmem_status_sum,
  output        io_memMMU_dmem_status_mxr,
  input         io_memMMU_dmem_loadPF,
  input         io_memMMU_dmem_storePF,
  input  [38:0] io_memMMU_dmem_addr,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input         _T_28,
  output        flushICache,
  output [63:0] satp,
  output        REG_6_valid,
  output [38:0] REG_6_pc,
  output        REG_6_isMissPredict,
  output [38:0] REG_6_actualTarget,
  output        REG_6_actualTaken,
  output [6:0]  REG_6_fuOpType,
  output [1:0]  REG_6_btbType,
  output        REG_6_isRVC,
  input         io_extra_mtip,
  output        amoReq,
  input         io_extra_meip_0,
  input         vmEnable,
  output [11:0] intrVec,
  input         _T_27,
  input         io_extra_msip,
  output        flushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
`endif // RANDOMIZE_REG_INIT
  wire  isu_clock; // @[Backend.scala 675:20]
  wire  isu_reset; // @[Backend.scala 675:20]
  wire  isu_io_in_0_ready; // @[Backend.scala 675:20]
  wire  isu_io_in_0_valid; // @[Backend.scala 675:20]
  wire [63:0] isu_io_in_0_bits_cf_instr; // @[Backend.scala 675:20]
  wire [38:0] isu_io_in_0_bits_cf_pc; // @[Backend.scala 675:20]
  wire [38:0] isu_io_in_0_bits_cf_pnpc; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_1; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_2; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_12; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_0; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_1; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_2; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_3; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_4; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_5; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_6; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_7; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_8; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_9; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_10; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_11; // @[Backend.scala 675:20]
  wire [3:0] isu_io_in_0_bits_cf_brIdx; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_crossPageIPFFix; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_ctrl_src1Type; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_ctrl_src2Type; // @[Backend.scala 675:20]
  wire [2:0] isu_io_in_0_bits_ctrl_fuType; // @[Backend.scala 675:20]
  wire [6:0] isu_io_in_0_bits_ctrl_fuOpType; // @[Backend.scala 675:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc1; // @[Backend.scala 675:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc2; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_ctrl_rfWen; // @[Backend.scala 675:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfDest; // @[Backend.scala 675:20]
  wire [63:0] isu_io_in_0_bits_data_imm; // @[Backend.scala 675:20]
  wire  isu_io_out_ready; // @[Backend.scala 675:20]
  wire  isu_io_out_valid; // @[Backend.scala 675:20]
  wire [63:0] isu_io_out_bits_cf_instr; // @[Backend.scala 675:20]
  wire [38:0] isu_io_out_bits_cf_pc; // @[Backend.scala 675:20]
  wire [38:0] isu_io_out_bits_cf_pnpc; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_exceptionVec_1; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_exceptionVec_2; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_exceptionVec_12; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_0; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_1; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_2; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_3; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_4; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_5; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_6; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_7; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_8; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_9; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_10; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_11; // @[Backend.scala 675:20]
  wire [3:0] isu_io_out_bits_cf_brIdx; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_crossPageIPFFix; // @[Backend.scala 675:20]
  wire [2:0] isu_io_out_bits_ctrl_fuType; // @[Backend.scala 675:20]
  wire [6:0] isu_io_out_bits_ctrl_fuOpType; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_ctrl_rfWen; // @[Backend.scala 675:20]
  wire [4:0] isu_io_out_bits_ctrl_rfDest; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_ctrl_permitLibLoad; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_ctrl_permitLibStore; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_ctrl_lsuIsLoad; // @[Backend.scala 675:20]
  wire [63:0] isu_io_out_bits_data_src1; // @[Backend.scala 675:20]
  wire [63:0] isu_io_out_bits_data_src2; // @[Backend.scala 675:20]
  wire [63:0] isu_io_out_bits_data_imm; // @[Backend.scala 675:20]
  wire [63:0] isu_io_out_bits_data_addr; // @[Backend.scala 675:20]
  wire  isu_io_wb_rfWen; // @[Backend.scala 675:20]
  wire [4:0] isu_io_wb_rfDest; // @[Backend.scala 675:20]
  wire [63:0] isu_io_wb_rfData; // @[Backend.scala 675:20]
  wire  isu_io_forward_valid; // @[Backend.scala 675:20]
  wire  isu_io_forward_wb_rfWen; // @[Backend.scala 675:20]
  wire [4:0] isu_io_forward_wb_rfDest; // @[Backend.scala 675:20]
  wire [63:0] isu_io_forward_wb_rfData; // @[Backend.scala 675:20]
  wire [2:0] isu_io_forward_fuType; // @[Backend.scala 675:20]
  wire  isu_io_flush; // @[Backend.scala 675:20]
  wire [63:0] isu_isuAddr_0; // @[Backend.scala 675:20]
  wire  isu_isu_perm_lib_ld; // @[Backend.scala 675:20]
  wire  isu_isu_perm_lib_st; // @[Backend.scala 675:20]
  wire  exu_clock; // @[Backend.scala 676:20]
  wire  exu_reset; // @[Backend.scala 676:20]
  wire  exu_io__in_ready; // @[Backend.scala 676:20]
  wire  exu_io__in_valid; // @[Backend.scala 676:20]
  wire [63:0] exu_io__in_bits_cf_instr; // @[Backend.scala 676:20]
  wire [38:0] exu_io__in_bits_cf_pc; // @[Backend.scala 676:20]
  wire [38:0] exu_io__in_bits_cf_pnpc; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_exceptionVec_1; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_exceptionVec_2; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_exceptionVec_12; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_0; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_1; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_2; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_3; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_4; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_5; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_6; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_7; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_8; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_9; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_10; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_11; // @[Backend.scala 676:20]
  wire [3:0] exu_io__in_bits_cf_brIdx; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_crossPageIPFFix; // @[Backend.scala 676:20]
  wire [2:0] exu_io__in_bits_ctrl_fuType; // @[Backend.scala 676:20]
  wire [6:0] exu_io__in_bits_ctrl_fuOpType; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_ctrl_rfWen; // @[Backend.scala 676:20]
  wire [4:0] exu_io__in_bits_ctrl_rfDest; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_ctrl_permitLibLoad; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_ctrl_permitLibStore; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_ctrl_lsuIsLoad; // @[Backend.scala 676:20]
  wire [63:0] exu_io__in_bits_data_src1; // @[Backend.scala 676:20]
  wire [63:0] exu_io__in_bits_data_src2; // @[Backend.scala 676:20]
  wire [63:0] exu_io__in_bits_data_imm; // @[Backend.scala 676:20]
  wire [63:0] exu_io__in_bits_data_addr; // @[Backend.scala 676:20]
  wire  exu_io__out_ready; // @[Backend.scala 676:20]
  wire  exu_io__out_valid; // @[Backend.scala 676:20]
  wire [38:0] exu_io__out_bits_decode_cf_pc; // @[Backend.scala 676:20]
  wire [38:0] exu_io__out_bits_decode_cf_redirect_target; // @[Backend.scala 676:20]
  wire  exu_io__out_bits_decode_cf_redirect_valid; // @[Backend.scala 676:20]
  wire [2:0] exu_io__out_bits_decode_ctrl_fuType; // @[Backend.scala 676:20]
  wire  exu_io__out_bits_decode_ctrl_rfWen; // @[Backend.scala 676:20]
  wire [4:0] exu_io__out_bits_decode_ctrl_rfDest; // @[Backend.scala 676:20]
  wire [63:0] exu_io__out_bits_commits_0; // @[Backend.scala 676:20]
  wire [63:0] exu_io__out_bits_commits_1; // @[Backend.scala 676:20]
  wire [63:0] exu_io__out_bits_commits_2; // @[Backend.scala 676:20]
  wire [63:0] exu_io__out_bits_commits_3; // @[Backend.scala 676:20]
  wire  exu_io__flush; // @[Backend.scala 676:20]
  wire  exu_io__dmem_req_ready; // @[Backend.scala 676:20]
  wire  exu_io__dmem_req_valid; // @[Backend.scala 676:20]
  wire [38:0] exu_io__dmem_req_bits_addr; // @[Backend.scala 676:20]
  wire [2:0] exu_io__dmem_req_bits_size; // @[Backend.scala 676:20]
  wire [3:0] exu_io__dmem_req_bits_cmd; // @[Backend.scala 676:20]
  wire [7:0] exu_io__dmem_req_bits_wmask; // @[Backend.scala 676:20]
  wire [63:0] exu_io__dmem_req_bits_wdata; // @[Backend.scala 676:20]
  wire  exu_io__dmem_resp_valid; // @[Backend.scala 676:20]
  wire [63:0] exu_io__dmem_resp_bits_rdata; // @[Backend.scala 676:20]
  wire  exu_io__forward_valid; // @[Backend.scala 676:20]
  wire  exu_io__forward_wb_rfWen; // @[Backend.scala 676:20]
  wire [4:0] exu_io__forward_wb_rfDest; // @[Backend.scala 676:20]
  wire [63:0] exu_io__forward_wb_rfData; // @[Backend.scala 676:20]
  wire [2:0] exu_io__forward_fuType; // @[Backend.scala 676:20]
  wire [1:0] exu_io__memMMU_imem_priviledgeMode; // @[Backend.scala 676:20]
  wire [1:0] exu_io__memMMU_dmem_priviledgeMode; // @[Backend.scala 676:20]
  wire  exu_io__memMMU_dmem_status_sum; // @[Backend.scala 676:20]
  wire  exu_io__memMMU_dmem_status_mxr; // @[Backend.scala 676:20]
  wire  exu_io__memMMU_dmem_loadPF; // @[Backend.scala 676:20]
  wire  exu_io__memMMU_dmem_storePF; // @[Backend.scala 676:20]
  wire [38:0] exu_io__memMMU_dmem_addr; // @[Backend.scala 676:20]
  wire  exu__T_28_0; // @[Backend.scala 676:20]
  wire  exu_flushICache; // @[Backend.scala 676:20]
  wire [63:0] exu_satp; // @[Backend.scala 676:20]
  wire  exu_REG_6_valid; // @[Backend.scala 676:20]
  wire [38:0] exu_REG_6_pc; // @[Backend.scala 676:20]
  wire  exu_REG_6_isMissPredict; // @[Backend.scala 676:20]
  wire [38:0] exu_REG_6_actualTarget; // @[Backend.scala 676:20]
  wire  exu_REG_6_actualTaken; // @[Backend.scala 676:20]
  wire [6:0] exu_REG_6_fuOpType; // @[Backend.scala 676:20]
  wire [1:0] exu_REG_6_btbType; // @[Backend.scala 676:20]
  wire  exu_REG_6_isRVC; // @[Backend.scala 676:20]
  wire  exu_io_in_valid; // @[Backend.scala 676:20]
  wire  exu_io_extra_mtip; // @[Backend.scala 676:20]
  wire  exu_amoReq; // @[Backend.scala 676:20]
  wire  exu_io_extra_meip_0; // @[Backend.scala 676:20]
  wire  exu_vmEnable; // @[Backend.scala 676:20]
  wire [63:0] exu_isuAddr; // @[Backend.scala 676:20]
  wire  exu_isuPermitLibLoad; // @[Backend.scala 676:20]
  wire  exu_isuPermitLibStore; // @[Backend.scala 676:20]
  wire [11:0] exu_intrVec; // @[Backend.scala 676:20]
  wire  exu__T_27_0; // @[Backend.scala 676:20]
  wire  exu_io_extra_msip; // @[Backend.scala 676:20]
  wire  exu_flushTLB; // @[Backend.scala 676:20]
  wire  exu_falseWire; // @[Backend.scala 676:20]
  wire  wbu_io__in_valid; // @[Backend.scala 677:20]
  wire [38:0] wbu_io__in_bits_decode_cf_pc; // @[Backend.scala 677:20]
  wire [38:0] wbu_io__in_bits_decode_cf_redirect_target; // @[Backend.scala 677:20]
  wire  wbu_io__in_bits_decode_cf_redirect_valid; // @[Backend.scala 677:20]
  wire [2:0] wbu_io__in_bits_decode_ctrl_fuType; // @[Backend.scala 677:20]
  wire  wbu_io__in_bits_decode_ctrl_rfWen; // @[Backend.scala 677:20]
  wire [4:0] wbu_io__in_bits_decode_ctrl_rfDest; // @[Backend.scala 677:20]
  wire [63:0] wbu_io__in_bits_commits_0; // @[Backend.scala 677:20]
  wire [63:0] wbu_io__in_bits_commits_1; // @[Backend.scala 677:20]
  wire [63:0] wbu_io__in_bits_commits_2; // @[Backend.scala 677:20]
  wire [63:0] wbu_io__in_bits_commits_3; // @[Backend.scala 677:20]
  wire  wbu_io__wb_rfWen; // @[Backend.scala 677:20]
  wire [4:0] wbu_io__wb_rfDest; // @[Backend.scala 677:20]
  wire [63:0] wbu_io__wb_rfData; // @[Backend.scala 677:20]
  wire [38:0] wbu_io__redirect_target; // @[Backend.scala 677:20]
  wire  wbu_io__redirect_valid; // @[Backend.scala 677:20]
  wire  wbu_io_in_valid; // @[Backend.scala 677:20]
  wire  wbu_falseWire_0; // @[Backend.scala 677:20]
  wire  _T = exu_io__out_ready & exu_io__out_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : REG; // @[Pipeline.scala 25:25 Pipeline.scala 25:33 Pipeline.scala 24:24]
  wire  _T_2 = isu_io_out_valid & exu_io__in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = isu_io_out_valid & exu_io__in_ready | _GEN_0; // @[Pipeline.scala 26:38 Pipeline.scala 26:46]
  reg [63:0] REG_1_cf_instr; // @[Reg.scala 27:20]
  reg [38:0] REG_1_cf_pc; // @[Reg.scala 27:20]
  reg [38:0] REG_1_cf_pnpc; // @[Reg.scala 27:20]
  reg  REG_1_cf_exceptionVec_1; // @[Reg.scala 27:20]
  reg  REG_1_cf_exceptionVec_2; // @[Reg.scala 27:20]
  reg  REG_1_cf_exceptionVec_12; // @[Reg.scala 27:20]
  reg  REG_1_cf_intrVec_0; // @[Reg.scala 27:20]
  reg  REG_1_cf_intrVec_1; // @[Reg.scala 27:20]
  reg  REG_1_cf_intrVec_2; // @[Reg.scala 27:20]
  reg  REG_1_cf_intrVec_3; // @[Reg.scala 27:20]
  reg  REG_1_cf_intrVec_4; // @[Reg.scala 27:20]
  reg  REG_1_cf_intrVec_5; // @[Reg.scala 27:20]
  reg  REG_1_cf_intrVec_6; // @[Reg.scala 27:20]
  reg  REG_1_cf_intrVec_7; // @[Reg.scala 27:20]
  reg  REG_1_cf_intrVec_8; // @[Reg.scala 27:20]
  reg  REG_1_cf_intrVec_9; // @[Reg.scala 27:20]
  reg  REG_1_cf_intrVec_10; // @[Reg.scala 27:20]
  reg  REG_1_cf_intrVec_11; // @[Reg.scala 27:20]
  reg [3:0] REG_1_cf_brIdx; // @[Reg.scala 27:20]
  reg  REG_1_cf_crossPageIPFFix; // @[Reg.scala 27:20]
  reg [2:0] REG_1_ctrl_fuType; // @[Reg.scala 27:20]
  reg [6:0] REG_1_ctrl_fuOpType; // @[Reg.scala 27:20]
  reg  REG_1_ctrl_rfWen; // @[Reg.scala 27:20]
  reg [4:0] REG_1_ctrl_rfDest; // @[Reg.scala 27:20]
  reg  REG_1_ctrl_permitLibLoad; // @[Reg.scala 27:20]
  reg  REG_1_ctrl_permitLibStore; // @[Reg.scala 27:20]
  reg  REG_1_ctrl_lsuIsLoad; // @[Reg.scala 27:20]
  reg [63:0] REG_1_data_src1; // @[Reg.scala 27:20]
  reg [63:0] REG_1_data_src2; // @[Reg.scala 27:20]
  reg [63:0] REG_1_data_imm; // @[Reg.scala 27:20]
  reg [63:0] REG_1_data_addr; // @[Reg.scala 27:20]
  reg  REG_2; // @[Pipeline.scala 24:24]
  wire  _T_5 = exu_io__out_valid; // @[Pipeline.scala 26:22]
  reg [38:0] REG_3_decode_cf_pc; // @[Reg.scala 27:20]
  reg [38:0] REG_3_decode_cf_redirect_target; // @[Reg.scala 27:20]
  reg  REG_3_decode_cf_redirect_valid; // @[Reg.scala 27:20]
  reg [2:0] REG_3_decode_ctrl_fuType; // @[Reg.scala 27:20]
  reg  REG_3_decode_ctrl_rfWen; // @[Reg.scala 27:20]
  reg [4:0] REG_3_decode_ctrl_rfDest; // @[Reg.scala 27:20]
  reg [63:0] REG_3_commits_0; // @[Reg.scala 27:20]
  reg [63:0] REG_3_commits_1; // @[Reg.scala 27:20]
  reg [63:0] REG_3_commits_2; // @[Reg.scala 27:20]
  reg [63:0] REG_3_commits_3; // @[Reg.scala 27:20]
  ysyx_210000_ISU isu ( // @[Backend.scala 675:20]
    .clock(isu_clock),
    .reset(isu_reset),
    .io_in_0_ready(isu_io_in_0_ready),
    .io_in_0_valid(isu_io_in_0_valid),
    .io_in_0_bits_cf_instr(isu_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(isu_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(isu_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(isu_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(isu_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(isu_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_0(isu_io_in_0_bits_cf_intrVec_0),
    .io_in_0_bits_cf_intrVec_1(isu_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_2(isu_io_in_0_bits_cf_intrVec_2),
    .io_in_0_bits_cf_intrVec_3(isu_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_4(isu_io_in_0_bits_cf_intrVec_4),
    .io_in_0_bits_cf_intrVec_5(isu_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_6(isu_io_in_0_bits_cf_intrVec_6),
    .io_in_0_bits_cf_intrVec_7(isu_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_8(isu_io_in_0_bits_cf_intrVec_8),
    .io_in_0_bits_cf_intrVec_9(isu_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_10(isu_io_in_0_bits_cf_intrVec_10),
    .io_in_0_bits_cf_intrVec_11(isu_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(isu_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossPageIPFFix(isu_io_in_0_bits_cf_crossPageIPFFix),
    .io_in_0_bits_ctrl_src1Type(isu_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(isu_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(isu_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(isu_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(isu_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(isu_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(isu_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(isu_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_data_imm(isu_io_in_0_bits_data_imm),
    .io_out_ready(isu_io_out_ready),
    .io_out_valid(isu_io_out_valid),
    .io_out_bits_cf_instr(isu_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(isu_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(isu_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(isu_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(isu_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(isu_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_0(isu_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(isu_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(isu_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(isu_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(isu_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(isu_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(isu_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(isu_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(isu_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(isu_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(isu_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(isu_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(isu_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossPageIPFFix(isu_io_out_bits_cf_crossPageIPFFix),
    .io_out_bits_ctrl_fuType(isu_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(isu_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfWen(isu_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(isu_io_out_bits_ctrl_rfDest),
    .io_out_bits_ctrl_permitLibLoad(isu_io_out_bits_ctrl_permitLibLoad),
    .io_out_bits_ctrl_permitLibStore(isu_io_out_bits_ctrl_permitLibStore),
    .io_out_bits_ctrl_lsuIsLoad(isu_io_out_bits_ctrl_lsuIsLoad),
    .io_out_bits_data_src1(isu_io_out_bits_data_src1),
    .io_out_bits_data_src2(isu_io_out_bits_data_src2),
    .io_out_bits_data_imm(isu_io_out_bits_data_imm),
    .io_out_bits_data_addr(isu_io_out_bits_data_addr),
    .io_wb_rfWen(isu_io_wb_rfWen),
    .io_wb_rfDest(isu_io_wb_rfDest),
    .io_wb_rfData(isu_io_wb_rfData),
    .io_forward_valid(isu_io_forward_valid),
    .io_forward_wb_rfWen(isu_io_forward_wb_rfWen),
    .io_forward_wb_rfDest(isu_io_forward_wb_rfDest),
    .io_forward_wb_rfData(isu_io_forward_wb_rfData),
    .io_forward_fuType(isu_io_forward_fuType),
    .io_flush(isu_io_flush),
    .isuAddr_0(isu_isuAddr_0),
    .isu_perm_lib_ld(isu_isu_perm_lib_ld),
    .isu_perm_lib_st(isu_isu_perm_lib_st)
  );
  ysyx_210000_EXU exu ( // @[Backend.scala 676:20]
    .clock(exu_clock),
    .reset(exu_reset),
    .io__in_ready(exu_io__in_ready),
    .io__in_valid(exu_io__in_valid),
    .io__in_bits_cf_instr(exu_io__in_bits_cf_instr),
    .io__in_bits_cf_pc(exu_io__in_bits_cf_pc),
    .io__in_bits_cf_pnpc(exu_io__in_bits_cf_pnpc),
    .io__in_bits_cf_exceptionVec_1(exu_io__in_bits_cf_exceptionVec_1),
    .io__in_bits_cf_exceptionVec_2(exu_io__in_bits_cf_exceptionVec_2),
    .io__in_bits_cf_exceptionVec_12(exu_io__in_bits_cf_exceptionVec_12),
    .io__in_bits_cf_intrVec_0(exu_io__in_bits_cf_intrVec_0),
    .io__in_bits_cf_intrVec_1(exu_io__in_bits_cf_intrVec_1),
    .io__in_bits_cf_intrVec_2(exu_io__in_bits_cf_intrVec_2),
    .io__in_bits_cf_intrVec_3(exu_io__in_bits_cf_intrVec_3),
    .io__in_bits_cf_intrVec_4(exu_io__in_bits_cf_intrVec_4),
    .io__in_bits_cf_intrVec_5(exu_io__in_bits_cf_intrVec_5),
    .io__in_bits_cf_intrVec_6(exu_io__in_bits_cf_intrVec_6),
    .io__in_bits_cf_intrVec_7(exu_io__in_bits_cf_intrVec_7),
    .io__in_bits_cf_intrVec_8(exu_io__in_bits_cf_intrVec_8),
    .io__in_bits_cf_intrVec_9(exu_io__in_bits_cf_intrVec_9),
    .io__in_bits_cf_intrVec_10(exu_io__in_bits_cf_intrVec_10),
    .io__in_bits_cf_intrVec_11(exu_io__in_bits_cf_intrVec_11),
    .io__in_bits_cf_brIdx(exu_io__in_bits_cf_brIdx),
    .io__in_bits_cf_crossPageIPFFix(exu_io__in_bits_cf_crossPageIPFFix),
    .io__in_bits_ctrl_fuType(exu_io__in_bits_ctrl_fuType),
    .io__in_bits_ctrl_fuOpType(exu_io__in_bits_ctrl_fuOpType),
    .io__in_bits_ctrl_rfWen(exu_io__in_bits_ctrl_rfWen),
    .io__in_bits_ctrl_rfDest(exu_io__in_bits_ctrl_rfDest),
    .io__in_bits_ctrl_permitLibLoad(exu_io__in_bits_ctrl_permitLibLoad),
    .io__in_bits_ctrl_permitLibStore(exu_io__in_bits_ctrl_permitLibStore),
    .io__in_bits_ctrl_lsuIsLoad(exu_io__in_bits_ctrl_lsuIsLoad),
    .io__in_bits_data_src1(exu_io__in_bits_data_src1),
    .io__in_bits_data_src2(exu_io__in_bits_data_src2),
    .io__in_bits_data_imm(exu_io__in_bits_data_imm),
    .io__in_bits_data_addr(exu_io__in_bits_data_addr),
    .io__out_ready(exu_io__out_ready),
    .io__out_valid(exu_io__out_valid),
    .io__out_bits_decode_cf_pc(exu_io__out_bits_decode_cf_pc),
    .io__out_bits_decode_cf_redirect_target(exu_io__out_bits_decode_cf_redirect_target),
    .io__out_bits_decode_cf_redirect_valid(exu_io__out_bits_decode_cf_redirect_valid),
    .io__out_bits_decode_ctrl_fuType(exu_io__out_bits_decode_ctrl_fuType),
    .io__out_bits_decode_ctrl_rfWen(exu_io__out_bits_decode_ctrl_rfWen),
    .io__out_bits_decode_ctrl_rfDest(exu_io__out_bits_decode_ctrl_rfDest),
    .io__out_bits_commits_0(exu_io__out_bits_commits_0),
    .io__out_bits_commits_1(exu_io__out_bits_commits_1),
    .io__out_bits_commits_2(exu_io__out_bits_commits_2),
    .io__out_bits_commits_3(exu_io__out_bits_commits_3),
    .io__flush(exu_io__flush),
    .io__dmem_req_ready(exu_io__dmem_req_ready),
    .io__dmem_req_valid(exu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(exu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(exu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(exu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(exu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(exu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(exu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(exu_io__dmem_resp_bits_rdata),
    .io__forward_valid(exu_io__forward_valid),
    .io__forward_wb_rfWen(exu_io__forward_wb_rfWen),
    .io__forward_wb_rfDest(exu_io__forward_wb_rfDest),
    .io__forward_wb_rfData(exu_io__forward_wb_rfData),
    .io__forward_fuType(exu_io__forward_fuType),
    .io__memMMU_imem_priviledgeMode(exu_io__memMMU_imem_priviledgeMode),
    .io__memMMU_dmem_priviledgeMode(exu_io__memMMU_dmem_priviledgeMode),
    .io__memMMU_dmem_status_sum(exu_io__memMMU_dmem_status_sum),
    .io__memMMU_dmem_status_mxr(exu_io__memMMU_dmem_status_mxr),
    .io__memMMU_dmem_loadPF(exu_io__memMMU_dmem_loadPF),
    .io__memMMU_dmem_storePF(exu_io__memMMU_dmem_storePF),
    .io__memMMU_dmem_addr(exu_io__memMMU_dmem_addr),
    ._T_28_0(exu__T_28_0),
    .flushICache(exu_flushICache),
    .satp(exu_satp),
    .REG_6_valid(exu_REG_6_valid),
    .REG_6_pc(exu_REG_6_pc),
    .REG_6_isMissPredict(exu_REG_6_isMissPredict),
    .REG_6_actualTarget(exu_REG_6_actualTarget),
    .REG_6_actualTaken(exu_REG_6_actualTaken),
    .REG_6_fuOpType(exu_REG_6_fuOpType),
    .REG_6_btbType(exu_REG_6_btbType),
    .REG_6_isRVC(exu_REG_6_isRVC),
    .io_in_valid(exu_io_in_valid),
    .io_extra_mtip(exu_io_extra_mtip),
    .amoReq(exu_amoReq),
    .io_extra_meip_0(exu_io_extra_meip_0),
    .vmEnable(exu_vmEnable),
    .isuAddr(exu_isuAddr),
    .isuPermitLibLoad(exu_isuPermitLibLoad),
    .isuPermitLibStore(exu_isuPermitLibStore),
    .intrVec(exu_intrVec),
    ._T_27_0(exu__T_27_0),
    .io_extra_msip(exu_io_extra_msip),
    .flushTLB(exu_flushTLB),
    .falseWire(exu_falseWire)
  );
  ysyx_210000_WBU wbu ( // @[Backend.scala 677:20]
    .io__in_valid(wbu_io__in_valid),
    .io__in_bits_decode_cf_pc(wbu_io__in_bits_decode_cf_pc),
    .io__in_bits_decode_cf_redirect_target(wbu_io__in_bits_decode_cf_redirect_target),
    .io__in_bits_decode_cf_redirect_valid(wbu_io__in_bits_decode_cf_redirect_valid),
    .io__in_bits_decode_ctrl_fuType(wbu_io__in_bits_decode_ctrl_fuType),
    .io__in_bits_decode_ctrl_rfWen(wbu_io__in_bits_decode_ctrl_rfWen),
    .io__in_bits_decode_ctrl_rfDest(wbu_io__in_bits_decode_ctrl_rfDest),
    .io__in_bits_commits_0(wbu_io__in_bits_commits_0),
    .io__in_bits_commits_1(wbu_io__in_bits_commits_1),
    .io__in_bits_commits_2(wbu_io__in_bits_commits_2),
    .io__in_bits_commits_3(wbu_io__in_bits_commits_3),
    .io__wb_rfWen(wbu_io__wb_rfWen),
    .io__wb_rfDest(wbu_io__wb_rfDest),
    .io__wb_rfData(wbu_io__wb_rfData),
    .io__redirect_target(wbu_io__redirect_target),
    .io__redirect_valid(wbu_io__redirect_valid),
    .io_in_valid(wbu_io_in_valid),
    .falseWire_0(wbu_falseWire_0)
  );
  assign io_in_0_ready = isu_io_in_0_ready; // @[Backend.scala 682:13]
  assign io_dmem_req_valid = exu_io__dmem_req_valid; // @[Backend.scala 694:11]
  assign io_dmem_req_bits_addr = exu_io__dmem_req_bits_addr; // @[Backend.scala 694:11]
  assign io_dmem_req_bits_size = exu_io__dmem_req_bits_size; // @[Backend.scala 694:11]
  assign io_dmem_req_bits_cmd = exu_io__dmem_req_bits_cmd; // @[Backend.scala 694:11]
  assign io_dmem_req_bits_wmask = exu_io__dmem_req_bits_wmask; // @[Backend.scala 694:11]
  assign io_dmem_req_bits_wdata = exu_io__dmem_req_bits_wdata; // @[Backend.scala 694:11]
  assign io_memMMU_imem_priviledgeMode = exu_io__memMMU_imem_priviledgeMode; // @[Backend.scala 692:18]
  assign io_memMMU_dmem_priviledgeMode = exu_io__memMMU_dmem_priviledgeMode; // @[Backend.scala 693:18]
  assign io_memMMU_dmem_status_sum = exu_io__memMMU_dmem_status_sum; // @[Backend.scala 693:18]
  assign io_memMMU_dmem_status_mxr = exu_io__memMMU_dmem_status_mxr; // @[Backend.scala 693:18]
  assign io_redirect_target = wbu_io__redirect_target; // @[Backend.scala 688:15]
  assign io_redirect_valid = wbu_io__redirect_valid; // @[Backend.scala 688:15]
  assign flushICache = exu_flushICache;
  assign satp = exu_satp;
  assign REG_6_valid = exu_REG_6_valid;
  assign REG_6_pc = exu_REG_6_pc;
  assign REG_6_isMissPredict = exu_REG_6_isMissPredict;
  assign REG_6_actualTarget = exu_REG_6_actualTarget;
  assign REG_6_actualTaken = exu_REG_6_actualTaken;
  assign REG_6_fuOpType = exu_REG_6_fuOpType;
  assign REG_6_btbType = exu_REG_6_btbType;
  assign REG_6_isRVC = exu_REG_6_isRVC;
  assign amoReq = exu_amoReq;
  assign intrVec = exu_intrVec;
  assign flushTLB = exu_flushTLB;
  assign isu_clock = clock;
  assign isu_reset = reset;
  assign isu_io_in_0_valid = io_in_0_valid; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_instr = io_in_0_bits_cf_instr; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_pc = io_in_0_bits_cf_pc; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_0 = io_in_0_bits_cf_intrVec_0; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_2 = io_in_0_bits_cf_intrVec_2; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_4 = io_in_0_bits_cf_intrVec_4; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_6 = io_in_0_bits_cf_intrVec_6; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_8 = io_in_0_bits_cf_intrVec_8; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_10 = io_in_0_bits_cf_intrVec_10; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_crossPageIPFFix = io_in_0_bits_cf_crossPageIPFFix; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_src1Type = io_in_0_bits_ctrl_src1Type; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_src2Type = io_in_0_bits_ctrl_src2Type; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_rfSrc1 = io_in_0_bits_ctrl_rfSrc1; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_rfSrc2 = io_in_0_bits_ctrl_rfSrc2; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_data_imm = io_in_0_bits_data_imm; // @[Backend.scala 682:13]
  assign isu_io_out_ready = exu_io__in_ready; // @[Pipeline.scala 29:16]
  assign isu_io_wb_rfWen = wbu_io__wb_rfWen; // @[Backend.scala 687:13]
  assign isu_io_wb_rfDest = wbu_io__wb_rfDest; // @[Backend.scala 687:13]
  assign isu_io_wb_rfData = wbu_io__wb_rfData; // @[Backend.scala 687:13]
  assign isu_io_forward_valid = exu_io__forward_valid; // @[Backend.scala 690:18]
  assign isu_io_forward_wb_rfWen = exu_io__forward_wb_rfWen; // @[Backend.scala 690:18]
  assign isu_io_forward_wb_rfDest = exu_io__forward_wb_rfDest; // @[Backend.scala 690:18]
  assign isu_io_forward_wb_rfData = exu_io__forward_wb_rfData; // @[Backend.scala 690:18]
  assign isu_io_forward_fuType = exu_io__forward_fuType; // @[Backend.scala 690:18]
  assign isu_io_flush = io_flush[0]; // @[Backend.scala 684:27]
  assign isu_isu_perm_lib_ld = exu_isuPermitLibLoad;
  assign isu_isu_perm_lib_st = exu_isuPermitLibStore;
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io__in_valid = REG; // @[Pipeline.scala 31:17]
  assign exu_io__in_bits_cf_instr = REG_1_cf_instr; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pc = REG_1_cf_pc; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pnpc = REG_1_cf_pnpc; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_1 = REG_1_cf_exceptionVec_1; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_2 = REG_1_cf_exceptionVec_2; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_12 = REG_1_cf_exceptionVec_12; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_0 = REG_1_cf_intrVec_0; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_1 = REG_1_cf_intrVec_1; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_2 = REG_1_cf_intrVec_2; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_3 = REG_1_cf_intrVec_3; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_4 = REG_1_cf_intrVec_4; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_5 = REG_1_cf_intrVec_5; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_6 = REG_1_cf_intrVec_6; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_7 = REG_1_cf_intrVec_7; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_8 = REG_1_cf_intrVec_8; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_9 = REG_1_cf_intrVec_9; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_10 = REG_1_cf_intrVec_10; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_11 = REG_1_cf_intrVec_11; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_brIdx = REG_1_cf_brIdx; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_crossPageIPFFix = REG_1_cf_crossPageIPFFix; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuType = REG_1_ctrl_fuType; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuOpType = REG_1_ctrl_fuOpType; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfWen = REG_1_ctrl_rfWen; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfDest = REG_1_ctrl_rfDest; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_permitLibLoad = REG_1_ctrl_permitLibLoad; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_permitLibStore = REG_1_ctrl_permitLibStore; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_lsuIsLoad = REG_1_ctrl_lsuIsLoad; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src1 = REG_1_data_src1; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src2 = REG_1_data_src2; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_imm = REG_1_data_imm; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_addr = REG_1_data_addr; // @[Pipeline.scala 30:16]
  assign exu_io__out_ready = 1'h1; // @[Pipeline.scala 29:16]
  assign exu_io__flush = io_flush[1]; // @[Backend.scala 685:27]
  assign exu_io__dmem_req_ready = io_dmem_req_ready; // @[Backend.scala 694:11]
  assign exu_io__dmem_resp_valid = io_dmem_resp_valid; // @[Backend.scala 694:11]
  assign exu_io__dmem_resp_bits_rdata = io_dmem_resp_bits_rdata; // @[Backend.scala 694:11]
  assign exu_io__memMMU_dmem_loadPF = io_memMMU_dmem_loadPF; // @[Backend.scala 693:18]
  assign exu_io__memMMU_dmem_storePF = io_memMMU_dmem_storePF; // @[Backend.scala 693:18]
  assign exu_io__memMMU_dmem_addr = io_memMMU_dmem_addr; // @[Backend.scala 693:18]
  assign exu__T_28_0 = _T_28;
  assign exu_io_in_valid = wbu_io_in_valid;
  assign exu_io_extra_mtip = io_extra_mtip;
  assign exu_io_extra_meip_0 = io_extra_meip_0;
  assign exu_vmEnable = vmEnable;
  assign exu_isuAddr = isu_isuAddr_0;
  assign exu__T_27_0 = _T_27;
  assign exu_io_extra_msip = io_extra_msip;
  assign exu_falseWire = wbu_falseWire_0;
  assign wbu_io__in_valid = REG_2; // @[Pipeline.scala 31:17]
  assign wbu_io__in_bits_decode_cf_pc = REG_3_decode_cf_pc; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_target = REG_3_decode_cf_redirect_target; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_valid = REG_3_decode_cf_redirect_valid; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_fuType = REG_3_decode_ctrl_fuType; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfWen = REG_3_decode_ctrl_rfWen; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfDest = REG_3_decode_ctrl_rfDest; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_0 = REG_3_commits_0; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_1 = REG_3_commits_1; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_2 = REG_3_commits_2; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_3 = REG_3_commits_3; // @[Pipeline.scala 30:16]
  always @(posedge clock) begin
    if (reset) begin // @[Pipeline.scala 24:24]
      REG <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (io_flush[0]) begin // @[Pipeline.scala 27:20]
      REG <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG <= _GEN_1;
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_instr <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_instr <= isu_io_out_bits_cf_instr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_pc <= 39'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_pc <= isu_io_out_bits_cf_pc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_pnpc <= 39'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_pnpc <= isu_io_out_bits_cf_pnpc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_exceptionVec_1 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_exceptionVec_1 <= isu_io_out_bits_cf_exceptionVec_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_exceptionVec_2 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_exceptionVec_2 <= isu_io_out_bits_cf_exceptionVec_2; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_exceptionVec_12 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_exceptionVec_12 <= isu_io_out_bits_cf_exceptionVec_12; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_intrVec_0 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_intrVec_0 <= isu_io_out_bits_cf_intrVec_0; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_intrVec_1 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_intrVec_1 <= isu_io_out_bits_cf_intrVec_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_intrVec_2 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_intrVec_2 <= isu_io_out_bits_cf_intrVec_2; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_intrVec_3 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_intrVec_3 <= isu_io_out_bits_cf_intrVec_3; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_intrVec_4 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_intrVec_4 <= isu_io_out_bits_cf_intrVec_4; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_intrVec_5 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_intrVec_5 <= isu_io_out_bits_cf_intrVec_5; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_intrVec_6 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_intrVec_6 <= isu_io_out_bits_cf_intrVec_6; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_intrVec_7 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_intrVec_7 <= isu_io_out_bits_cf_intrVec_7; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_intrVec_8 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_intrVec_8 <= isu_io_out_bits_cf_intrVec_8; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_intrVec_9 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_intrVec_9 <= isu_io_out_bits_cf_intrVec_9; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_intrVec_10 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_intrVec_10 <= isu_io_out_bits_cf_intrVec_10; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_intrVec_11 <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_intrVec_11 <= isu_io_out_bits_cf_intrVec_11; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_brIdx <= 4'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_brIdx <= isu_io_out_bits_cf_brIdx; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_cf_crossPageIPFFix <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_cf_crossPageIPFFix <= isu_io_out_bits_cf_crossPageIPFFix; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_ctrl_fuType <= 3'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_ctrl_fuType <= isu_io_out_bits_ctrl_fuType; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_ctrl_fuOpType <= 7'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_ctrl_fuOpType <= isu_io_out_bits_ctrl_fuOpType; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_ctrl_rfWen <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_ctrl_rfWen <= isu_io_out_bits_ctrl_rfWen; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_ctrl_rfDest <= 5'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_ctrl_rfDest <= isu_io_out_bits_ctrl_rfDest; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_ctrl_permitLibLoad <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_ctrl_permitLibLoad <= isu_io_out_bits_ctrl_permitLibLoad; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_ctrl_permitLibStore <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_ctrl_permitLibStore <= isu_io_out_bits_ctrl_permitLibStore; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_ctrl_lsuIsLoad <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_ctrl_lsuIsLoad <= isu_io_out_bits_ctrl_lsuIsLoad; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_data_src1 <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_data_src1 <= isu_io_out_bits_data_src1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_data_src2 <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_data_src2 <= isu_io_out_bits_data_src2; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_data_imm <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_data_imm <= isu_io_out_bits_data_imm; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_data_addr <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_data_addr <= isu_io_out_bits_data_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Pipeline.scala 24:24]
      REG_2 <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (io_flush[1]) begin // @[Pipeline.scala 27:20]
      REG_2 <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG_2 <= _T_5;
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_decode_cf_pc <= 39'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_decode_cf_pc <= exu_io__out_bits_decode_cf_pc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_decode_cf_redirect_target <= 39'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_decode_cf_redirect_target <= exu_io__out_bits_decode_cf_redirect_target; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_decode_cf_redirect_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_decode_cf_redirect_valid <= exu_io__out_bits_decode_cf_redirect_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_decode_ctrl_fuType <= 3'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_decode_ctrl_fuType <= exu_io__out_bits_decode_ctrl_fuType; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_decode_ctrl_rfWen <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_decode_ctrl_rfWen <= exu_io__out_bits_decode_ctrl_rfWen; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_decode_ctrl_rfDest <= 5'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_decode_ctrl_rfDest <= exu_io__out_bits_decode_ctrl_rfDest; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_commits_0 <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_commits_0 <= exu_io__out_bits_commits_0; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_commits_1 <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_commits_1 <= exu_io__out_bits_commits_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_commits_2 <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_commits_2 <= exu_io__out_bits_commits_2; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_commits_3 <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_commits_3 <= exu_io__out_bits_commits_3; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  REG_1_cf_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  REG_1_cf_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  REG_1_cf_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  REG_1_cf_exceptionVec_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1_cf_exceptionVec_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  REG_1_cf_exceptionVec_12 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  REG_1_cf_intrVec_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  REG_1_cf_intrVec_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  REG_1_cf_intrVec_2 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  REG_1_cf_intrVec_3 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG_1_cf_intrVec_4 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  REG_1_cf_intrVec_5 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  REG_1_cf_intrVec_6 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  REG_1_cf_intrVec_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  REG_1_cf_intrVec_8 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  REG_1_cf_intrVec_9 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  REG_1_cf_intrVec_10 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  REG_1_cf_intrVec_11 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  REG_1_cf_brIdx = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  REG_1_cf_crossPageIPFFix = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  REG_1_ctrl_fuType = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  REG_1_ctrl_fuOpType = _RAND_22[6:0];
  _RAND_23 = {1{`RANDOM}};
  REG_1_ctrl_rfWen = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  REG_1_ctrl_rfDest = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  REG_1_ctrl_permitLibLoad = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  REG_1_ctrl_permitLibStore = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  REG_1_ctrl_lsuIsLoad = _RAND_27[0:0];
  _RAND_28 = {2{`RANDOM}};
  REG_1_data_src1 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  REG_1_data_src2 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  REG_1_data_imm = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  REG_1_data_addr = _RAND_31[63:0];
  _RAND_32 = {1{`RANDOM}};
  REG_2 = _RAND_32[0:0];
  _RAND_33 = {2{`RANDOM}};
  REG_3_decode_cf_pc = _RAND_33[38:0];
  _RAND_34 = {2{`RANDOM}};
  REG_3_decode_cf_redirect_target = _RAND_34[38:0];
  _RAND_35 = {1{`RANDOM}};
  REG_3_decode_cf_redirect_valid = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  REG_3_decode_ctrl_fuType = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  REG_3_decode_ctrl_rfWen = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  REG_3_decode_ctrl_rfDest = _RAND_38[4:0];
  _RAND_39 = {2{`RANDOM}};
  REG_3_commits_0 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  REG_3_commits_1 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  REG_3_commits_2 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  REG_3_commits_3 = _RAND_42[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_LockingArbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [2:0]  io_in_0_bits_size,
  input  [3:0]  io_in_0_bits_cmd,
  input  [7:0]  io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [2:0]  io_in_1_bits_size,
  input  [3:0]  io_in_1_bits_cmd,
  input  [7:0]  io_in_1_bits_wmask,
  input  [63:0] io_in_1_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata,
  output        io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] value; // @[Counter.scala 60:40]
  reg  REG; // @[Arbiter.scala 46:22]
  wire  _T = value != 3'h0; // @[Arbiter.scala 47:34]
  wire  _T_3 = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[Crossbar.scala 100:62]
  wire  _T_4 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _value_T_1 = value + 3'h1; // @[Counter.scala 76:24]
  wire  choice = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 88:27 Arbiter.scala 88:36]
  wire  _T_7 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_9 = _T ? ~REG : 1'h1; // @[Arbiter.scala 57:22]
  wire  _T_12 = _T ? REG : _T_7; // @[Arbiter.scala 57:22]
  assign io_in_0_ready = _T_9 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_in_1_ready = _T_12 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16 Arbiter.scala 41:16]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_size = io_chosen ? io_in_1_bits_size : io_in_0_bits_size; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_cmd = io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_wmask = io_chosen ? io_in_1_bits_wmask : io_in_0_bits_wmask; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_wdata = io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_chosen = _T ? REG : choice; // @[Arbiter.scala 55:19 Arbiter.scala 55:31 Arbiter.scala 40:13]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 60:40]
      value <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_4 & _T_3) begin // @[Arbiter.scala 50:39]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (_T_4 & _T_3) begin // @[Arbiter.scala 50:39]
      REG <= io_chosen; // @[Arbiter.scala 51:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  REG = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_SimpleBusCrossbarNto1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [31:0] io_in_0_req_bits_addr,
  input  [2:0]  io_in_0_req_bits_size,
  input  [3:0]  io_in_0_req_bits_cmd,
  input  [7:0]  io_in_0_req_bits_wmask,
  input  [63:0] io_in_0_req_bits_wdata,
  input         io_in_0_resp_ready,
  output        io_in_0_resp_valid,
  output [3:0]  io_in_0_resp_bits_cmd,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [31:0] io_in_1_req_bits_addr,
  input  [2:0]  io_in_1_req_bits_size,
  input  [3:0]  io_in_1_req_bits_cmd,
  input  [7:0]  io_in_1_req_bits_wmask,
  input  [63:0] io_in_1_req_bits_wdata,
  input         io_in_1_resp_ready,
  output        io_in_1_resp_valid,
  output [3:0]  io_in_1_resp_bits_cmd,
  output [63:0] io_in_1_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[Crossbar.scala 101:24]
  wire  inputArb_reset; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_in_0_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_in_1_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_1_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_out_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_chosen; // @[Crossbar.scala 101:24]
  reg [1:0] state; // @[Crossbar.scala 98:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  reg  inflightSrc; // @[Crossbar.scala 105:28]
  wire  _T_14 = state == 2'h0; // @[Crossbar.scala 109:47]
  wire  _T_18 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_19 = inputArb_io_out_ready & inputArb_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_25 = inputArb_io_out_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_26 = inputArb_io_out_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire [1:0] _GEN_4 = _T_25 | _T_26 ? 2'h2 : state; // @[Crossbar.scala 124:80 Crossbar.scala 124:88 Crossbar.scala 98:22]
  wire  _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_29 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_30 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_32 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_9 = _T_29 ? 2'h0 : state; // @[Crossbar.scala 128:50 Crossbar.scala 128:58 Crossbar.scala 98:22]
  ysyx_210000_LockingArbiter inputArb ( // @[Crossbar.scala 101:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_size(inputArb_io_in_0_bits_size),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_size(inputArb_io_in_1_bits_size),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(inputArb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[Crossbar.scala 102:68]
  assign io_in_0_resp_valid = ~inflightSrc & io_out_resp_valid; // @[Crossbar.scala 115:13 Crossbar.scala 115:13 Crossbar.scala 113:26]
  assign io_in_0_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[Crossbar.scala 102:68]
  assign io_in_1_resp_valid = inflightSrc & io_out_resp_valid; // @[Crossbar.scala 115:13 Crossbar.scala 115:13 Crossbar.scala 113:26]
  assign io_in_1_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[Crossbar.scala 109:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[Crossbar.scala 107:19]
  assign io_out_resp_ready = inflightSrc ? io_in_1_resp_ready : io_in_0_resp_ready; // @[Crossbar.scala 116:13 Crossbar.scala 116:13]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_size = io_in_0_req_bits_size; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_size = io_in_1_req_bits_size; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_wmask = io_in_1_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_out_ready = io_out_req_ready & _T_14; // @[Crossbar.scala 110:37]
  always @(posedge clock) begin
    if (reset) begin // @[Crossbar.scala 98:22]
      state <= 2'h0; // @[Crossbar.scala 98:22]
    end else if (_T_18) begin // @[Conditional.scala 40:58]
      if (_T_19) begin // @[Crossbar.scala 121:29]
        if (_T_4) begin // @[Crossbar.scala 123:38]
          state <= 2'h1; // @[Crossbar.scala 123:46]
        end else begin
          state <= _GEN_4;
        end
      end
    end else if (_T_28) begin // @[Conditional.scala 39:67]
      if (_T_29 & _T_30) begin // @[Crossbar.scala 127:82]
        state <= 2'h0; // @[Crossbar.scala 127:90]
      end
    end else if (_T_32) begin // @[Conditional.scala 39:67]
      state <= _GEN_9;
    end
    if (reset) begin // @[Crossbar.scala 105:28]
      inflightSrc <= 1'h0; // @[Crossbar.scala 105:28]
    end else if (_T_18) begin // @[Conditional.scala 40:58]
      if (_T_19) begin // @[Crossbar.scala 121:29]
        inflightSrc <= inputArb_io_chosen; // @[Crossbar.scala 122:21]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(inputArb_io_out_valid & ~_T_4 & _T_1) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:104 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[Crossbar.scala 104:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(inputArb_io_out_valid & ~_T_4 & _T_1) | reset)) begin
          $fatal; // @[Crossbar.scala 104:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_LockingArbiter_1(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [2:0]  io_in_0_bits_size,
  input  [3:0]  io_in_0_bits_cmd,
  input  [7:0]  io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [3:0]  io_in_1_bits_cmd,
  input  [63:0] io_in_1_bits_wdata,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_addr,
  input  [3:0]  io_in_2_bits_cmd,
  input  [63:0] io_in_2_bits_wdata,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_addr,
  input  [2:0]  io_in_3_bits_size,
  input  [3:0]  io_in_3_bits_cmd,
  input  [7:0]  io_in_3_bits_wmask,
  input  [63:0] io_in_3_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata,
  output [1:0]  io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_1 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16 Arbiter.scala 41:16]
  wire  _GEN_2 = 2'h2 == io_chosen ? io_in_2_valid : _GEN_1; // @[Arbiter.scala 41:16 Arbiter.scala 41:16]
  wire [63:0] _GEN_5 = 2'h1 == io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [63:0] _GEN_6 = 2'h2 == io_chosen ? io_in_2_bits_wdata : _GEN_5; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [7:0] _GEN_9 = 2'h1 == io_chosen ? 8'hff : io_in_0_bits_wmask; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [7:0] _GEN_10 = 2'h2 == io_chosen ? 8'hff : _GEN_9; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [3:0] _GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [3:0] _GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_cmd : _GEN_13; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [2:0] _GEN_17 = 2'h1 == io_chosen ? 3'h3 : io_in_0_bits_size; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [2:0] _GEN_18 = 2'h2 == io_chosen ? 3'h3 : _GEN_17; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [31:0] _GEN_21 = 2'h1 == io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  wire [31:0] _GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_addr : _GEN_21; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  reg [2:0] value; // @[Counter.scala 60:40]
  reg [1:0] REG; // @[Arbiter.scala 46:22]
  wire  _T = value != 3'h0; // @[Arbiter.scala 47:34]
  wire  _T_3 = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[Crossbar.scala 100:62]
  wire  _T_4 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _value_T_1 = value + 3'h1; // @[Counter.scala 76:24]
  wire [1:0] _GEN_27 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 88:27 Arbiter.scala 88:36]
  wire [1:0] _GEN_28 = io_in_1_valid ? 2'h1 : _GEN_27; // @[Arbiter.scala 88:27 Arbiter.scala 88:36]
  wire [1:0] choice = io_in_0_valid ? 2'h0 : _GEN_28; // @[Arbiter.scala 88:27 Arbiter.scala 88:36]
  wire  _T_9 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_10 = ~(io_in_0_valid | io_in_1_valid); // @[Arbiter.scala 31:78]
  wire  _T_11 = ~(io_in_0_valid | io_in_1_valid | io_in_2_valid); // @[Arbiter.scala 31:78]
  wire  _T_13 = _T ? REG == 2'h0 : 1'h1; // @[Arbiter.scala 57:22]
  wire  _T_16 = _T ? REG == 2'h1 : _T_9; // @[Arbiter.scala 57:22]
  wire  _T_19 = _T ? REG == 2'h2 : _T_10; // @[Arbiter.scala 57:22]
  wire  _T_22 = _T ? REG == 2'h3 : _T_11; // @[Arbiter.scala 57:22]
  assign io_in_0_ready = _T_13 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_in_1_ready = _T_16 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_in_2_ready = _T_19 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_in_3_ready = _T_22 & io_out_ready; // @[Arbiter.scala 57:56]
  assign io_out_valid = 2'h3 == io_chosen ? io_in_3_valid : _GEN_2; // @[Arbiter.scala 41:16 Arbiter.scala 41:16]
  assign io_out_bits_addr = 2'h3 == io_chosen ? io_in_3_bits_addr : _GEN_22; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_size = 2'h3 == io_chosen ? io_in_3_bits_size : _GEN_18; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_cmd = 2'h3 == io_chosen ? io_in_3_bits_cmd : _GEN_14; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_wmask = 2'h3 == io_chosen ? io_in_3_bits_wmask : _GEN_10; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_out_bits_wdata = 2'h3 == io_chosen ? io_in_3_bits_wdata : _GEN_6; // @[Arbiter.scala 42:15 Arbiter.scala 42:15]
  assign io_chosen = _T ? REG : choice; // @[Arbiter.scala 55:19 Arbiter.scala 55:31 Arbiter.scala 40:13]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 60:40]
      value <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_4 & _T_3) begin // @[Arbiter.scala 50:39]
      value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (_T_4 & _T_3) begin // @[Arbiter.scala 50:39]
      REG <= io_chosen; // @[Arbiter.scala 51:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  REG = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_SimpleBusCrossbarNto1_1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [31:0] io_in_0_req_bits_addr,
  input  [2:0]  io_in_0_req_bits_size,
  input  [3:0]  io_in_0_req_bits_cmd,
  input  [7:0]  io_in_0_req_bits_wmask,
  input  [63:0] io_in_0_req_bits_wdata,
  output        io_in_0_resp_valid,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [31:0] io_in_1_req_bits_addr,
  input  [3:0]  io_in_1_req_bits_cmd,
  input  [63:0] io_in_1_req_bits_wdata,
  output        io_in_1_resp_valid,
  output [63:0] io_in_1_resp_bits_rdata,
  output        io_in_2_req_ready,
  input         io_in_2_req_valid,
  input  [31:0] io_in_2_req_bits_addr,
  input  [3:0]  io_in_2_req_bits_cmd,
  input  [63:0] io_in_2_req_bits_wdata,
  output        io_in_2_resp_valid,
  output [63:0] io_in_2_resp_bits_rdata,
  output        io_in_3_req_ready,
  input         io_in_3_req_valid,
  input  [31:0] io_in_3_req_bits_addr,
  input  [2:0]  io_in_3_req_bits_size,
  input  [3:0]  io_in_3_req_bits_cmd,
  input  [7:0]  io_in_3_req_bits_wmask,
  input  [63:0] io_in_3_req_bits_wdata,
  input         io_in_3_resp_ready,
  output        io_in_3_resp_valid,
  output [3:0]  io_in_3_resp_bits_cmd,
  output [63:0] io_in_3_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[Crossbar.scala 101:24]
  wire  inputArb_reset; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_in_0_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_2_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_2_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_2_bits_addr; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_2_bits_cmd; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_2_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_3_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_3_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_3_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_in_3_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_3_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_3_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_3_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_out_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[Crossbar.scala 101:24]
  wire [1:0] inputArb_io_chosen; // @[Crossbar.scala 101:24]
  reg [1:0] state; // @[Crossbar.scala 98:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_4 = ~inputArb_io_out_bits_cmd[0] & ~inputArb_io_out_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  reg [1:0] inflightSrc; // @[Crossbar.scala 105:28]
  wire  _T_14 = state == 2'h0; // @[Crossbar.scala 109:47]
  wire  _T_18 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_19 = inputArb_io_out_ready & inputArb_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_25 = inputArb_io_out_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_26 = inputArb_io_out_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire [1:0] _GEN_8 = _T_25 | _T_26 ? 2'h2 : state; // @[Crossbar.scala 124:80 Crossbar.scala 124:88 Crossbar.scala 98:22]
  wire  _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_29 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_30 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_32 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_13 = _T_29 ? 2'h0 : state; // @[Crossbar.scala 128:50 Crossbar.scala 128:58 Crossbar.scala 98:22]
  ysyx_210000_LockingArbiter_1 inputArb ( // @[Crossbar.scala 101:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_size(inputArb_io_in_0_bits_size),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_in_2_ready(inputArb_io_in_2_ready),
    .io_in_2_valid(inputArb_io_in_2_valid),
    .io_in_2_bits_addr(inputArb_io_in_2_bits_addr),
    .io_in_2_bits_cmd(inputArb_io_in_2_bits_cmd),
    .io_in_2_bits_wdata(inputArb_io_in_2_bits_wdata),
    .io_in_3_ready(inputArb_io_in_3_ready),
    .io_in_3_valid(inputArb_io_in_3_valid),
    .io_in_3_bits_addr(inputArb_io_in_3_bits_addr),
    .io_in_3_bits_size(inputArb_io_in_3_bits_size),
    .io_in_3_bits_cmd(inputArb_io_in_3_bits_cmd),
    .io_in_3_bits_wmask(inputArb_io_in_3_bits_wmask),
    .io_in_3_bits_wdata(inputArb_io_in_3_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[Crossbar.scala 102:68]
  assign io_in_0_resp_valid = 2'h0 == inflightSrc & io_out_resp_valid; // @[Crossbar.scala 115:13 Crossbar.scala 115:13 Crossbar.scala 113:26]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[Crossbar.scala 102:68]
  assign io_in_1_resp_valid = 2'h1 == inflightSrc & io_out_resp_valid; // @[Crossbar.scala 115:13 Crossbar.scala 115:13 Crossbar.scala 113:26]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_2_req_ready = inputArb_io_in_2_ready; // @[Crossbar.scala 102:68]
  assign io_in_2_resp_valid = 2'h2 == inflightSrc & io_out_resp_valid; // @[Crossbar.scala 115:13 Crossbar.scala 115:13 Crossbar.scala 113:26]
  assign io_in_2_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_3_req_ready = inputArb_io_in_3_ready; // @[Crossbar.scala 102:68]
  assign io_in_3_resp_valid = 2'h3 == inflightSrc & io_out_resp_valid; // @[Crossbar.scala 115:13 Crossbar.scala 115:13 Crossbar.scala 113:26]
  assign io_in_3_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_3_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_out_req_valid = inputArb_io_out_valid & state == 2'h0; // @[Crossbar.scala 109:37]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[Crossbar.scala 107:19]
  assign io_out_resp_ready = 2'h3 == inflightSrc ? io_in_3_resp_ready : 1'h1; // @[Crossbar.scala 116:13 Crossbar.scala 116:13]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_size = io_in_0_req_bits_size; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_valid = io_in_2_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_bits_addr = io_in_2_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_bits_cmd = io_in_2_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_bits_wdata = io_in_2_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_valid = io_in_3_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_addr = io_in_3_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_size = io_in_3_req_bits_size; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_cmd = io_in_3_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_wmask = io_in_3_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_wdata = io_in_3_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_out_ready = io_out_req_ready & _T_14; // @[Crossbar.scala 110:37]
  always @(posedge clock) begin
    if (reset) begin // @[Crossbar.scala 98:22]
      state <= 2'h0; // @[Crossbar.scala 98:22]
    end else if (_T_18) begin // @[Conditional.scala 40:58]
      if (_T_19) begin // @[Crossbar.scala 121:29]
        if (_T_4) begin // @[Crossbar.scala 123:38]
          state <= 2'h1; // @[Crossbar.scala 123:46]
        end else begin
          state <= _GEN_8;
        end
      end
    end else if (_T_28) begin // @[Conditional.scala 39:67]
      if (_T_29 & _T_30) begin // @[Crossbar.scala 127:82]
        state <= 2'h0; // @[Crossbar.scala 127:90]
      end
    end else if (_T_32) begin // @[Conditional.scala 39:67]
      state <= _GEN_13;
    end
    if (reset) begin // @[Crossbar.scala 105:28]
      inflightSrc <= 2'h0; // @[Crossbar.scala 105:28]
    end else if (_T_18) begin // @[Conditional.scala 40:58]
      if (_T_19) begin // @[Crossbar.scala 121:29]
        inflightSrc <= inputArb_io_chosen; // @[Crossbar.scala 122:21]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(inputArb_io_out_valid & ~_T_4 & _T_1) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Crossbar.scala:104 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[Crossbar.scala 104:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(inputArb_io_out_valid & ~_T_4 & _T_1) | reset)) begin
          $fatal; // @[Crossbar.scala 104:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_MMIOBridge(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] state; // @[NutCore.scala 125:22]
  wire  _T = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg [31:0] in_reqLatch_addr; // @[Reg.scala 27:20]
  wire  _T_1 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = _T_1 & state == 8'h2; // @[NutCore.scala 127:72]
  reg [63:0] REG_rdata; // @[Reg.scala 27:20]
  wire [63:0] _GEN_5 = _T_3 ? io_out_resp_bits_rdata : REG_rdata; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _T_6 = _T_1 & state == 8'h4; // @[NutCore.scala 128:72]
  reg [63:0] REG_1_rdata; // @[Reg.scala 27:20]
  wire [63:0] _GEN_7 = _T_6 ? io_out_resp_bits_rdata : REG_1_rdata; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  reg  normal; // @[NutCore.scala 129:23]
  wire  _T_9 = io_in_req_bits_size == 3'h3; // @[NutCore.scala 132:38]
  wire  in_sel = ~(io_in_req_bits_size == 3'h3); // @[NutCore.scala 132:16]
  wire  _T_10 = 8'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_16 = 8'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_17 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_18 = 8'h2 == state; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_16 = _T_1 ? 8'h3 : state; // @[NutCore.scala 153:33 NutCore.scala 155:15 NutCore.scala 125:22]
  wire  _T_20 = 8'h3 == state; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_17 = _T_17 ? 8'h4 : state; // @[NutCore.scala 159:32 NutCore.scala 160:15 NutCore.scala 125:22]
  wire  _T_22 = 8'h4 == state; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_18 = _T_1 ? 8'h5 : state; // @[NutCore.scala 164:33 NutCore.scala 165:15 NutCore.scala 125:22]
  wire  _T_24 = 8'h5 == state; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_19 = io_in_resp_valid ? 8'h0 : state; // @[NutCore.scala 169:32 NutCore.scala 170:15 NutCore.scala 125:22]
  wire  _T_26 = 8'h6 == state; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_20 = _T_17 ? 8'h7 : state; // @[NutCore.scala 176:32 NutCore.scala 177:15 NutCore.scala 125:22]
  wire  _T_28 = 8'h7 == state; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_22 = _T_28 ? _GEN_18 : state; // @[Conditional.scala 39:67 NutCore.scala 125:22]
  wire [7:0] _GEN_23 = _T_26 ? _GEN_20 : _GEN_22; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_24 = _T_24 ? _GEN_19 : _GEN_23; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_25 = _T_22 ? _GEN_18 : _GEN_24; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_26 = _T_20 ? _GEN_17 : _GEN_25; // @[Conditional.scala 39:67]
  wire  _T_30 = state == 8'h0; // @[NutCore.scala 187:58]
  wire [31:0] hi = _GEN_7[31:0]; // @[NutCore.scala 190:88]
  wire [31:0] lo = _GEN_5[31:0]; // @[NutCore.scala 190:116]
  wire [63:0] _T_35 = {hi,lo}; // @[Cat.scala 30:58]
  wire  _T_37 = state == 8'h1; // @[NutCore.scala 192:30]
  wire [28:0] hi_1 = in_reqLatch_addr[31:3]; // @[NutCore.scala 194:103]
  wire [31:0] _T_45 = {hi_1,3'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_48 = _T_45 + 32'h4; // @[NutCore.scala 194:158]
  wire [31:0] _T_49 = _T_37 ? _T_45 : _T_48; // @[NutCore.scala 194:64]
  assign io_in_req_ready = in_sel ? io_out_req_ready : state == 8'h0; // @[NutCore.scala 187:25]
  assign io_in_resp_valid = normal ? io_out_resp_valid : state == 8'h5; // @[NutCore.scala 188:26]
  assign io_in_resp_bits_rdata = normal ? io_out_resp_bits_rdata : _T_35; // @[NutCore.scala 190:31]
  assign io_out_req_valid = state == 8'h1 | state == 8'h3 | _T_30 & io_in_req_valid & in_sel; // @[NutCore.scala 192:64]
  assign io_out_req_bits_addr = in_sel ? io_in_req_bits_addr : _T_49; // @[NutCore.scala 194:31]
  assign io_out_req_bits_size = in_sel ? io_in_req_bits_size : 3'h2; // @[NutCore.scala 195:30]
  assign io_out_resp_ready = 1'h1; // @[NutCore.scala 199:27]
  always @(posedge clock) begin
    if (reset) begin // @[NutCore.scala 125:22]
      state <= 8'h0; // @[NutCore.scala 125:22]
    end else if (_T_10) begin // @[Conditional.scala 40:58]
      if (_T) begin // @[NutCore.scala 136:31]
        if (_T_9) begin // @[NutCore.scala 137:48]
          state <= 8'h1; // @[NutCore.scala 138:17]
        end
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      if (_T_17) begin // @[NutCore.scala 147:32]
        state <= 8'h2; // @[NutCore.scala 149:15]
      end
    end else if (_T_18) begin // @[Conditional.scala 39:67]
      state <= _GEN_16;
    end else begin
      state <= _GEN_26;
    end
    if (reset) begin // @[Reg.scala 27:20]
      in_reqLatch_addr <= 32'h0; // @[Reg.scala 27:20]
    end else if (_T) begin // @[Reg.scala 28:19]
      in_reqLatch_addr <= io_in_req_bits_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_rdata <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_3) begin // @[Reg.scala 28:19]
      REG_rdata <= io_out_resp_bits_rdata; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_rdata <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_6) begin // @[Reg.scala 28:19]
      REG_1_rdata <= io_out_resp_bits_rdata; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[NutCore.scala 129:23]
      normal <= 1'h0; // @[NutCore.scala 129:23]
    end else if (_T_10) begin // @[Conditional.scala 40:58]
      if (_T) begin // @[NutCore.scala 136:31]
        if (_T_9) begin // @[NutCore.scala 137:48]
          normal <= 1'h0; // @[NutCore.scala 139:18]
        end else begin
          normal <= 1'h1; // @[NutCore.scala 142:18]
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & _T & in_sel & ~reset) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NutCore.scala:141 assert(false.B)\n"); // @[NutCore.scala 141:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10 & _T & in_sel & ~reset) begin
          $fatal; // @[NutCore.scala 141:17]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  in_reqLatch_addr = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  REG_rdata = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  REG_1_rdata = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  normal = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_EmbeddedTLBExec(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [38:0]  io_in_bits_addr,
  input  [2:0]   io_in_bits_size,
  input  [86:0]  io_in_bits_user,
  input          io_out_ready,
  output         io_out_valid,
  output [31:0]  io_out_bits_addr,
  output [2:0]   io_out_bits_size,
  output [86:0]  io_out_bits_user,
  input  [120:0] io_md_0,
  input  [120:0] io_md_1,
  input  [120:0] io_md_2,
  input  [120:0] io_md_3,
  output         io_mdWrite_wen,
  output [3:0]   io_mdWrite_waymask,
  output [120:0] io_mdWrite_wdata,
  input          io_mdReady,
  input          io_mem_req_ready,
  output         io_mem_req_valid,
  output [31:0]  io_mem_req_bits_addr,
  output [3:0]   io_mem_req_bits_cmd,
  output [63:0]  io_mem_req_bits_wdata,
  output         io_mem_resp_ready,
  input          io_mem_resp_valid,
  input  [63:0]  io_mem_resp_bits_rdata,
  input          io_flush,
  input  [63:0]  io_satp,
  input  [1:0]   io_pf_priviledgeMode,
  output         io_pf_loadPF,
  output         io_pf_storePF,
  output         io_ipf,
  output         io_isFinish
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[EmbeddedTLB.scala 193:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[EmbeddedTLB.scala 193:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[EmbeddedTLB.scala 193:54]
  wire [19:0] satp_ppn = io_satp[19:0]; // @[EmbeddedTLB.scala 195:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[EmbeddedTLB.scala 195:30]
  wire [26:0] _T_43 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[EmbeddedTLB.scala 204:201]
  wire [26:0] _T_44 = {9'h1ff,io_md_0[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_45 = _T_44 & io_md_0[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_47 = _T_44 & _T_43; // @[TLB.scala 131:84]
  wire  _T_48 = _T_45 == _T_47; // @[TLB.scala 131:48]
  wire  _T_49 = io_md_0[52] & io_md_0[93:78] == satp_asid & _T_48; // @[EmbeddedTLB.scala 204:132]
  wire [26:0] _T_85 = {9'h1ff,io_md_1[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_86 = _T_85 & io_md_1[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_88 = _T_85 & _T_43; // @[TLB.scala 131:84]
  wire  _T_89 = _T_86 == _T_88; // @[TLB.scala 131:48]
  wire  _T_90 = io_md_1[52] & io_md_1[93:78] == satp_asid & _T_89; // @[EmbeddedTLB.scala 204:132]
  wire [26:0] _T_126 = {9'h1ff,io_md_2[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_127 = _T_126 & io_md_2[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_129 = _T_126 & _T_43; // @[TLB.scala 131:84]
  wire  _T_130 = _T_127 == _T_129; // @[TLB.scala 131:48]
  wire  _T_131 = io_md_2[52] & io_md_2[93:78] == satp_asid & _T_130; // @[EmbeddedTLB.scala 204:132]
  wire [26:0] _T_167 = {9'h1ff,io_md_3[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_168 = _T_167 & io_md_3[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_170 = _T_167 & _T_43; // @[TLB.scala 131:84]
  wire  _T_171 = _T_168 == _T_170; // @[TLB.scala 131:48]
  wire  _T_172 = io_md_3[52] & io_md_3[93:78] == satp_asid & _T_171; // @[EmbeddedTLB.scala 204:132]
  wire [3:0] hitVec = {_T_172,_T_131,_T_90,_T_49}; // @[EmbeddedTLB.scala 204:211]
  wire  _T_173 = |hitVec; // @[EmbeddedTLB.scala 205:35]
  wire  hit = io_in_valid & |hitVec; // @[EmbeddedTLB.scala 205:25]
  wire  miss = io_in_valid & ~_T_173; // @[EmbeddedTLB.scala 206:26]
  reg [63:0] REG; // @[LFSR64.scala 25:23]
  wire  hi_5 = REG[0] ^ REG[1] ^ REG[3] ^ REG[4]; // @[LFSR64.scala 26:43]
  wire [62:0] lo_1 = REG[63:1]; // @[LFSR64.scala 28:51]
  wire [63:0] _T_183 = {hi_5,lo_1}; // @[Cat.scala 30:58]
  wire [3:0] victimWaymask = 4'h1 << REG[1:0]; // @[EmbeddedTLB.scala 208:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[EmbeddedTLB.scala 209:20]
  wire [120:0] _T_190 = waymask[0] ? io_md_0 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_191 = waymask[1] ? io_md_1 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_192 = waymask[2] ? io_md_2 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_193 = waymask[3] ? io_md_3 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_194 = _T_190 | _T_191; // @[Mux.scala 27:72]
  wire [120:0] _T_195 = _T_194 | _T_192; // @[Mux.scala 27:72]
  wire [120:0] _T_196 = _T_195 | _T_193; // @[Mux.scala 27:72]
  wire [7:0] hitMeta_flag = _T_196[59:52]; // @[EmbeddedTLB.scala 215:70]
  wire [17:0] hitMeta_mask = _T_196[77:60]; // @[EmbeddedTLB.scala 215:70]
  wire [15:0] hitMeta_asid = _T_196[93:78]; // @[EmbeddedTLB.scala 215:70]
  wire [31:0] hitData_pteaddr = _T_196[31:0]; // @[EmbeddedTLB.scala 216:70]
  wire [19:0] hitData_ppn = _T_196[51:32]; // @[EmbeddedTLB.scala 216:70]
  wire  hitFlag_v = hitMeta_flag[0]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_r = hitMeta_flag[1]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_g = hitMeta_flag[5]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[EmbeddedTLB.scala 217:38]
  wire  _T_241 = io_pf_priviledgeMode == 2'h0; // @[EmbeddedTLB.scala 226:62]
  wire  _T_246 = io_pf_priviledgeMode == 2'h1; // @[EmbeddedTLB.scala 226:110]
  wire  hitCheck = hit & ~(io_pf_priviledgeMode == 2'h0 & ~hitFlag_u) & ~(io_pf_priviledgeMode == 2'h1 & hitFlag_u); // @[EmbeddedTLB.scala 226:87]
  wire  hitExec = hitCheck & hitFlag_x; // @[EmbeddedTLB.scala 227:26]
  wire  hitinstrPF = ~hitExec & hit; // @[EmbeddedTLB.scala 239:52]
  wire  _T_235 = io_pf_loadPF | io_pf_storePF; // @[Bundle.scala 133:23]
  wire  _T_237 = ~_T_235; // @[EmbeddedTLB.scala 221:84]
  wire  hitWB = hit & ~hitFlag_a & ~hitinstrPF & ~_T_235; // @[EmbeddedTLB.scala 221:81]
  wire [7:0] _T_239 = {hitFlag_d,hitFlag_a,hitFlag_g,hitFlag_u,hitFlag_x,hitFlag_w,hitFlag_r,hitFlag_v}; // @[EmbeddedTLB.scala 222:79]
  wire [7:0] hitRefillFlag = 8'h40 | _T_239; // @[EmbeddedTLB.scala 222:69]
  wire [39:0] _T_240 = {10'h0,hitData_ppn,2'h0,hitRefillFlag}; // @[Cat.scala 30:58]
  reg [39:0] hitWBStore; // @[Reg.scala 27:20]
  reg [2:0] state; // @[EmbeddedTLB.scala 247:22]
  reg [1:0] level; // @[EmbeddedTLB.scala 248:22]
  reg [63:0] memRespStore; // @[EmbeddedTLB.scala 250:29]
  reg [17:0] missMaskStore; // @[EmbeddedTLB.scala 252:30]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[EmbeddedTLB.scala 255:49]
  wire [19:0] memRdata_ppn = io_mem_resp_bits_rdata[29:10]; // @[EmbeddedTLB.scala 255:49]
  reg [31:0] raddr; // @[EmbeddedTLB.scala 256:22]
  wire  _T_267 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_2 = _T_267 | alreadyOutFire; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  reg  needFlush; // @[EmbeddedTLB.scala 260:26]
  wire  isFlush = needFlush | io_flush; // @[EmbeddedTLB.scala 262:27]
  wire  _GEN_3 = io_flush & state != 3'h0 | needFlush; // @[EmbeddedTLB.scala 263:40 EmbeddedTLB.scala 263:52 EmbeddedTLB.scala 260:26]
  wire  _GEN_4 = _T_267 & needFlush ? 1'h0 : _GEN_3; // @[EmbeddedTLB.scala 264:37 EmbeddedTLB.scala 264:49]
  reg  missIPF; // @[EmbeddedTLB.scala 266:24]
  wire  _T_272 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_273 = ~io_flush; // @[EmbeddedTLB.scala 271:13]
  wire [31:0] _T_277 = {satp_ppn,vpn_vpn2,3'h0}; // @[Cat.scala 30:58]
  wire  _T_278 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_279 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_15 = _T_279 ? 3'h2 : state; // @[EmbeddedTLB.scala 288:38 EmbeddedTLB.scala 288:46 EmbeddedTLB.scala 247:22]
  wire  _GEN_17 = isFlush ? 1'h0 : _GEN_4; // @[EmbeddedTLB.scala 285:22 EmbeddedTLB.scala 287:19]
  wire  _T_280 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [7:0] _T_281 = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,memRdata_flag_w,
    memRdata_flag_r,memRdata_flag_v}; // @[EmbeddedTLB.scala 292:44]
  wire  _T_290 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_293 = level == 2'h3; // @[EmbeddedTLB.scala 297:58]
  wire  _T_294 = level == 2'h2; // @[EmbeddedTLB.scala 297:73]
  wire [8:0] lo_5 = _T_293 ? vpn_vpn1 : vpn_vpn0; // @[EmbeddedTLB.scala 311:50]
  wire [31:0] _T_314 = {memRdata_ppn,lo_5,3'h0}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_18 = ~_T_281[0] | ~_T_281[1] & _T_281[2] ? 3'h4 : 3'h1; // @[EmbeddedTLB.scala 298:60 EmbeddedTLB.scala 299:43 EmbeddedTLB.scala 310:19]
  wire  _GEN_19 = ~_T_281[0] | ~_T_281[1] & _T_281[2] | missIPF; // @[EmbeddedTLB.scala 298:60 EmbeddedTLB.scala 300:45 EmbeddedTLB.scala 266:24]
  wire [31:0] _GEN_20 = ~_T_281[0] | ~_T_281[1] & _T_281[2] ? raddr : _T_314; // @[EmbeddedTLB.scala 298:60 EmbeddedTLB.scala 256:22 EmbeddedTLB.scala 311:19]
  wire  _T_327 = _T_281[0] & ~(_T_241 & ~_T_281[4]) & ~(_T_246 & _T_281[4]); // @[EmbeddedTLB.scala 314:87]
  wire  _T_328 = _T_327 & _T_281[3]; // @[EmbeddedTLB.scala 315:36]
  wire  _T_333 = ~_T_281[6]; // @[EmbeddedTLB.scala 318:60]
  wire [7:0] _T_340 = {_T_281[7],_T_281[6],_T_281[5],_T_281[4],_T_281[3],_T_281[2],_T_281[1],_T_281[0]}; // @[EmbeddedTLB.scala 320:79]
  wire [7:0] _T_341 = 8'h40 | _T_340; // @[EmbeddedTLB.scala 320:68]
  wire [63:0] _T_342 = io_mem_resp_bits_rdata | 64'h40; // @[EmbeddedTLB.scala 321:50]
  wire [2:0] _T_344 = _T_333 ? 3'h3 : 3'h4; // @[EmbeddedTLB.scala 325:27]
  wire  _GEN_21 = ~_T_328 | missIPF; // @[EmbeddedTLB.scala 323:30 EmbeddedTLB.scala 323:40 EmbeddedTLB.scala 266:24]
  wire [2:0] _GEN_22 = ~_T_328 ? 3'h4 : _T_344; // @[EmbeddedTLB.scala 323:30 EmbeddedTLB.scala 323:58 EmbeddedTLB.scala 325:21]
  wire  _GEN_23 = ~_T_328 ? 1'h0 : 1'h1; // @[EmbeddedTLB.scala 323:30 EmbeddedTLB.scala 326:30]
  wire [17:0] _T_347 = _T_294 ? 18'h3fe00 : 18'h3ffff; // @[EmbeddedTLB.scala 339:59]
  wire [17:0] _T_348 = _T_293 ? 18'h0 : _T_347; // @[EmbeddedTLB.scala 339:26]
  wire [7:0] _GEN_24 = level != 2'h0 ? _T_341 : 8'h0; // @[EmbeddedTLB.scala 313:36 EmbeddedTLB.scala 320:26]
  wire [63:0] _GEN_25 = level != 2'h0 ? _T_342 : memRespStore; // @[EmbeddedTLB.scala 313:36 EmbeddedTLB.scala 321:24 EmbeddedTLB.scala 250:29]
  wire  _GEN_26 = level != 2'h0 ? _GEN_21 : missIPF; // @[EmbeddedTLB.scala 313:36 EmbeddedTLB.scala 266:24]
  wire [2:0] _GEN_27 = level != 2'h0 ? _GEN_22 : state; // @[EmbeddedTLB.scala 313:36 EmbeddedTLB.scala 247:22]
  wire  _GEN_28 = level != 2'h0 & _GEN_23; // @[EmbeddedTLB.scala 313:36]
  wire [17:0] _GEN_29 = level != 2'h0 ? _T_348 : 18'h3ffff; // @[EmbeddedTLB.scala 313:36 EmbeddedTLB.scala 339:20]
  wire [17:0] _GEN_37 = ~(_T_281[1] | _T_281[3]) & (level == 2'h3 | level == 2'h2) ? 18'h3ffff : _GEN_29; // @[EmbeddedTLB.scala 297:82]
  wire [17:0] _GEN_45 = isFlush ? 18'h3ffff : _GEN_37; // @[EmbeddedTLB.scala 294:24]
  wire [17:0] _GEN_54 = _T_290 ? _GEN_45 : 18'h3ffff; // @[EmbeddedTLB.scala 293:33]
  wire [17:0] _GEN_77 = _T_280 ? _GEN_54 : 18'h3ffff; // @[Conditional.scala 39:67]
  wire [17:0] _GEN_88 = _T_278 ? 18'h3ffff : _GEN_77; // @[Conditional.scala 39:67]
  wire [17:0] missMask = _T_272 ? 18'h3ffff : _GEN_88; // @[Conditional.scala 40:58]
  wire [17:0] _GEN_30 = level != 2'h0 ? missMask : missMaskStore; // @[EmbeddedTLB.scala 313:36 EmbeddedTLB.scala 340:25 EmbeddedTLB.scala 252:30]
  wire [2:0] _GEN_31 = ~(_T_281[1] | _T_281[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_18 : _GEN_27; // @[EmbeddedTLB.scala 297:82]
  wire  _GEN_32 = ~(_T_281[1] | _T_281[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_19 : _GEN_26; // @[EmbeddedTLB.scala 297:82]
  wire [31:0] _GEN_33 = ~(_T_281[1] | _T_281[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_20 : raddr; // @[EmbeddedTLB.scala 297:82 EmbeddedTLB.scala 256:22]
  wire [7:0] _GEN_34 = ~(_T_281[1] | _T_281[3]) & (level == 2'h3 | level == 2'h2) ? 8'h0 : _GEN_24; // @[EmbeddedTLB.scala 297:82]
  wire [63:0] _GEN_35 = ~(_T_281[1] | _T_281[3]) & (level == 2'h3 | level == 2'h2) ? memRespStore : _GEN_25; // @[EmbeddedTLB.scala 297:82 EmbeddedTLB.scala 250:29]
  wire  _GEN_36 = ~(_T_281[1] | _T_281[3]) & (level == 2'h3 | level == 2'h2) ? 1'h0 : _GEN_28; // @[EmbeddedTLB.scala 297:82]
  wire [17:0] _GEN_38 = ~(_T_281[1] | _T_281[3]) & (level == 2'h3 | level == 2'h2) ? missMaskStore : _GEN_30; // @[EmbeddedTLB.scala 297:82 EmbeddedTLB.scala 252:30]
  wire [2:0] _GEN_39 = isFlush ? 3'h0 : _GEN_31; // @[EmbeddedTLB.scala 294:24 EmbeddedTLB.scala 295:17]
  wire  _GEN_40 = isFlush ? missIPF : _GEN_32; // @[EmbeddedTLB.scala 294:24 EmbeddedTLB.scala 266:24]
  wire [31:0] _GEN_41 = isFlush ? raddr : _GEN_33; // @[EmbeddedTLB.scala 294:24 EmbeddedTLB.scala 256:22]
  wire [7:0] _GEN_42 = isFlush ? 8'h0 : _GEN_34; // @[EmbeddedTLB.scala 294:24]
  wire [63:0] _GEN_43 = isFlush ? memRespStore : _GEN_35; // @[EmbeddedTLB.scala 294:24 EmbeddedTLB.scala 250:29]
  wire  _GEN_44 = isFlush ? 1'h0 : _GEN_36; // @[EmbeddedTLB.scala 294:24]
  wire [17:0] _GEN_46 = isFlush ? missMaskStore : _GEN_38; // @[EmbeddedTLB.scala 294:24 EmbeddedTLB.scala 252:30]
  wire [1:0] _T_350 = level - 2'h1; // @[EmbeddedTLB.scala 342:24]
  wire [2:0] _GEN_47 = _T_290 ? _GEN_39 : state; // @[EmbeddedTLB.scala 293:33 EmbeddedTLB.scala 247:22]
  wire  _GEN_48 = _T_290 ? _GEN_17 : _GEN_4; // @[EmbeddedTLB.scala 293:33]
  wire  _GEN_49 = _T_290 ? _GEN_40 : missIPF; // @[EmbeddedTLB.scala 293:33 EmbeddedTLB.scala 266:24]
  wire [31:0] _GEN_50 = _T_290 ? _GEN_41 : raddr; // @[EmbeddedTLB.scala 293:33 EmbeddedTLB.scala 256:22]
  wire [7:0] _GEN_51 = _T_290 ? _GEN_42 : 8'h0; // @[EmbeddedTLB.scala 293:33]
  wire [63:0] _GEN_52 = _T_290 ? _GEN_43 : memRespStore; // @[EmbeddedTLB.scala 293:33 EmbeddedTLB.scala 250:29]
  wire  _GEN_53 = _T_290 & _GEN_44; // @[EmbeddedTLB.scala 293:33]
  wire [17:0] _GEN_55 = _T_290 ? _GEN_46 : missMaskStore; // @[EmbeddedTLB.scala 293:33 EmbeddedTLB.scala 252:30]
  wire [1:0] _GEN_56 = _T_290 ? _T_350 : level; // @[EmbeddedTLB.scala 293:33 EmbeddedTLB.scala 342:15 EmbeddedTLB.scala 248:22]
  wire  _T_351 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_57 = _T_279 ? 3'h4 : state; // @[EmbeddedTLB.scala 350:38 EmbeddedTLB.scala 350:46 EmbeddedTLB.scala 247:22]
  wire [2:0] _GEN_58 = isFlush ? 3'h0 : _GEN_57; // @[EmbeddedTLB.scala 347:22 EmbeddedTLB.scala 348:15]
  wire  _T_353 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_59 = _T_267 | io_flush | alreadyOutFire ? 3'h0 : state; // @[EmbeddedTLB.scala 353:73 EmbeddedTLB.scala 354:13 EmbeddedTLB.scala 247:22]
  wire  _GEN_60 = _T_267 | io_flush | alreadyOutFire ? 1'h0 : missIPF; // @[EmbeddedTLB.scala 353:73 EmbeddedTLB.scala 355:15 EmbeddedTLB.scala 266:24]
  wire  _GEN_61 = _T_267 | io_flush | alreadyOutFire ? 1'h0 : _GEN_2; // @[EmbeddedTLB.scala 353:73 EmbeddedTLB.scala 356:22]
  wire  _T_357 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_62 = _T_357 ? 3'h0 : state; // @[Conditional.scala 39:67 EmbeddedTLB.scala 360:13 EmbeddedTLB.scala 247:22]
  wire [2:0] _GEN_63 = _T_353 ? _GEN_59 : _GEN_62; // @[Conditional.scala 39:67]
  wire  _GEN_64 = _T_353 ? _GEN_60 : missIPF; // @[Conditional.scala 39:67 EmbeddedTLB.scala 266:24]
  wire  _GEN_65 = _T_353 ? _GEN_61 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_66 = _T_351 ? _GEN_58 : _GEN_63; // @[Conditional.scala 39:67]
  wire  _GEN_67 = _T_351 ? _GEN_17 : _GEN_4; // @[Conditional.scala 39:67]
  wire  _GEN_68 = _T_351 ? missIPF : _GEN_64; // @[Conditional.scala 39:67 EmbeddedTLB.scala 266:24]
  wire  _GEN_69 = _T_351 ? _GEN_2 : _GEN_65; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_74 = _T_280 ? _GEN_51 : 8'h0; // @[Conditional.scala 39:67]
  wire  _GEN_87 = _T_278 ? 1'h0 : _T_280 & _GEN_53; // @[Conditional.scala 39:67]
  wire  missMetaRefill = _T_272 ? 1'h0 : _GEN_87; // @[Conditional.scala 40:58]
  wire  cmd = state == 3'h3; // @[EmbeddedTLB.scala 365:23]
  wire  _T_364 = ~isFlush; // @[EmbeddedTLB.scala 367:77]
  wire  _T_368 = state == 3'h0; // @[EmbeddedTLB.scala 371:82]
  reg  REG_7; // @[EmbeddedTLB.scala 371:33]
  reg [3:0] REG_9; // @[EmbeddedTLB.scala 372:65]
  reg [26:0] hi_hi_hi; // @[EmbeddedTLB.scala 372:94]
  reg [15:0] hi_hi_lo; // @[EmbeddedTLB.scala 373:19]
  reg [17:0] hi_lo_4; // @[EmbeddedTLB.scala 373:77]
  reg [7:0] lo_hi_hi; // @[EmbeddedTLB.scala 374:19]
  reg [19:0] lo_hi_lo; // @[EmbeddedTLB.scala 374:82]
  reg [31:0] lo_lo_3; // @[EmbeddedTLB.scala 375:22]
  wire [59:0] lo_8 = {lo_hi_hi,lo_hi_lo,lo_lo_3}; // @[Cat.scala 30:58]
  wire [60:0] hi_16 = {hi_hi_hi,hi_hi_lo,hi_lo_4}; // @[Cat.scala 30:58]
  wire [31:0] _T_384 = {hitData_ppn,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_385 = {2'h3,hitMeta_mask,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_386 = _T_384 & _T_385; // @[BitUtils.scala 32:13]
  wire [31:0] _T_387 = ~_T_385; // @[BitUtils.scala 32:38]
  wire [31:0] _T_388 = io_in_bits_addr[31:0] & _T_387; // @[BitUtils.scala 32:36]
  wire [31:0] _T_389 = _T_386 | _T_388; // @[BitUtils.scala 32:25]
  wire [31:0] _T_402 = {memRespStore[29:10],12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_403 = {2'h3,missMaskStore,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_404 = _T_402 & _T_403; // @[BitUtils.scala 32:13]
  wire [31:0] _T_405 = ~_T_403; // @[BitUtils.scala 32:38]
  wire [31:0] _T_406 = io_in_bits_addr[31:0] & _T_405; // @[BitUtils.scala 32:36]
  wire [31:0] _T_407 = _T_404 | _T_406; // @[BitUtils.scala 32:25]
  wire  _T_409 = ~hitWB; // @[EmbeddedTLB.scala 380:45]
  wire  _T_416 = hit & ~hitWB ? _T_237 : state == 3'h4; // @[EmbeddedTLB.scala 380:37]
  assign io_in_ready = io_out_ready & _T_368 & ~miss & _T_409 & io_mdReady & _T_237; // @[EmbeddedTLB.scala 382:86]
  assign io_out_valid = io_in_valid & _T_416; // @[EmbeddedTLB.scala 380:31]
  assign io_out_bits_addr = hit ? _T_389 : _T_407; // @[EmbeddedTLB.scala 379:26]
  assign io_out_bits_size = io_in_bits_size; // @[EmbeddedTLB.scala 378:15]
  assign io_out_bits_user = io_in_bits_user; // @[EmbeddedTLB.scala 378:15]
  assign io_mdWrite_wen = REG_7; // @[TLB.scala 214:14]
  assign io_mdWrite_waymask = REG_9; // @[TLB.scala 216:18]
  assign io_mdWrite_wdata = {hi_16,lo_8}; // @[Cat.scala 30:58]
  assign io_mem_req_valid = (state == 3'h1 | cmd) & ~isFlush; // @[EmbeddedTLB.scala 367:74]
  assign io_mem_req_bits_addr = hitWB ? hitData_pteaddr : raddr; // @[EmbeddedTLB.scala 366:35]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[EmbeddedTLB.scala 365:23]
  assign io_mem_req_bits_wdata = hitWB ? {{24'd0}, hitWBStore} : memRespStore; // @[EmbeddedTLB.scala 366:138]
  assign io_mem_resp_ready = 1'h1; // @[EmbeddedTLB.scala 368:21]
  assign io_pf_loadPF = 1'h0; // @[EmbeddedTLB.scala 236:16]
  assign io_pf_storePF = 1'h0; // @[EmbeddedTLB.scala 237:17]
  assign io_ipf = hit ? hitinstrPF : missIPF; // @[EmbeddedTLB.scala 384:16]
  assign io_isFinish = _T_267 | _T_235; // @[EmbeddedTLB.scala 385:32]
  always @(posedge clock) begin
    if (reset) begin // @[LFSR64.scala 25:23]
      REG <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG == 64'h0) begin // @[LFSR64.scala 28:18]
      REG <= 64'h1;
    end else begin
      REG <= _T_183;
    end
    if (reset) begin // @[Reg.scala 27:20]
      hitWBStore <= 40'h0; // @[Reg.scala 27:20]
    end else if (hitWB) begin // @[Reg.scala 28:19]
      hitWBStore <= _T_240; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[EmbeddedTLB.scala 247:22]
      state <= 3'h0; // @[EmbeddedTLB.scala 247:22]
    end else if (_T_272) begin // @[Conditional.scala 40:58]
      if (~io_flush & hitWB) begin // @[EmbeddedTLB.scala 271:32]
        state <= 3'h3; // @[EmbeddedTLB.scala 272:15]
      end else if (miss & _T_273) begin // @[EmbeddedTLB.scala 275:37]
        state <= 3'h1; // @[EmbeddedTLB.scala 276:15]
      end
    end else if (_T_278) begin // @[Conditional.scala 39:67]
      if (isFlush) begin // @[EmbeddedTLB.scala 285:22]
        state <= 3'h0; // @[EmbeddedTLB.scala 286:15]
      end else begin
        state <= _GEN_15;
      end
    end else if (_T_280) begin // @[Conditional.scala 39:67]
      state <= _GEN_47;
    end else begin
      state <= _GEN_66;
    end
    if (reset) begin // @[EmbeddedTLB.scala 248:22]
      level <= 2'h3; // @[EmbeddedTLB.scala 248:22]
    end else if (_T_272) begin // @[Conditional.scala 40:58]
      if (!(~io_flush & hitWB)) begin // @[EmbeddedTLB.scala 271:32]
        if (miss & _T_273) begin // @[EmbeddedTLB.scala 275:37]
          level <= 2'h3; // @[EmbeddedTLB.scala 278:15]
        end
      end
    end else if (!(_T_278)) begin // @[Conditional.scala 39:67]
      if (_T_280) begin // @[Conditional.scala 39:67]
        level <= _GEN_56;
      end
    end
    if (reset) begin // @[EmbeddedTLB.scala 250:29]
      memRespStore <= 64'h0; // @[EmbeddedTLB.scala 250:29]
    end else if (!(_T_272)) begin // @[Conditional.scala 40:58]
      if (!(_T_278)) begin // @[Conditional.scala 39:67]
        if (_T_280) begin // @[Conditional.scala 39:67]
          memRespStore <= _GEN_52;
        end
      end
    end
    if (reset) begin // @[EmbeddedTLB.scala 252:30]
      missMaskStore <= 18'h0; // @[EmbeddedTLB.scala 252:30]
    end else if (!(_T_272)) begin // @[Conditional.scala 40:58]
      if (!(_T_278)) begin // @[Conditional.scala 39:67]
        if (_T_280) begin // @[Conditional.scala 39:67]
          missMaskStore <= _GEN_55;
        end
      end
    end
    if (reset) begin // @[EmbeddedTLB.scala 256:22]
      raddr <= 32'h0; // @[EmbeddedTLB.scala 256:22]
    end else if (_T_272) begin // @[Conditional.scala 40:58]
      if (!(~io_flush & hitWB)) begin // @[EmbeddedTLB.scala 271:32]
        if (miss & _T_273) begin // @[EmbeddedTLB.scala 275:37]
          raddr <= _T_277; // @[EmbeddedTLB.scala 277:15]
        end
      end
    end else if (!(_T_278)) begin // @[Conditional.scala 39:67]
      if (_T_280) begin // @[Conditional.scala 39:67]
        raddr <= _GEN_50;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      alreadyOutFire <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_272) begin // @[Conditional.scala 40:58]
      if (~io_flush & hitWB) begin // @[EmbeddedTLB.scala 271:32]
        alreadyOutFire <= 1'h0; // @[EmbeddedTLB.scala 274:24]
      end else if (miss & _T_273) begin // @[EmbeddedTLB.scala 275:37]
        alreadyOutFire <= 1'h0; // @[EmbeddedTLB.scala 280:24]
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else if (_T_278) begin // @[Conditional.scala 39:67]
      alreadyOutFire <= _GEN_2;
    end else if (_T_280) begin // @[Conditional.scala 39:67]
      alreadyOutFire <= _GEN_2;
    end else begin
      alreadyOutFire <= _GEN_69;
    end
    if (reset) begin // @[EmbeddedTLB.scala 260:26]
      needFlush <= 1'h0; // @[EmbeddedTLB.scala 260:26]
    end else if (_T_272) begin // @[Conditional.scala 40:58]
      if (~io_flush & hitWB) begin // @[EmbeddedTLB.scala 271:32]
        needFlush <= 1'h0; // @[EmbeddedTLB.scala 273:19]
      end else if (miss & _T_273) begin // @[EmbeddedTLB.scala 275:37]
        needFlush <= 1'h0; // @[EmbeddedTLB.scala 279:19]
      end else begin
        needFlush <= _GEN_4;
      end
    end else if (_T_278) begin // @[Conditional.scala 39:67]
      if (isFlush) begin // @[EmbeddedTLB.scala 285:22]
        needFlush <= 1'h0; // @[EmbeddedTLB.scala 287:19]
      end else begin
        needFlush <= _GEN_4;
      end
    end else if (_T_280) begin // @[Conditional.scala 39:67]
      needFlush <= _GEN_48;
    end else begin
      needFlush <= _GEN_67;
    end
    if (reset) begin // @[EmbeddedTLB.scala 266:24]
      missIPF <= 1'h0; // @[EmbeddedTLB.scala 266:24]
    end else if (!(_T_272)) begin // @[Conditional.scala 40:58]
      if (!(_T_278)) begin // @[Conditional.scala 39:67]
        if (_T_280) begin // @[Conditional.scala 39:67]
          missIPF <= _GEN_49;
        end else begin
          missIPF <= _GEN_68;
        end
      end
    end
    if (reset) begin // @[EmbeddedTLB.scala 371:33]
      REG_7 <= 1'h0; // @[EmbeddedTLB.scala 371:33]
    end else begin
      REG_7 <= missMetaRefill & _T_364 | hitWB & state == 3'h0 & _T_364; // @[EmbeddedTLB.scala 371:33]
    end
    if (reset) begin // @[EmbeddedTLB.scala 372:65]
      REG_9 <= 4'h0; // @[EmbeddedTLB.scala 372:65]
    end else if (hit) begin // @[EmbeddedTLB.scala 209:20]
      REG_9 <= hitVec;
    end else begin
      REG_9 <= victimWaymask;
    end
    if (reset) begin // @[EmbeddedTLB.scala 372:94]
      hi_hi_hi <= 27'h0; // @[EmbeddedTLB.scala 372:94]
    end else begin
      hi_hi_hi <= _T_43; // @[EmbeddedTLB.scala 372:94]
    end
    if (reset) begin // @[EmbeddedTLB.scala 373:19]
      hi_hi_lo <= 16'h0; // @[EmbeddedTLB.scala 373:19]
    end else if (hitWB) begin // @[EmbeddedTLB.scala 373:23]
      hi_hi_lo <= hitMeta_asid;
    end else begin
      hi_hi_lo <= satp_asid;
    end
    if (reset) begin // @[EmbeddedTLB.scala 373:77]
      hi_lo_4 <= 18'h0; // @[EmbeddedTLB.scala 373:77]
    end else if (hitWB) begin // @[EmbeddedTLB.scala 373:81]
      hi_lo_4 <= hitMeta_mask;
    end else if (_T_272) begin // @[Conditional.scala 40:58]
      hi_lo_4 <= 18'h3ffff;
    end else if (_T_278) begin // @[Conditional.scala 39:67]
      hi_lo_4 <= 18'h3ffff;
    end else begin
      hi_lo_4 <= _GEN_77;
    end
    if (reset) begin // @[EmbeddedTLB.scala 374:19]
      lo_hi_hi <= 8'h0; // @[EmbeddedTLB.scala 374:19]
    end else if (hitWB) begin // @[EmbeddedTLB.scala 374:23]
      lo_hi_hi <= hitRefillFlag;
    end else if (_T_272) begin // @[Conditional.scala 40:58]
      lo_hi_hi <= 8'h0;
    end else if (_T_278) begin // @[Conditional.scala 39:67]
      lo_hi_hi <= 8'h0;
    end else begin
      lo_hi_hi <= _GEN_74;
    end
    if (reset) begin // @[EmbeddedTLB.scala 374:82]
      lo_hi_lo <= 20'h0; // @[EmbeddedTLB.scala 374:82]
    end else if (hitWB) begin // @[EmbeddedTLB.scala 374:86]
      lo_hi_lo <= hitData_ppn;
    end else begin
      lo_hi_lo <= memRdata_ppn;
    end
    if (reset) begin // @[EmbeddedTLB.scala 375:22]
      lo_lo_3 <= 32'h0; // @[EmbeddedTLB.scala 375:22]
    end else if (hitWB) begin // @[EmbeddedTLB.scala 366:35]
      lo_lo_3 <= hitData_pteaddr;
    end else begin
      lo_lo_3 <= raddr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  REG = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  hitWBStore = _RAND_1[39:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  level = _RAND_3[1:0];
  _RAND_4 = {2{`RANDOM}};
  memRespStore = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  missMaskStore = _RAND_5[17:0];
  _RAND_6 = {1{`RANDOM}};
  raddr = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  alreadyOutFire = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  needFlush = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  missIPF = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  REG_7 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG_9 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  hi_hi_hi = _RAND_12[26:0];
  _RAND_13 = {1{`RANDOM}};
  hi_hi_lo = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  hi_lo_4 = _RAND_14[17:0];
  _RAND_15 = {1{`RANDOM}};
  lo_hi_hi = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  lo_hi_lo = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  lo_lo_3 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_EmbeddedTLBMD(
  input          clock,
  input          reset,
  output [120:0] io_tlbmd_0,
  output [120:0] io_tlbmd_1,
  output [120:0] io_tlbmd_2,
  output [120:0] io_tlbmd_3,
  input          io_write_wen,
  input  [3:0]   io_write_waymask,
  input  [120:0] io_write_wdata,
  output         io_ready
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [120:0] tlbmd_0 [0:0]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_0_MPORT_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0_MPORT_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_0_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0_MPORT_1_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0_MPORT_1_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0_MPORT_1_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_1 [0:0]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_1_MPORT_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1_MPORT_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_1_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1_MPORT_1_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1_MPORT_1_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1_MPORT_1_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_2 [0:0]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_2_MPORT_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2_MPORT_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_2_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2_MPORT_1_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2_MPORT_1_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2_MPORT_1_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_3 [0:0]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_3_MPORT_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3_MPORT_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_3_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3_MPORT_1_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3_MPORT_1_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3_MPORT_1_en; // @[EmbeddedTLB.scala 38:18]
  reg  resetState; // @[EmbeddedTLB.scala 42:27]
  wire  _GEN_1 = resetState ? 1'h0 : resetState; // @[EmbeddedTLB.scala 44:22 EmbeddedTLB.scala 44:35 EmbeddedTLB.scala 42:27]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[EmbeddedTLB.scala 53:20]
  assign tlbmd_0_MPORT_addr = 1'h0;
  assign tlbmd_0_MPORT_data = tlbmd_0[tlbmd_0_MPORT_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_0_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_0_MPORT_1_addr = 1'h0;
  assign tlbmd_0_MPORT_1_mask = waymask[0];
  assign tlbmd_0_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_1_MPORT_addr = 1'h0;
  assign tlbmd_1_MPORT_data = tlbmd_1[tlbmd_1_MPORT_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_1_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_1_MPORT_1_addr = 1'h0;
  assign tlbmd_1_MPORT_1_mask = waymask[1];
  assign tlbmd_1_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_2_MPORT_addr = 1'h0;
  assign tlbmd_2_MPORT_data = tlbmd_2[tlbmd_2_MPORT_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_2_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_2_MPORT_1_addr = 1'h0;
  assign tlbmd_2_MPORT_1_mask = waymask[2];
  assign tlbmd_2_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_3_MPORT_addr = 1'h0;
  assign tlbmd_3_MPORT_data = tlbmd_3[tlbmd_3_MPORT_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_3_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_3_MPORT_1_addr = 1'h0;
  assign tlbmd_3_MPORT_1_mask = waymask[3];
  assign tlbmd_3_MPORT_1_en = resetState | io_write_wen;
  assign io_tlbmd_0 = tlbmd_0_MPORT_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_1 = tlbmd_1_MPORT_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_2 = tlbmd_2_MPORT_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_3 = tlbmd_3_MPORT_data; // @[EmbeddedTLB.scala 39:12]
  assign io_ready = ~resetState; // @[EmbeddedTLB.scala 59:15]
  always @(posedge clock) begin
    if(tlbmd_0_MPORT_1_en & tlbmd_0_MPORT_1_mask) begin
      tlbmd_0[tlbmd_0_MPORT_1_addr] <= tlbmd_0_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_1_MPORT_1_en & tlbmd_1_MPORT_1_mask) begin
      tlbmd_1[tlbmd_1_MPORT_1_addr] <= tlbmd_1_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_2_MPORT_1_en & tlbmd_2_MPORT_1_mask) begin
      tlbmd_2[tlbmd_2_MPORT_1_addr] <= tlbmd_2_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_3_MPORT_1_en & tlbmd_3_MPORT_1_mask) begin
      tlbmd_3[tlbmd_3_MPORT_1_addr] <= tlbmd_3_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
    end
    resetState <= reset | _GEN_1; // @[EmbeddedTLB.scala 42:27 EmbeddedTLB.scala 42:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[120:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_EmbeddedTLB(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [86:0] io_in_req_bits_user,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output [86:0] io_in_resp_bits_user,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [86:0] io_out_req_bits_user,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input  [86:0] io_out_resp_bits_user,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  input         io_mem_resp_valid,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_flush,
  input  [1:0]  io_csrMMU_priviledgeMode,
  input         io_cacheEmpty,
  output        io_ipf,
  input  [63:0] CSRSATP,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [95:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_reset; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_in_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_in_valid; // @[EmbeddedTLB.scala 80:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [2:0] tlbExec_io_in_bits_size; // @[EmbeddedTLB.scala 80:23]
  wire [86:0] tlbExec_io_in_bits_user; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_out_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_out_valid; // @[EmbeddedTLB.scala 80:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [2:0] tlbExec_io_out_bits_size; // @[EmbeddedTLB.scala 80:23]
  wire [86:0] tlbExec_io_out_bits_user; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_0; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_1; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_2; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_3; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mdReady; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_req_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 80:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_resp_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_resp_valid; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_flush; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_satp; // @[EmbeddedTLB.scala 80:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_ipf; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_isFinish; // @[EmbeddedTLB.scala 80:23]
  wire  mdTLB_clock; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_reset; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_0; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_1; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_2; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_3; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_io_write_wen; // @[EmbeddedTLB.scala 82:21]
  wire [3:0] mdTLB_io_write_waymask; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_write_wdata; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_io_ready; // @[EmbeddedTLB.scala 82:21]
  reg [120:0] REG__0; // @[Reg.scala 27:20]
  reg [120:0] REG__1; // @[Reg.scala 27:20]
  reg [120:0] REG__2; // @[Reg.scala 27:20]
  reg [120:0] REG__3; // @[Reg.scala 27:20]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[EmbeddedTLB.scala 114:26]
  wire  vmEnable = CSRSATP[63:60] == 4'h8 & io_csrMMU_priviledgeMode < 2'h3; // @[EmbeddedTLB.scala 102:57]
  reg  REG_1; // @[EmbeddedTLB.scala 105:24]
  wire  _GEN_4 = tlbExec_io_isFinish ? 1'h0 : REG_1; // @[EmbeddedTLB.scala 106:25 EmbeddedTLB.scala 106:33 EmbeddedTLB.scala 105:24]
  wire  _GEN_5 = mdUpdate & vmEnable | _GEN_4; // @[EmbeddedTLB.scala 107:50 EmbeddedTLB.scala 107:58]
  reg [38:0] REG_2_addr; // @[Reg.scala 27:20]
  reg [2:0] REG_2_size; // @[Reg.scala 27:20]
  reg [86:0] REG_2_user; // @[Reg.scala 27:20]
  wire  _GEN_13 = ~vmEnable | io_out_req_ready; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 124:26 EmbeddedTLB.scala 136:23]
  wire  _GEN_14 = ~vmEnable ? io_in_req_valid : tlbExec_io_out_valid; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 126:22 EmbeddedTLB.scala 136:23]
  wire  _T_17 = tlbExec_io_ipf & vmEnable; // @[EmbeddedTLB.scala 152:26]
  ysyx_210000_EmbeddedTLBExec tlbExec ( // @[EmbeddedTLB.scala 80:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_size(tlbExec_io_in_bits_size),
    .io_in_bits_user(tlbExec_io_in_bits_user),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_size(tlbExec_io_out_bits_size),
    .io_out_bits_user(tlbExec_io_out_bits_user),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_flush(tlbExec_io_flush),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_ipf(tlbExec_io_ipf),
    .io_isFinish(tlbExec_io_isFinish)
  );
  ysyx_210000_EmbeddedTLBMD mdTLB ( // @[EmbeddedTLB.scala 82:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_ready(mdTLB_io_ready)
  );
  assign io_in_req_ready = ~vmEnable ? io_out_req_ready : tlbExec_io_in_ready; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 127:21 EmbeddedTLB.scala 110:16]
  assign io_in_resp_valid = _T_17 & io_cacheEmpty | io_out_resp_valid; // @[EmbeddedTLB.scala 157:56 EmbeddedTLB.scala 158:24 EmbeddedTLB.scala 138:15]
  assign io_in_resp_bits_rdata = _T_17 & io_cacheEmpty ? 64'h0 : io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 157:56 EmbeddedTLB.scala 159:29 EmbeddedTLB.scala 138:15]
  assign io_in_resp_bits_user = _T_17 & io_cacheEmpty ? tlbExec_io_in_bits_user : io_out_resp_bits_user; // @[EmbeddedTLB.scala 157:56 EmbeddedTLB.scala 161:34 EmbeddedTLB.scala 138:15]
  assign io_out_req_valid = tlbExec_io_ipf & vmEnable ? 1'h0 : _GEN_14; // @[EmbeddedTLB.scala 152:39 EmbeddedTLB.scala 154:24]
  assign io_out_req_bits_addr = ~vmEnable ? io_in_req_bits_addr[31:0] : tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 128:26 EmbeddedTLB.scala 136:23]
  assign io_out_req_bits_size = ~vmEnable ? 3'h3 : tlbExec_io_out_bits_size; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 129:26 EmbeddedTLB.scala 136:23]
  assign io_out_req_bits_user = ~vmEnable ? io_in_req_bits_user : tlbExec_io_out_bits_user; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 133:32 EmbeddedTLB.scala 136:23]
  assign io_out_resp_ready = io_in_resp_ready; // @[EmbeddedTLB.scala 138:15]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 87:18]
  assign io_ipf = _T_17 & io_cacheEmpty & tlbExec_io_ipf; // @[EmbeddedTLB.scala 157:56 EmbeddedTLB.scala 162:14 EmbeddedTLB.scala 94:10]
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = REG_1; // @[EmbeddedTLB.scala 112:17]
  assign tlbExec_io_in_bits_addr = REG_2_addr; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_size = REG_2_size; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_user = REG_2_user; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_out_ready = tlbExec_io_ipf & vmEnable ? io_cacheEmpty & io_in_resp_ready : _GEN_13; // @[EmbeddedTLB.scala 152:39 EmbeddedTLB.scala 153:28]
  assign tlbExec_io_md_0 = REG__0; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_1 = REG__1; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_2 = REG__2; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_3 = REG__3; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[EmbeddedTLB.scala 90:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_flush = io_flush; // @[EmbeddedTLB.scala 85:20]
  assign tlbExec_io_satp = CSRSATP; // @[EmbeddedTLB.scala 86:19]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 88:17]
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[EmbeddedTLB.scala 99:31]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 92:18]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      REG__0 <= 121'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG__0 <= mdTLB_io_tlbmd_0; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG__1 <= 121'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG__1 <= mdTLB_io_tlbmd_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG__2 <= 121'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG__2 <= mdTLB_io_tlbmd_2; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG__3 <= 121'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG__3 <= mdTLB_io_tlbmd_3; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[EmbeddedTLB.scala 105:24]
      REG_1 <= 1'h0; // @[EmbeddedTLB.scala 105:24]
    end else if (io_flush) begin // @[EmbeddedTLB.scala 108:20]
      REG_1 <= 1'h0; // @[EmbeddedTLB.scala 108:28]
    end else begin
      REG_1 <= _GEN_5;
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_2_addr <= 39'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG_2_addr <= io_in_req_bits_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_2_size <= 3'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG_2_size <= 3'h3; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_2_user <= 87'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG_2_user <= io_in_req_bits_user; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  REG__0 = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  REG__1 = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  REG__2 = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  REG__3 = _RAND_3[120:0];
  _RAND_4 = {1{`RANDOM}};
  REG_1 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  REG_2_addr = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  REG_2_size = _RAND_6[2:0];
  _RAND_7 = {3{`RANDOM}};
  REG_2_user = _RAND_7[86:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_CacheStage1(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [86:0] io_in_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [86:0] io_out_bits_req_user,
  input         io_metaReadBus_req_ready,
  output        io_metaReadBus_req_valid,
  output [3:0]  io_metaReadBus_req_bits_setIdx,
  input  [21:0] io_metaReadBus_resp_data_0_tag,
  input         io_metaReadBus_resp_data_0_valid,
  input  [21:0] io_metaReadBus_resp_data_1_tag,
  input         io_metaReadBus_resp_data_1_valid,
  input  [21:0] io_metaReadBus_resp_data_2_tag,
  input         io_metaReadBus_resp_data_2_valid,
  input  [21:0] io_metaReadBus_resp_data_3_tag,
  input         io_metaReadBus_resp_data_3_valid,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [6:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data
);
  wire  _T_26 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = (~io_in_valid | _T_26) & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 134:78]
  assign io_out_valid = io_in_valid & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 133:59]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[Cache.scala 132:19]
  assign io_out_bits_req_size = io_in_bits_size; // @[Cache.scala 132:19]
  assign io_out_bits_req_user = io_in_bits_user; // @[Cache.scala 132:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 128:34]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[9:6]; // @[Cache.scala 79:45]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 128:34]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[9:6],io_in_bits_addr[5:3]}; // @[Cat.scala 30:58]
endmodule
module ysyx_210000_CacheStage2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [86:0] io_in_bits_req_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [86:0] io_out_bits_req_user,
  output [21:0] io_out_bits_metas_0_tag,
  output [21:0] io_out_bits_metas_1_tag,
  output [21:0] io_out_bits_metas_2_tag,
  output [21:0] io_out_bits_metas_3_tag,
  output [63:0] io_out_bits_datas_0_data,
  output [63:0] io_out_bits_datas_1_data,
  output [63:0] io_out_bits_datas_2_data,
  output [63:0] io_out_bits_datas_3_data,
  output        io_out_bits_hit,
  output [3:0]  io_out_bits_waymask,
  output        io_out_bits_mmio,
  output        io_out_bits_isForwardData,
  output [63:0] io_out_bits_forwardData_data_data,
  output [3:0]  io_out_bits_forwardData_waymask,
  input  [21:0] io_metaReadResp_0_tag,
  input         io_metaReadResp_0_valid,
  input  [21:0] io_metaReadResp_1_tag,
  input         io_metaReadResp_1_valid,
  input  [21:0] io_metaReadResp_2_tag,
  input         io_metaReadResp_2_valid,
  input  [21:0] io_metaReadResp_3_tag,
  input         io_metaReadResp_3_valid,
  input  [63:0] io_dataReadResp_0_data,
  input  [63:0] io_dataReadResp_1_data,
  input  [63:0] io_dataReadResp_2_data,
  input  [63:0] io_dataReadResp_3_data,
  input         io_metaWriteBus_req_valid,
  input  [3:0]  io_metaWriteBus_req_bits_setIdx,
  input  [21:0] io_metaWriteBus_req_bits_data_tag,
  input  [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_dataWriteBus_req_valid,
  input  [6:0]  io_dataWriteBus_req_bits_setIdx,
  input  [63:0] io_dataWriteBus_req_bits_data_data,
  input  [3:0]  io_dataWriteBus_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 162:31]
  wire [3:0] addr_index = io_in_bits_req_addr[9:6]; // @[Cache.scala 162:31]
  wire [21:0] addr_tag = io_in_bits_req_addr[31:10]; // @[Cache.scala 162:31]
  wire  isForwardMeta = io_in_valid & io_metaWriteBus_req_valid & io_metaWriteBus_req_bits_setIdx == addr_index; // @[Cache.scala 164:64]
  reg  isForwardMetaReg; // @[Cache.scala 165:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[Cache.scala 166:24 Cache.scala 166:43 Cache.scala 165:33]
  wire  _T_10 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_11 = ~io_in_valid; // @[Cache.scala 167:25]
  wire  _T_12 = _T_10 | ~io_in_valid; // @[Cache.scala 167:22]
  reg [21:0] forwardMetaReg_data_tag; // @[Reg.scala 27:20]
  reg  forwardMetaReg_data_valid; // @[Reg.scala 27:20]
  reg [3:0] forwardMetaReg_waymask; // @[Reg.scala 27:20]
  wire [3:0] _GEN_2 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _GEN_4 = isForwardMeta | forwardMetaReg_data_valid; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [21:0] _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[Cache.scala 171:42]
  wire  forwardWaymask_0 = _GEN_2[0]; // @[Cache.scala 173:61]
  wire  forwardWaymask_1 = _GEN_2[1]; // @[Cache.scala 173:61]
  wire  forwardWaymask_2 = _GEN_2[2]; // @[Cache.scala 173:61]
  wire  forwardWaymask_3 = _GEN_2[3]; // @[Cache.scala 173:61]
  wire [21:0] metaWay_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 175:22]
  wire  metaWay_0_valid = pickForwardMeta & forwardWaymask_0 ? _GEN_4 : io_metaReadResp_0_valid; // @[Cache.scala 175:22]
  wire [21:0] metaWay_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 175:22]
  wire  metaWay_1_valid = pickForwardMeta & forwardWaymask_1 ? _GEN_4 : io_metaReadResp_1_valid; // @[Cache.scala 175:22]
  wire [21:0] metaWay_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 175:22]
  wire  metaWay_2_valid = pickForwardMeta & forwardWaymask_2 ? _GEN_4 : io_metaReadResp_2_valid; // @[Cache.scala 175:22]
  wire [21:0] metaWay_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 175:22]
  wire  metaWay_3_valid = pickForwardMeta & forwardWaymask_3 ? _GEN_4 : io_metaReadResp_3_valid; // @[Cache.scala 175:22]
  wire  _T_23 = metaWay_0_valid & metaWay_0_tag == addr_tag & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_26 = metaWay_1_valid & metaWay_1_tag == addr_tag & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_29 = metaWay_2_valid & metaWay_2_tag == addr_tag & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_32 = metaWay_3_valid & metaWay_3_tag == addr_tag & io_in_valid; // @[Cache.scala 178:73]
  wire [3:0] hitVec = {_T_32,_T_29,_T_26,_T_23}; // @[Cache.scala 178:90]
  reg [63:0] REG; // @[LFSR64.scala 25:23]
  wire  hi_1 = REG[0] ^ REG[1] ^ REG[3] ^ REG[4]; // @[LFSR64.scala 26:43]
  wire [62:0] lo_1 = REG[63:1]; // @[LFSR64.scala 28:51]
  wire [63:0] _T_40 = {hi_1,lo_1}; // @[Cat.scala 30:58]
  wire [3:0] victimWaymask = 4'h1 << REG[1:0]; // @[Cache.scala 179:42]
  wire  _T_43 = ~metaWay_0_valid; // @[Cache.scala 181:45]
  wire  _T_44 = ~metaWay_1_valid; // @[Cache.scala 181:45]
  wire  _T_45 = ~metaWay_2_valid; // @[Cache.scala 181:45]
  wire  _T_46 = ~metaWay_3_valid; // @[Cache.scala 181:45]
  wire [3:0] invalidVec = {_T_46,_T_45,_T_44,_T_43}; // @[Cache.scala 181:56]
  wire  hasInvalidWay = |invalidVec; // @[Cache.scala 182:34]
  wire [1:0] _T_50 = invalidVec >= 4'h2 ? 2'h2 : 2'h1; // @[Cache.scala 185:8]
  wire [2:0] _T_51 = invalidVec >= 4'h4 ? 3'h4 : {{1'd0}, _T_50}; // @[Cache.scala 184:8]
  wire [3:0] refillInvalidWaymask = invalidVec >= 4'h8 ? 4'h8 : {{1'd0}, _T_51}; // @[Cache.scala 183:33]
  wire [3:0] _T_52 = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[Cache.scala 188:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _T_52; // @[Cache.scala 188:20]
  wire [1:0] _T_57 = waymask[0] + waymask[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_59 = waymask[2] + waymask[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_61 = _T_57 + _T_59; // @[Bitwise.scala 47:55]
  wire  _T_63 = _T_61 > 3'h1; // @[Cache.scala 189:26]
  wire  _T_127 = io_in_bits_req_addr < 32'h10000000; // @[NutCore.scala 115:32]
  wire  _T_131 = io_in_bits_req_addr >= 32'h10000000 & io_in_bits_req_addr < 32'h80000000; // @[NutCore.scala 115:24]
  wire [6:0] _T_141 = {addr_index,addr_wordIndex}; // @[Cat.scala 30:58]
  wire  _T_143 = io_dataWriteBus_req_valid & io_dataWriteBus_req_bits_setIdx == _T_141; // @[Cache.scala 205:13]
  wire  isForwardData = io_in_valid & _T_143; // @[Cache.scala 204:35]
  reg  isForwardDataReg; // @[Cache.scala 207:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[Cache.scala 208:24 Cache.scala 208:43 Cache.scala 207:33]
  reg [63:0] forwardDataReg_data_data; // @[Reg.scala 27:20]
  reg [3:0] forwardDataReg_waymask; // @[Reg.scala 27:20]
  wire  _T_150 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = _T_11 | _T_150; // @[Cache.scala 216:31]
  assign io_out_valid = io_in_valid; // @[Cache.scala 215:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[Cache.scala 214:19]
  assign io_out_bits_req_size = io_in_bits_req_size; // @[Cache.scala 214:19]
  assign io_out_bits_req_user = io_in_bits_req_user; // @[Cache.scala 214:19]
  assign io_out_bits_metas_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 175:22]
  assign io_out_bits_metas_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 175:22]
  assign io_out_bits_metas_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 175:22]
  assign io_out_bits_metas_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 175:22]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[Cache.scala 201:21]
  assign io_out_bits_hit = io_in_valid & |hitVec; // @[Cache.scala 199:34]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _T_52; // @[Cache.scala 188:20]
  assign io_out_bits_mmio = _T_127 | _T_131; // @[NutCore.scala 116:15]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[Cache.scala 211:49]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data :
    forwardDataReg_data_data; // @[Cache.scala 212:33]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[Cache.scala 212:33]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 165:33]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 165:33]
    end else if (_T_10 | ~io_in_valid) begin // @[Cache.scala 167:39]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 167:58]
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (reset) begin // @[Reg.scala 27:20]
      forwardMetaReg_data_tag <= 22'h0; // @[Reg.scala 27:20]
    end else if (isForwardMeta) begin // @[Reg.scala 28:19]
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      forwardMetaReg_data_valid <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      forwardMetaReg_data_valid <= _GEN_4;
    end
    if (reset) begin // @[Reg.scala 27:20]
      forwardMetaReg_waymask <= 4'h0; // @[Reg.scala 27:20]
    end else if (isForwardMeta) begin // @[Reg.scala 28:19]
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      REG <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG == 64'h0) begin // @[LFSR64.scala 28:18]
      REG <= 64'h1;
    end else begin
      REG <= _T_40;
    end
    if (reset) begin // @[Cache.scala 207:33]
      isForwardDataReg <= 1'h0; // @[Cache.scala 207:33]
    end else if (_T_12) begin // @[Cache.scala 209:39]
      isForwardDataReg <= 1'h0; // @[Cache.scala 209:58]
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (reset) begin // @[Reg.scala 27:20]
      forwardDataReg_data_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (isForwardData) begin // @[Reg.scala 28:19]
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      forwardDataReg_waymask <= 4'h0; // @[Reg.scala 27:20]
    end else if (isForwardData) begin // @[Reg.scala 28:19]
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask; // @[Reg.scala 28:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_in_valid & _T_63) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:196 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[Cache.scala 196:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_valid & _T_63) | reset)) begin
          $fatal; // @[Cache.scala 196:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  REG = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  isForwardDataReg = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_Arbiter(
  input         io_in_0_valid,
  input  [3:0]  io_in_0_bits_setIdx,
  input  [21:0] io_in_0_bits_data_tag,
  input         io_in_0_bits_data_dirty,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [3:0]  io_in_1_bits_setIdx,
  input  [21:0] io_in_1_bits_data_tag,
  input         io_in_1_bits_data_dirty,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [3:0]  io_out_bits_setIdx,
  output [21:0] io_out_bits_data_tag,
  output        io_out_bits_data_dirty,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  assign io_out_bits_data_tag = io_in_0_valid ? io_in_0_bits_data_tag : io_in_1_bits_data_tag; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  assign io_out_bits_data_dirty = io_in_0_valid ? io_in_0_bits_data_dirty : io_in_1_bits_data_dirty; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
endmodule
module ysyx_210000_Arbiter_1(
  input         io_in_0_valid,
  input  [6:0]  io_in_0_bits_setIdx,
  input  [63:0] io_in_0_bits_data_data,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [6:0]  io_in_1_bits_setIdx,
  input  [63:0] io_in_1_bits_data_data,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [6:0]  io_out_bits_setIdx,
  output [63:0] io_out_bits_data_data,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  assign io_out_bits_data_data = io_in_0_valid ? io_in_0_bits_data_data : io_in_1_bits_data_data; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
endmodule
module ysyx_210000_CacheStage3(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [86:0] io_in_bits_req_user,
  input  [21:0] io_in_bits_metas_0_tag,
  input  [21:0] io_in_bits_metas_1_tag,
  input  [21:0] io_in_bits_metas_2_tag,
  input  [21:0] io_in_bits_metas_3_tag,
  input  [63:0] io_in_bits_datas_0_data,
  input  [63:0] io_in_bits_datas_1_data,
  input  [63:0] io_in_bits_datas_2_data,
  input  [63:0] io_in_bits_datas_3_data,
  input         io_in_bits_hit,
  input  [3:0]  io_in_bits_waymask,
  input         io_in_bits_mmio,
  input         io_in_bits_isForwardData,
  input  [63:0] io_in_bits_forwardData_data_data,
  input  [3:0]  io_in_bits_forwardData_waymask,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_rdata,
  output [86:0] io_out_bits_user,
  output        io_isFinish,
  input         io_flush,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [6:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  output        io_dataWriteBus_req_valid,
  output [6:0]  io_dataWriteBus_req_bits_setIdx,
  output [63:0] io_dataWriteBus_req_bits_data_data,
  output [3:0]  io_dataWriteBus_req_bits_waymask,
  output        io_metaWriteBus_req_valid,
  output [3:0]  io_metaWriteBus_req_bits_setIdx,
  output [21:0] io_metaWriteBus_req_bits_data_tag,
  output        io_metaWriteBus_req_bits_data_dirty,
  output [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  output        io_mem_resp_ready,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output        io_mmio_resp_ready,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_cohResp_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 241:28]
  wire [21:0] metaWriteArb_io_in_0_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_0_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_valid; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 241:28]
  wire [21:0] metaWriteArb_io_in_1_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_valid; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 241:28]
  wire [21:0] metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[Cache.scala 241:28]
  wire  dataWriteArb_io_in_0_valid; // @[Cache.scala 242:28]
  wire [6:0] dataWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_in_1_valid; // @[Cache.scala 242:28]
  wire [6:0] dataWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_out_valid; // @[Cache.scala 242:28]
  wire [6:0] dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[Cache.scala 242:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 245:31]
  wire [3:0] addr_index = io_in_bits_req_addr[9:6]; // @[Cache.scala 245:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[Cache.scala 246:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[Cache.scala 247:25]
  wire  miss = io_in_valid & ~io_in_bits_hit; // @[Cache.scala 248:26]
  wire [21:0] _T_26 = io_in_bits_waymask[0] ? io_in_bits_metas_0_tag : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_27 = io_in_bits_waymask[1] ? io_in_bits_metas_1_tag : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_28 = io_in_bits_waymask[2] ? io_in_bits_metas_2_tag : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_29 = io_in_bits_waymask[3] ? io_in_bits_metas_3_tag : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_30 = _T_26 | _T_27; // @[Mux.scala 27:72]
  wire [21:0] _T_31 = _T_30 | _T_28; // @[Mux.scala 27:72]
  wire [21:0] meta_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  wire  useForwardData = io_in_bits_isForwardData & io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[Cache.scala 260:49]
  wire [63:0] _T_43 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_44 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_47 = _T_43 | _T_44; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = _T_47 | _T_45; // @[Mux.scala 27:72]
  wire [63:0] _T_49 = _T_48 | _T_46; // @[Mux.scala 27:72]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _T_49; // @[Cache.scala 262:21]
  wire  _T_70 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg [3:0] state; // @[Cache.scala 281:22]
  reg  needFlush; // @[Cache.scala 282:26]
  wire  _GEN_1 = io_flush & state != 4'h0 | needFlush; // @[Cache.scala 284:41 Cache.scala 284:53 Cache.scala 282:26]
  reg [2:0] value_1; // @[Counter.scala 60:40]
  reg [2:0] value_2; // @[Counter.scala 60:40]
  reg [1:0] state2; // @[Cache.scala 291:23]
  wire  _T_95 = state == 4'h3; // @[Cache.scala 293:39]
  wire  _T_96 = state == 4'h8; // @[Cache.scala 293:66]
  wire [2:0] lo_2 = _T_96 ? value_1 : value_2; // @[Cache.scala 294:33]
  wire  _T_102 = state2 == 2'h1; // @[Cache.scala 295:105]
  reg [63:0] dataWay_0_data; // @[Reg.scala 27:20]
  reg [63:0] dataWay_1_data; // @[Reg.scala 27:20]
  reg [63:0] dataWay_2_data; // @[Reg.scala 27:20]
  reg [63:0] dataWay_3_data; // @[Reg.scala 27:20]
  wire [63:0] _T_107 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_108 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_109 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_110 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_111 = _T_107 | _T_108; // @[Mux.scala 27:72]
  wire [63:0] _T_112 = _T_111 | _T_109; // @[Mux.scala 27:72]
  wire  _T_114 = 2'h0 == state2; // @[Conditional.scala 37:30]
  wire  _T_115 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_116 = 2'h1 == state2; // @[Conditional.scala 37:30]
  wire  _T_117 = 2'h2 == state2; // @[Conditional.scala 37:30]
  wire  _T_118 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_8 = _T_118 | io_cohResp_valid ? 2'h0 : state2; // @[Cache.scala 301:100 Cache.scala 301:109 Cache.scala 291:23]
  wire [28:0] hi_1 = io_in_bits_req_addr[31:3]; // @[Cache.scala 305:44]
  wire [31:0] raddr = {hi_1,3'h0}; // @[Cat.scala 30:58]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[Cat.scala 30:58]
  wire  _T_123 = state == 4'h1; // @[Cache.scala 309:23]
  wire [2:0] _T_125 = value_2 == 3'h7 ? 3'h7 : 3'h3; // @[Cache.scala 310:8]
  wire [2:0] cmd = state == 4'h1 ? 3'h2 : _T_125; // @[Cache.scala 309:16]
  wire  _T_131 = state2 == 2'h2; // @[Cache.scala 316:89]
  reg  afterFirstRead; // @[Cache.scala 323:31]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_12 = _T_70 | alreadyOutFire; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _T_137 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_139 = state == 4'h2; // @[Cache.scala 325:70]
  wire  readingFirst = ~afterFirstRead & _T_137 & state == 4'h2; // @[Cache.scala 325:60]
  wire  _T_142 = mmio ? state == 4'h6 : readingFirst; // @[Cache.scala 328:39]
  reg [63:0] inRdataRegDemand; // @[Reg.scala 27:20]
  wire  _T_143 = state == 4'h0; // @[Cache.scala 331:31]
  wire  _T_171 = 4'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_182 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_183 = io_mmio_req_ready & io_mmio_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_184 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire  _T_185 = io_mmio_resp_ready & io_mmio_resp_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_26 = _T_185 ? 4'h7 : state; // @[Cache.scala 360:50 Cache.scala 360:58 Cache.scala 281:22]
  wire  _T_186 = 4'h8 == state; // @[Conditional.scala 37:30]
  wire [2:0] _value_T_7 = value_1 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_27 = io_cohResp_valid ? _value_T_7 : value_1; // @[Cache.scala 363:48 Counter.scala 76:15 Counter.scala 60:40]
  wire  _T_195 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_29 = _T_118 ? 4'h2 : state; // @[Cache.scala 367:50 Cache.scala 368:13 Cache.scala 281:22]
  wire [2:0] _GEN_30 = _T_118 ? addr_wordIndex : value_1; // @[Cache.scala 367:50 Cache.scala 369:25 Counter.scala 60:40]
  wire  _T_197 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_201 = io_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [3:0] _GEN_32 = _T_201 ? 4'h7 : state; // @[Cache.scala 377:46 Cache.scala 377:54 Cache.scala 281:22]
  wire  _GEN_33 = _T_137 | afterFirstRead; // @[Cache.scala 373:33 Cache.scala 374:24 Cache.scala 323:31]
  wire [2:0] _GEN_34 = _T_137 ? _value_T_7 : value_1; // @[Cache.scala 373:33 Counter.scala 76:15 Counter.scala 60:40]
  wire [3:0] _GEN_36 = _T_137 ? _GEN_32 : state; // @[Cache.scala 373:33 Cache.scala 281:22]
  wire  _T_202 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _value_T_11 = value_2 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_37 = _T_118 ? _value_T_11 : value_2; // @[Cache.scala 382:32 Counter.scala 76:15 Counter.scala 60:40]
  wire  _T_205 = io_mem_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire [3:0] _GEN_38 = _T_205 & _T_118 ? 4'h4 : state; // @[Cache.scala 383:65 Cache.scala 383:73 Cache.scala 281:22]
  wire  _T_208 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_39 = _T_137 ? 4'h1 : state; // @[Cache.scala 386:53 Cache.scala 386:61 Cache.scala 281:22]
  wire  _T_210 = 4'h7 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_40 = _T_70 | needFlush | alreadyOutFire ? 4'h0 : state; // @[Cache.scala 387:76 Cache.scala 387:84 Cache.scala 281:22]
  wire [3:0] _GEN_41 = _T_210 ? _GEN_40 : state; // @[Conditional.scala 39:67 Cache.scala 281:22]
  wire [3:0] _GEN_42 = _T_208 ? _GEN_39 : _GEN_41; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_43 = _T_202 ? _GEN_37 : value_2; // @[Conditional.scala 39:67 Counter.scala 60:40]
  wire [3:0] _GEN_44 = _T_202 ? _GEN_38 : _GEN_42; // @[Conditional.scala 39:67]
  wire  _GEN_45 = _T_197 ? _GEN_33 : afterFirstRead; // @[Conditional.scala 39:67 Cache.scala 323:31]
  wire [2:0] _GEN_46 = _T_197 ? _GEN_34 : value_1; // @[Conditional.scala 39:67 Counter.scala 60:40]
  wire [3:0] _GEN_48 = _T_197 ? _GEN_36 : _GEN_44; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_49 = _T_197 ? value_2 : _GEN_43; // @[Conditional.scala 39:67 Counter.scala 60:40]
  wire [3:0] _GEN_50 = _T_195 ? _GEN_29 : _GEN_48; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_51 = _T_195 ? _GEN_30 : _GEN_46; // @[Conditional.scala 39:67]
  wire  _GEN_52 = _T_195 ? afterFirstRead : _GEN_45; // @[Conditional.scala 39:67 Cache.scala 323:31]
  wire [2:0] _GEN_54 = _T_195 ? value_2 : _GEN_49; // @[Conditional.scala 39:67 Counter.scala 60:40]
  wire [2:0] _GEN_55 = _T_186 ? _GEN_27 : _GEN_51; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_56 = _T_186 ? state : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_186 ? afterFirstRead : _GEN_52; // @[Conditional.scala 39:67 Cache.scala 323:31]
  wire [2:0] _GEN_59 = _T_186 ? value_2 : _GEN_54; // @[Conditional.scala 39:67 Counter.scala 60:40]
  wire  dataRefillWriteBus_req_valid = _T_139 & _T_137; // @[Cache.scala 392:39]
  wire  _T_247 = state == 4'h7; // @[Cache.scala 434:48]
  wire  _T_266 = mmio ? _T_247 : afterFirstRead & ~alreadyOutFire; // @[Cache.scala 435:45]
  wire  _T_267 = hit | _T_266; // @[Cache.scala 435:28]
  ysyx_210000_Arbiter metaWriteArb ( // @[Cache.scala 241:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_dirty(metaWriteArb_io_in_0_bits_data_dirty),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  ysyx_210000_Arbiter_1 dataWriteArb ( // @[Cache.scala 242:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = io_out_ready & _T_143 & ~miss; // @[Cache.scala 446:70]
  assign io_out_valid = io_in_valid & _T_267; // @[Cache.scala 433:31]
  assign io_out_bits_rdata = hit ? dataRead : inRdataRegDemand; // @[Cache.scala 427:29]
  assign io_out_bits_user = io_in_bits_req_user; // @[Cache.scala 430:56]
  assign io_isFinish = hit ? _T_70 : _T_247 & _GEN_12; // @[Cache.scala 443:8]
  assign io_dataReadBus_req_valid = (state == 4'h3 | state == 4'h8) & state2 == 2'h0; // @[Cache.scala 293:81]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,lo_2}; // @[Cat.scala 30:58]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[Cache.scala 397:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 397:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[Cache.scala 397:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[Cache.scala 397:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[Cache.scala 407:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 407:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 407:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 407:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[Cache.scala 407:23]
  assign io_mem_req_valid = _T_123 | _T_95 & state2 == 2'h2; // @[Cache.scala 316:48]
  assign io_mem_req_bits_addr = _T_123 ? raddr : waddr; // @[Cache.scala 311:35]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[Cache.scala 309:16]
  assign io_mem_req_bits_wdata = _T_112 | _T_110; // @[Mux.scala 27:72]
  assign io_mem_resp_ready = 1'h1; // @[Cache.scala 315:21]
  assign io_mmio_req_valid = state == 4'h5; // @[Cache.scala 321:31]
  assign io_mmio_req_bits_addr = io_in_bits_req_addr; // @[Cache.scala 319:20]
  assign io_mmio_req_bits_size = io_in_bits_req_size; // @[Cache.scala 319:20]
  assign io_mmio_resp_ready = 1'h1; // @[Cache.scala 320:22]
  assign io_cohResp_valid = _T_96 & _T_131; // @[Cache.scala 332:46]
  assign metaWriteArb_io_in_0_valid = 1'h0; // @[Cache.scala 276:22]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[9:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_0_bits_data_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  assign metaWriteArb_io_in_0_bits_data_dirty = 1'h0; // @[Cache.scala 277:16 Cache.scala 97:16]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 275:29 SRAMTemplate.scala 90:24]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_req_valid & _T_201; // @[Cache.scala 400:61]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[9:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:10]; // @[Cache.scala 245:31]
  assign metaWriteArb_io_in_1_bits_data_dirty = 1'h0; // @[Cache.scala 401:85]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 399:32 SRAMTemplate.scala 90:24]
  assign dataWriteArb_io_in_0_valid = 1'h0; // @[Cache.scala 270:22]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,addr_wordIndex}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_0_bits_data_data = useForwardData ? io_in_bits_forwardData_data_data : _T_49; // @[Cache.scala 262:21]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 271:29 SRAMTemplate.scala 90:24]
  assign dataWriteArb_io_in_1_valid = _T_139 & _T_137; // @[Cache.scala 392:39]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,value_1}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_1_bits_data_data = io_mem_resp_bits_rdata; // @[BitUtils.scala 32:25]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 391:32 SRAMTemplate.scala 90:24]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 281:22]
      state <= 4'h0; // @[Cache.scala 281:22]
    end else if (_T_171) begin // @[Conditional.scala 40:58]
      if ((miss | mmio) & ~io_flush) begin // @[Cache.scala 354:49]
        if (mmio) begin // @[Cache.scala 355:21]
          state <= 4'h5;
        end else begin
          state <= 4'h1;
        end
      end
    end else if (_T_182) begin // @[Conditional.scala 39:67]
      if (_T_183) begin // @[Cache.scala 359:48]
        state <= 4'h6; // @[Cache.scala 359:56]
      end
    end else if (_T_184) begin // @[Conditional.scala 39:67]
      state <= _GEN_26;
    end else begin
      state <= _GEN_56;
    end
    if (reset) begin // @[Cache.scala 282:26]
      needFlush <= 1'h0; // @[Cache.scala 282:26]
    end else if (_T_70 & needFlush) begin // @[Cache.scala 285:37]
      needFlush <= 1'h0; // @[Cache.scala 285:49]
    end else begin
      needFlush <= _GEN_1;
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 3'h0; // @[Counter.scala 60:40]
    end else if (!(_T_171)) begin // @[Conditional.scala 40:58]
      if (!(_T_182)) begin // @[Conditional.scala 39:67]
        if (!(_T_184)) begin // @[Conditional.scala 39:67]
          value_1 <= _GEN_55;
        end
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_2 <= 3'h0; // @[Counter.scala 60:40]
    end else if (!(_T_171)) begin // @[Conditional.scala 40:58]
      if (!(_T_182)) begin // @[Conditional.scala 39:67]
        if (!(_T_184)) begin // @[Conditional.scala 39:67]
          value_2 <= _GEN_59;
        end
      end
    end
    if (reset) begin // @[Cache.scala 291:23]
      state2 <= 2'h0; // @[Cache.scala 291:23]
    end else if (_T_114) begin // @[Conditional.scala 40:58]
      if (_T_115) begin // @[Cache.scala 299:53]
        state2 <= 2'h1; // @[Cache.scala 299:62]
      end
    end else if (_T_116) begin // @[Conditional.scala 39:67]
      state2 <= 2'h2; // @[Cache.scala 300:35]
    end else if (_T_117) begin // @[Conditional.scala 39:67]
      state2 <= _GEN_8;
    end
    if (reset) begin // @[Reg.scala 27:20]
      dataWay_0_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_102) begin // @[Reg.scala 28:19]
      dataWay_0_data <= io_dataReadBus_resp_data_0_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      dataWay_1_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_102) begin // @[Reg.scala 28:19]
      dataWay_1_data <= io_dataReadBus_resp_data_1_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      dataWay_2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_102) begin // @[Reg.scala 28:19]
      dataWay_2_data <= io_dataReadBus_resp_data_2_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      dataWay_3_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_102) begin // @[Reg.scala 28:19]
      dataWay_3_data <= io_dataReadBus_resp_data_3_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Cache.scala 323:31]
      afterFirstRead <= 1'h0; // @[Cache.scala 323:31]
    end else if (_T_171) begin // @[Conditional.scala 40:58]
      afterFirstRead <= 1'h0; // @[Cache.scala 343:22]
    end else if (!(_T_182)) begin // @[Conditional.scala 39:67]
      if (!(_T_184)) begin // @[Conditional.scala 39:67]
        afterFirstRead <= _GEN_57;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      alreadyOutFire <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_171) begin // @[Conditional.scala 40:58]
      alreadyOutFire <= 1'h0; // @[Cache.scala 344:22]
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (reset) begin // @[Reg.scala 27:20]
      inRdataRegDemand <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_142) begin // @[Reg.scala 28:19]
      if (mmio) begin // @[Cache.scala 326:39]
        inRdataRegDemand <= io_mmio_resp_bits_rdata;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:252 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"
            ); // @[Cache.scala 252:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fatal; // @[Cache.scala 252:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  needFlush = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_SRAMTemplate_1(
  input         clock,
  input         reset,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [3:0]  io_rreq_bits_setIdx,
  output [21:0] io_rresp_data_0_tag,
  output        io_rresp_data_0_valid,
  output        io_rresp_data_0_dirty,
  output [21:0] io_rresp_data_1_tag,
  output        io_rresp_data_1_valid,
  output        io_rresp_data_1_dirty,
  output [21:0] io_rresp_data_2_tag,
  output        io_rresp_data_2_valid,
  output        io_rresp_data_2_dirty,
  output [21:0] io_rresp_data_3_tag,
  output        io_rresp_data_3_valid,
  output        io_rresp_data_3_dirty,
  input         io_wreq_valid,
  input  [3:0]  io_wreq_bits_setIdx,
  input  [21:0] io_wreq_bits_data_tag,
  input         io_wreq_bits_data_dirty,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [3:0] array_RW0_addr; // @[SRAMTemplate.scala 128:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 128:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 128:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 128:26]
  wire [23:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 128:26]
  wire [23:0] array_RW0_wdata_1; // @[SRAMTemplate.scala 128:26]
  wire [23:0] array_RW0_wdata_2; // @[SRAMTemplate.scala 128:26]
  wire [23:0] array_RW0_wdata_3; // @[SRAMTemplate.scala 128:26]
  wire [23:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 128:26]
  wire [23:0] array_RW0_rdata_1; // @[SRAMTemplate.scala 128:26]
  wire [23:0] array_RW0_rdata_2; // @[SRAMTemplate.scala 128:26]
  wire [23:0] array_RW0_rdata_3; // @[SRAMTemplate.scala 128:26]
  wire  array_RW0_wmask_0; // @[SRAMTemplate.scala 128:26]
  wire  array_RW0_wmask_1; // @[SRAMTemplate.scala 128:26]
  wire  array_RW0_wmask_2; // @[SRAMTemplate.scala 128:26]
  wire  array_RW0_wmask_3; // @[SRAMTemplate.scala 128:26]
  reg  REG; // @[SRAMTemplate.scala 132:30]
  reg [3:0] REG_1; // @[Counter.scala 60:40]
  wire  _T = REG_1 == 4'hf; // @[Counter.scala 72:24]
  wire [3:0] _T_2 = REG_1 + 4'h1; // @[Counter.scala 76:24]
  wire  _GEN_1 = REG & _T; // @[Counter.scala 118:17 Counter.scala 118:24]
  wire  _GEN_2 = _GEN_1 ? 1'h0 : REG; // @[SRAMTemplate.scala 134:24 SRAMTemplate.scala 134:38 SRAMTemplate.scala 132:30]
  wire  wen = io_wreq_valid | REG; // @[SRAMTemplate.scala 140:52]
  wire  _T_3 = ~wen; // @[SRAMTemplate.scala 141:41]
  wire  realRen = io_rreq_valid & ~wen; // @[SRAMTemplate.scala 141:38]
  wire [3:0] setIdx = REG ? REG_1 : io_wreq_bits_setIdx; // @[SRAMTemplate.scala 143:19]
  wire [23:0] _T_4 = {io_wreq_bits_data_tag,1'h1,io_wreq_bits_data_dirty}; // @[SRAMTemplate.scala 144:78]
  wire [3:0] waymask = REG ? 4'hf : io_wreq_bits_waymask; // @[SRAMTemplate.scala 145:20]
  wire [23:0] _WIRE_3 = array_RW0_rdata_0;
  wire [23:0] _WIRE_4 = array_RW0_rdata_1;
  wire [23:0] _WIRE_5 = array_RW0_rdata_2;
  wire [23:0] _WIRE_6 = array_RW0_rdata_3;
  ysyx_210000_array_0 array ( // @[SRAMTemplate.scala 128:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_wdata_1(array_RW0_wdata_1),
    .RW0_wdata_2(array_RW0_wdata_2),
    .RW0_wdata_3(array_RW0_wdata_3),
    .RW0_rdata_0(array_RW0_rdata_0),
    .RW0_rdata_1(array_RW0_rdata_1),
    .RW0_rdata_2(array_RW0_rdata_2),
    .RW0_rdata_3(array_RW0_rdata_3),
    .RW0_wmask_0(array_RW0_wmask_0),
    .RW0_wmask_1(array_RW0_wmask_1),
    .RW0_wmask_2(array_RW0_wmask_2),
    .RW0_wmask_3(array_RW0_wmask_3)
  );
  assign io_rreq_ready = ~REG & _T_3; // @[SRAMTemplate.scala 153:33]
  assign io_rresp_data_0_tag = _WIRE_3[23:2]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_0_valid = _WIRE_3[1]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_0_dirty = _WIRE_3[0]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_1_tag = _WIRE_4[23:2]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_1_valid = _WIRE_4[1]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_1_dirty = _WIRE_4[0]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_2_tag = _WIRE_5[23:2]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_2_valid = _WIRE_5[1]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_2_dirty = _WIRE_5[0]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_3_tag = _WIRE_6[23:2]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_3_valid = _WIRE_6[1]; // @[SRAMTemplate.scala 150:78]
  assign io_rresp_data_3_dirty = _WIRE_6[0]; // @[SRAMTemplate.scala 150:78]
  assign array_RW0_wdata_0 = REG ? 24'h0 : _T_4; // @[SRAMTemplate.scala 144:22]
  assign array_RW0_wdata_1 = REG ? 24'h0 : _T_4; // @[SRAMTemplate.scala 144:22]
  assign array_RW0_wdata_2 = REG ? 24'h0 : _T_4; // @[SRAMTemplate.scala 144:22]
  assign array_RW0_wdata_3 = REG ? 24'h0 : _T_4; // @[SRAMTemplate.scala 144:22]
  assign array_RW0_wmask_0 = waymask[0]; // @[SRAMTemplate.scala 147:51]
  assign array_RW0_wmask_1 = waymask[1]; // @[SRAMTemplate.scala 147:51]
  assign array_RW0_wmask_2 = waymask[2]; // @[SRAMTemplate.scala 147:51]
  assign array_RW0_wmask_3 = waymask[3]; // @[SRAMTemplate.scala 147:51]
  assign array_RW0_wmode = io_wreq_valid | REG; // @[SRAMTemplate.scala 140:52]
  assign array_RW0_clk = clock;
  assign array_RW0_en = realRen | wen;
  assign array_RW0_addr = wen ? setIdx : io_rreq_bits_setIdx;
  always @(posedge clock) begin
    REG <= reset | _GEN_2; // @[SRAMTemplate.scala 132:30 SRAMTemplate.scala 132:30]
    if (reset) begin // @[Counter.scala 60:40]
      REG_1 <= 4'h0; // @[Counter.scala 60:40]
    end else if (REG) begin // @[Counter.scala 118:17]
      REG_1 <= _T_2; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_Arbiter_2(
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [3:0] io_in_0_bits_setIdx,
  input        io_out_ready,
  output       io_out_valid,
  output [3:0] io_out_bits_setIdx
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_bits_setIdx; // @[Arbiter.scala 124:15]
endmodule
module ysyx_210000_SRAMTemplateWithArbiter(
  input         clock,
  input         reset,
  output        io_r0_req_ready,
  input         io_r0_req_valid,
  input  [3:0]  io_r0_req_bits_setIdx,
  output [21:0] io_r0_resp_data_0_tag,
  output        io_r0_resp_data_0_valid,
  output        io_r0_resp_data_0_dirty,
  output [21:0] io_r0_resp_data_1_tag,
  output        io_r0_resp_data_1_valid,
  output        io_r0_resp_data_1_dirty,
  output [21:0] io_r0_resp_data_2_tag,
  output        io_r0_resp_data_2_valid,
  output        io_r0_resp_data_2_dirty,
  output [21:0] io_r0_resp_data_3_tag,
  output        io_r0_resp_data_3_valid,
  output        io_r0_resp_data_3_dirty,
  input         io_wreq_valid,
  input  [3:0]  io_wreq_bits_setIdx,
  input  [21:0] io_wreq_bits_data_tag,
  input         io_wreq_bits_data_dirty,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 351:24]
  wire  ram_reset; // @[SRAMTemplate.scala 351:24]
  wire  ram_io_rreq_ready; // @[SRAMTemplate.scala 351:24]
  wire  ram_io_rreq_valid; // @[SRAMTemplate.scala 351:24]
  wire [3:0] ram_io_rreq_bits_setIdx; // @[SRAMTemplate.scala 351:24]
  wire [21:0] ram_io_rresp_data_0_tag; // @[SRAMTemplate.scala 351:24]
  wire  ram_io_rresp_data_0_valid; // @[SRAMTemplate.scala 351:24]
  wire  ram_io_rresp_data_0_dirty; // @[SRAMTemplate.scala 351:24]
  wire [21:0] ram_io_rresp_data_1_tag; // @[SRAMTemplate.scala 351:24]
  wire  ram_io_rresp_data_1_valid; // @[SRAMTemplate.scala 351:24]
  wire  ram_io_rresp_data_1_dirty; // @[SRAMTemplate.scala 351:24]
  wire [21:0] ram_io_rresp_data_2_tag; // @[SRAMTemplate.scala 351:24]
  wire  ram_io_rresp_data_2_valid; // @[SRAMTemplate.scala 351:24]
  wire  ram_io_rresp_data_2_dirty; // @[SRAMTemplate.scala 351:24]
  wire [21:0] ram_io_rresp_data_3_tag; // @[SRAMTemplate.scala 351:24]
  wire  ram_io_rresp_data_3_valid; // @[SRAMTemplate.scala 351:24]
  wire  ram_io_rresp_data_3_dirty; // @[SRAMTemplate.scala 351:24]
  wire  ram_io_wreq_valid; // @[SRAMTemplate.scala 351:24]
  wire [3:0] ram_io_wreq_bits_setIdx; // @[SRAMTemplate.scala 351:24]
  wire [21:0] ram_io_wreq_bits_data_tag; // @[SRAMTemplate.scala 351:24]
  wire  ram_io_wreq_bits_data_dirty; // @[SRAMTemplate.scala 351:24]
  wire [3:0] ram_io_wreq_bits_waymask; // @[SRAMTemplate.scala 351:24]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 355:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 355:23]
  wire [3:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 355:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 355:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 355:23]
  wire [3:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 355:23]
  wire  _T = io_r0_req_ready & io_r0_req_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[SRAMTemplate.scala 361:58]
  reg [21:0] REG_1_0_tag; // @[Reg.scala 27:20]
  reg  REG_1_0_valid; // @[Reg.scala 27:20]
  reg  REG_1_0_dirty; // @[Reg.scala 27:20]
  reg [21:0] REG_1_1_tag; // @[Reg.scala 27:20]
  reg  REG_1_1_valid; // @[Reg.scala 27:20]
  reg  REG_1_1_dirty; // @[Reg.scala 27:20]
  reg [21:0] REG_1_2_tag; // @[Reg.scala 27:20]
  reg  REG_1_2_valid; // @[Reg.scala 27:20]
  reg  REG_1_2_dirty; // @[Reg.scala 27:20]
  reg [21:0] REG_1_3_tag; // @[Reg.scala 27:20]
  reg  REG_1_3_valid; // @[Reg.scala 27:20]
  reg  REG_1_3_dirty; // @[Reg.scala 27:20]
  ysyx_210000_SRAMTemplate_1 ram ( // @[SRAMTemplate.scala 351:24]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_rreq_ready(ram_io_rreq_ready),
    .io_rreq_valid(ram_io_rreq_valid),
    .io_rreq_bits_setIdx(ram_io_rreq_bits_setIdx),
    .io_rresp_data_0_tag(ram_io_rresp_data_0_tag),
    .io_rresp_data_0_valid(ram_io_rresp_data_0_valid),
    .io_rresp_data_0_dirty(ram_io_rresp_data_0_dirty),
    .io_rresp_data_1_tag(ram_io_rresp_data_1_tag),
    .io_rresp_data_1_valid(ram_io_rresp_data_1_valid),
    .io_rresp_data_1_dirty(ram_io_rresp_data_1_dirty),
    .io_rresp_data_2_tag(ram_io_rresp_data_2_tag),
    .io_rresp_data_2_valid(ram_io_rresp_data_2_valid),
    .io_rresp_data_2_dirty(ram_io_rresp_data_2_dirty),
    .io_rresp_data_3_tag(ram_io_rresp_data_3_tag),
    .io_rresp_data_3_valid(ram_io_rresp_data_3_valid),
    .io_rresp_data_3_dirty(ram_io_rresp_data_3_dirty),
    .io_wreq_valid(ram_io_wreq_valid),
    .io_wreq_bits_setIdx(ram_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(ram_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(ram_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(ram_io_wreq_bits_waymask)
  );
  ysyx_210000_Arbiter_2 readArb ( // @[SRAMTemplate.scala 355:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 356:17]
  assign io_r0_resp_data_0_tag = REG ? ram_io_rresp_data_0_tag : REG_1_0_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_0_valid = REG ? ram_io_rresp_data_0_valid : REG_1_0_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_0_dirty = REG ? ram_io_rresp_data_0_dirty : REG_1_0_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_tag = REG ? ram_io_rresp_data_1_tag : REG_1_1_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_valid = REG ? ram_io_rresp_data_1_valid : REG_1_1_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_dirty = REG ? ram_io_rresp_data_1_dirty : REG_1_1_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_tag = REG ? ram_io_rresp_data_2_tag : REG_1_2_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_valid = REG ? ram_io_rresp_data_2_valid : REG_1_2_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_dirty = REG ? ram_io_rresp_data_2_dirty : REG_1_2_dirty; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_tag = REG ? ram_io_rresp_data_3_tag : REG_1_3_tag; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_valid = REG ? ram_io_rresp_data_3_valid : REG_1_3_valid; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_dirty = REG ? ram_io_rresp_data_3_dirty : REG_1_3_dirty; // @[Hold.scala 23:48]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_rreq_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 357:16]
  assign ram_io_rreq_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 357:16]
  assign ram_io_wreq_valid = io_wreq_valid; // @[SRAMTemplate.scala 353:12]
  assign ram_io_wreq_bits_setIdx = io_wreq_bits_setIdx; // @[SRAMTemplate.scala 353:12]
  assign ram_io_wreq_bits_data_tag = io_wreq_bits_data_tag; // @[SRAMTemplate.scala 353:12]
  assign ram_io_wreq_bits_data_dirty = io_wreq_bits_data_dirty; // @[SRAMTemplate.scala 353:12]
  assign ram_io_wreq_bits_waymask = io_wreq_bits_waymask; // @[SRAMTemplate.scala 353:12]
  assign readArb_io_in_0_valid = io_r0_req_valid; // @[SRAMTemplate.scala 356:17]
  assign readArb_io_in_0_bits_setIdx = io_r0_req_bits_setIdx; // @[SRAMTemplate.scala 356:17]
  assign readArb_io_out_ready = ram_io_rreq_ready; // @[SRAMTemplate.scala 357:16]
  always @(posedge clock) begin
    if (reset) begin // @[SRAMTemplate.scala 361:58]
      REG <= 1'h0; // @[SRAMTemplate.scala 361:58]
    end else begin
      REG <= _T; // @[SRAMTemplate.scala 361:58]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_0_tag <= 22'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_0_tag <= ram_io_rresp_data_0_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_0_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_0_valid <= ram_io_rresp_data_0_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_0_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_0_dirty <= ram_io_rresp_data_0_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_1_tag <= 22'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_1_tag <= ram_io_rresp_data_1_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_1_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_1_valid <= ram_io_rresp_data_1_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_1_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_1_dirty <= ram_io_rresp_data_1_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_2_tag <= 22'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_2_tag <= ram_io_rresp_data_2_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_2_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_2_valid <= ram_io_rresp_data_2_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_2_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_2_dirty <= ram_io_rresp_data_2_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_3_tag <= 22'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_3_tag <= ram_io_rresp_data_3_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_3_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_3_valid <= ram_io_rresp_data_3_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_3_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_3_dirty <= ram_io_rresp_data_3_dirty; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1_0_tag = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  REG_1_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  REG_1_0_dirty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_1_1_tag = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1_1_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  REG_1_1_dirty = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  REG_1_2_tag = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  REG_1_2_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  REG_1_2_dirty = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  REG_1_3_tag = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  REG_1_3_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  REG_1_3_dirty = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_SRAMWrapper(
  input          clock,
  input          reset,
  output [127:0] io_Q,
  input          io_CLK,
  input          io_CEN,
  input          io_WEN,
  input  [127:0] io_BWEN,
  input  [6:0]   io_A,
  input  [127:0] io_D
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [127:0] sram_lo_Q; // @[SRAMTemplate.scala 55:23]
  wire  sram_lo_CLK; // @[SRAMTemplate.scala 55:23]
  wire  sram_lo_CEN; // @[SRAMTemplate.scala 55:23]
  wire  sram_lo_WEN; // @[SRAMTemplate.scala 55:23]
  wire [127:0] sram_lo_BWEN; // @[SRAMTemplate.scala 55:23]
  wire [5:0] sram_lo_A; // @[SRAMTemplate.scala 55:23]
  wire [127:0] sram_lo_D; // @[SRAMTemplate.scala 55:23]
  wire [127:0] sram_hi_Q; // @[SRAMTemplate.scala 56:23]
  wire  sram_hi_CLK; // @[SRAMTemplate.scala 56:23]
  wire  sram_hi_CEN; // @[SRAMTemplate.scala 56:23]
  wire  sram_hi_WEN; // @[SRAMTemplate.scala 56:23]
  wire [127:0] sram_hi_BWEN; // @[SRAMTemplate.scala 56:23]
  wire [5:0] sram_hi_A; // @[SRAMTemplate.scala 56:23]
  wire [127:0] sram_hi_D; // @[SRAMTemplate.scala 56:23]
  reg  REG; // @[SRAMTemplate.scala 71:22]
  S011HD1P_X32Y2D128_BW sram_lo ( // @[SRAMTemplate.scala 55:23]
    .Q(sram_lo_Q),
    .CLK(sram_lo_CLK),
    .CEN(sram_lo_CEN),
    .WEN(sram_lo_WEN),
    .BWEN(sram_lo_BWEN),
    .A(sram_lo_A),
    .D(sram_lo_D)
  );
  S011HD1P_X32Y2D128_BW sram_hi ( // @[SRAMTemplate.scala 56:23]
    .Q(sram_hi_Q),
    .CLK(sram_hi_CLK),
    .CEN(sram_hi_CEN),
    .WEN(sram_hi_WEN),
    .BWEN(sram_hi_BWEN),
    .A(sram_hi_A),
    .D(sram_hi_D)
  );
  assign io_Q = REG ? sram_hi_Q : sram_lo_Q; // @[SRAMTemplate.scala 71:14]
  assign sram_lo_CLK = io_CLK; // @[SRAMTemplate.scala 57:18]
  assign sram_lo_CEN = io_A[6] | io_CEN; // @[SRAMTemplate.scala 58:29]
  assign sram_lo_WEN = io_WEN; // @[SRAMTemplate.scala 59:18]
  assign sram_lo_BWEN = io_BWEN; // @[SRAMTemplate.scala 60:19]
  assign sram_lo_A = io_A[5:0]; // @[SRAMTemplate.scala 61:23]
  assign sram_lo_D = io_D; // @[SRAMTemplate.scala 62:16]
  assign sram_hi_CLK = io_CLK; // @[SRAMTemplate.scala 64:18]
  assign sram_hi_CEN = ~io_A[6] | io_CEN; // @[SRAMTemplate.scala 65:30]
  assign sram_hi_WEN = io_WEN; // @[SRAMTemplate.scala 66:18]
  assign sram_hi_BWEN = io_BWEN; // @[SRAMTemplate.scala 67:19]
  assign sram_hi_A = io_A[5:0]; // @[SRAMTemplate.scala 68:23]
  assign sram_hi_D = io_D; // @[SRAMTemplate.scala 69:16]
  always @(posedge clock) begin
    if (reset) begin // @[SRAMTemplate.scala 71:22]
      REG <= 1'h0; // @[SRAMTemplate.scala 71:22]
    end else begin
      REG <= io_A[6]; // @[SRAMTemplate.scala 71:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_DataSRAMTemplate(
  input         clock,
  input         reset,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [6:0]  io_rreq_bits_setIdx,
  output [63:0] io_rresp_data_0_data,
  output [63:0] io_rresp_data_1_data,
  output [63:0] io_rresp_data_2_data,
  output [63:0] io_rresp_data_3_data,
  input         io_wreq_valid,
  input  [6:0]  io_wreq_bits_setIdx,
  input  [63:0] io_wreq_bits_data_data,
  input  [3:0]  io_wreq_bits_waymask
);
  wire  sram_0_clock; // @[SRAMTemplate.scala 288:32]
  wire  sram_0_reset; // @[SRAMTemplate.scala 288:32]
  wire [127:0] sram_0_io_Q; // @[SRAMTemplate.scala 288:32]
  wire  sram_0_io_CLK; // @[SRAMTemplate.scala 288:32]
  wire  sram_0_io_CEN; // @[SRAMTemplate.scala 288:32]
  wire  sram_0_io_WEN; // @[SRAMTemplate.scala 288:32]
  wire [127:0] sram_0_io_BWEN; // @[SRAMTemplate.scala 288:32]
  wire [6:0] sram_0_io_A; // @[SRAMTemplate.scala 288:32]
  wire [127:0] sram_0_io_D; // @[SRAMTemplate.scala 288:32]
  wire  sram_1_clock; // @[SRAMTemplate.scala 288:32]
  wire  sram_1_reset; // @[SRAMTemplate.scala 288:32]
  wire [127:0] sram_1_io_Q; // @[SRAMTemplate.scala 288:32]
  wire  sram_1_io_CLK; // @[SRAMTemplate.scala 288:32]
  wire  sram_1_io_CEN; // @[SRAMTemplate.scala 288:32]
  wire  sram_1_io_WEN; // @[SRAMTemplate.scala 288:32]
  wire [127:0] sram_1_io_BWEN; // @[SRAMTemplate.scala 288:32]
  wire [6:0] sram_1_io_A; // @[SRAMTemplate.scala 288:32]
  wire [127:0] sram_1_io_D; // @[SRAMTemplate.scala 288:32]
  wire  realRen = io_rreq_valid & ~io_wreq_valid; // @[SRAMTemplate.scala 301:38]
  wire  hi = |io_wreq_bits_waymask[3:2]; // @[OneHot.scala 32:14]
  wire [1:0] _T_10 = io_wreq_bits_waymask[3:2] | io_wreq_bits_waymask[1:0]; // @[OneHot.scala 32:28]
  wire  lo = _T_10[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] _T_11 = {hi,lo}; // @[Cat.scala 30:58]
  wire [63:0] lo_2 = _T_10[0] ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] hi_2 = lo ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [127:0] _T_31 = {hi_2,lo_2}; // @[Cat.scala 30:58]
  wire [255:0] _T_44 = {sram_1_io_Q,sram_0_io_Q}; // @[Cat.scala 30:58]
  ysyx_210000_SRAMWrapper sram_0 ( // @[SRAMTemplate.scala 288:32]
    .clock(sram_0_clock),
    .reset(sram_0_reset),
    .io_Q(sram_0_io_Q),
    .io_CLK(sram_0_io_CLK),
    .io_CEN(sram_0_io_CEN),
    .io_WEN(sram_0_io_WEN),
    .io_BWEN(sram_0_io_BWEN),
    .io_A(sram_0_io_A),
    .io_D(sram_0_io_D)
  );
  ysyx_210000_SRAMWrapper sram_1 ( // @[SRAMTemplate.scala 288:32]
    .clock(sram_1_clock),
    .reset(sram_1_reset),
    .io_Q(sram_1_io_Q),
    .io_CLK(sram_1_io_CLK),
    .io_CEN(sram_1_io_CEN),
    .io_WEN(sram_1_io_WEN),
    .io_BWEN(sram_1_io_BWEN),
    .io_A(sram_1_io_A),
    .io_D(sram_1_io_D)
  );
  assign io_rreq_ready = ~io_wreq_valid; // @[SRAMTemplate.scala 325:53]
  assign io_rresp_data_0_data = _T_44[63:0]; // @[SRAMTemplate.scala 322:53]
  assign io_rresp_data_1_data = _T_44[127:64]; // @[SRAMTemplate.scala 322:53]
  assign io_rresp_data_2_data = _T_44[191:128]; // @[SRAMTemplate.scala 322:53]
  assign io_rresp_data_3_data = _T_44[255:192]; // @[SRAMTemplate.scala 322:53]
  assign sram_0_clock = clock;
  assign sram_0_reset = reset;
  assign sram_0_io_CLK = clock; // @[SRAMTemplate.scala 309:21]
  assign sram_0_io_CEN = ~(io_wreq_valid | realRen); // @[SRAMTemplate.scala 312:32]
  assign sram_0_io_WEN = ~(io_wreq_valid & ~_T_11[1]); // @[SRAMTemplate.scala 315:32]
  assign sram_0_io_BWEN = ~_T_31; // @[SRAMTemplate.scala 318:33]
  assign sram_0_io_A = io_wreq_valid ? io_wreq_bits_setIdx : io_rreq_bits_setIdx; // @[SRAMTemplate.scala 310:25]
  assign sram_0_io_D = {io_wreq_bits_data_data,io_wreq_bits_data_data}; // @[Cat.scala 30:58]
  assign sram_1_clock = clock;
  assign sram_1_reset = reset;
  assign sram_1_io_CLK = clock; // @[SRAMTemplate.scala 309:21]
  assign sram_1_io_CEN = ~(io_wreq_valid | realRen); // @[SRAMTemplate.scala 312:32]
  assign sram_1_io_WEN = ~(io_wreq_valid & _T_11[1]); // @[SRAMTemplate.scala 315:32]
  assign sram_1_io_BWEN = ~_T_31; // @[SRAMTemplate.scala 318:33]
  assign sram_1_io_A = io_wreq_valid ? io_wreq_bits_setIdx : io_rreq_bits_setIdx; // @[SRAMTemplate.scala 310:25]
  assign sram_1_io_D = {io_wreq_bits_data_data,io_wreq_bits_data_data}; // @[Cat.scala 30:58]
endmodule
module ysyx_210000_Arbiter_3(
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [6:0] io_in_0_bits_setIdx,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input  [6:0] io_in_1_bits_setIdx,
  input        io_out_ready,
  output       io_out_valid,
  output [6:0] io_out_bits_setIdx
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
endmodule
module ysyx_210000_SRAMTemplateWithArbiter_1(
  input         clock,
  input         reset,
  output        io_r0_req_ready,
  input         io_r0_req_valid,
  input  [6:0]  io_r0_req_bits_setIdx,
  output [63:0] io_r0_resp_data_0_data,
  output [63:0] io_r0_resp_data_1_data,
  output [63:0] io_r0_resp_data_2_data,
  output [63:0] io_r0_resp_data_3_data,
  output        io_r1_req_ready,
  input         io_r1_req_valid,
  input  [6:0]  io_r1_req_bits_setIdx,
  output [63:0] io_r1_resp_data_0_data,
  output [63:0] io_r1_resp_data_1_data,
  output [63:0] io_r1_resp_data_2_data,
  output [63:0] io_r1_resp_data_3_data,
  input         io_wreq_valid,
  input  [6:0]  io_wreq_bits_setIdx,
  input  [63:0] io_wreq_bits_data_data,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 350:31]
  wire  ram_reset; // @[SRAMTemplate.scala 350:31]
  wire  ram_io_rreq_ready; // @[SRAMTemplate.scala 350:31]
  wire  ram_io_rreq_valid; // @[SRAMTemplate.scala 350:31]
  wire [6:0] ram_io_rreq_bits_setIdx; // @[SRAMTemplate.scala 350:31]
  wire [63:0] ram_io_rresp_data_0_data; // @[SRAMTemplate.scala 350:31]
  wire [63:0] ram_io_rresp_data_1_data; // @[SRAMTemplate.scala 350:31]
  wire [63:0] ram_io_rresp_data_2_data; // @[SRAMTemplate.scala 350:31]
  wire [63:0] ram_io_rresp_data_3_data; // @[SRAMTemplate.scala 350:31]
  wire  ram_io_wreq_valid; // @[SRAMTemplate.scala 350:31]
  wire [6:0] ram_io_wreq_bits_setIdx; // @[SRAMTemplate.scala 350:31]
  wire [63:0] ram_io_wreq_bits_data_data; // @[SRAMTemplate.scala 350:31]
  wire [3:0] ram_io_wreq_bits_waymask; // @[SRAMTemplate.scala 350:31]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 355:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 355:23]
  wire [6:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 355:23]
  wire  readArb_io_in_1_ready; // @[SRAMTemplate.scala 355:23]
  wire  readArb_io_in_1_valid; // @[SRAMTemplate.scala 355:23]
  wire [6:0] readArb_io_in_1_bits_setIdx; // @[SRAMTemplate.scala 355:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 355:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 355:23]
  wire [6:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 355:23]
  wire  _T = io_r0_req_ready & io_r0_req_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[SRAMTemplate.scala 361:58]
  reg [63:0] REG_1_0_data; // @[Reg.scala 27:20]
  reg [63:0] REG_1_1_data; // @[Reg.scala 27:20]
  reg [63:0] REG_1_2_data; // @[Reg.scala 27:20]
  reg [63:0] REG_1_3_data; // @[Reg.scala 27:20]
  wire  _T_2 = io_r1_req_ready & io_r1_req_valid; // @[Decoupled.scala 40:37]
  reg  REG_2; // @[SRAMTemplate.scala 361:58]
  reg [63:0] REG_3_0_data; // @[Reg.scala 27:20]
  reg [63:0] REG_3_1_data; // @[Reg.scala 27:20]
  reg [63:0] REG_3_2_data; // @[Reg.scala 27:20]
  reg [63:0] REG_3_3_data; // @[Reg.scala 27:20]
  ysyx_210000_DataSRAMTemplate ram ( // @[SRAMTemplate.scala 350:31]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_rreq_ready(ram_io_rreq_ready),
    .io_rreq_valid(ram_io_rreq_valid),
    .io_rreq_bits_setIdx(ram_io_rreq_bits_setIdx),
    .io_rresp_data_0_data(ram_io_rresp_data_0_data),
    .io_rresp_data_1_data(ram_io_rresp_data_1_data),
    .io_rresp_data_2_data(ram_io_rresp_data_2_data),
    .io_rresp_data_3_data(ram_io_rresp_data_3_data),
    .io_wreq_valid(ram_io_wreq_valid),
    .io_wreq_bits_setIdx(ram_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(ram_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(ram_io_wreq_bits_waymask)
  );
  ysyx_210000_Arbiter_3 readArb ( // @[SRAMTemplate.scala 355:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_in_1_ready(readArb_io_in_1_ready),
    .io_in_1_valid(readArb_io_in_1_valid),
    .io_in_1_bits_setIdx(readArb_io_in_1_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 356:17]
  assign io_r0_resp_data_0_data = REG ? ram_io_rresp_data_0_data : REG_1_0_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_1_data = REG ? ram_io_rresp_data_1_data : REG_1_1_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_2_data = REG ? ram_io_rresp_data_2_data : REG_1_2_data; // @[Hold.scala 23:48]
  assign io_r0_resp_data_3_data = REG ? ram_io_rresp_data_3_data : REG_1_3_data; // @[Hold.scala 23:48]
  assign io_r1_req_ready = readArb_io_in_1_ready; // @[SRAMTemplate.scala 356:17]
  assign io_r1_resp_data_0_data = REG_2 ? ram_io_rresp_data_0_data : REG_3_0_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_1_data = REG_2 ? ram_io_rresp_data_1_data : REG_3_1_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_2_data = REG_2 ? ram_io_rresp_data_2_data : REG_3_2_data; // @[Hold.scala 23:48]
  assign io_r1_resp_data_3_data = REG_2 ? ram_io_rresp_data_3_data : REG_3_3_data; // @[Hold.scala 23:48]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_rreq_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 357:16]
  assign ram_io_rreq_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 357:16]
  assign ram_io_wreq_valid = io_wreq_valid; // @[SRAMTemplate.scala 353:12]
  assign ram_io_wreq_bits_setIdx = io_wreq_bits_setIdx; // @[SRAMTemplate.scala 353:12]
  assign ram_io_wreq_bits_data_data = io_wreq_bits_data_data; // @[SRAMTemplate.scala 353:12]
  assign ram_io_wreq_bits_waymask = io_wreq_bits_waymask; // @[SRAMTemplate.scala 353:12]
  assign readArb_io_in_0_valid = io_r0_req_valid; // @[SRAMTemplate.scala 356:17]
  assign readArb_io_in_0_bits_setIdx = io_r0_req_bits_setIdx; // @[SRAMTemplate.scala 356:17]
  assign readArb_io_in_1_valid = io_r1_req_valid; // @[SRAMTemplate.scala 356:17]
  assign readArb_io_in_1_bits_setIdx = io_r1_req_bits_setIdx; // @[SRAMTemplate.scala 356:17]
  assign readArb_io_out_ready = ram_io_rreq_ready; // @[SRAMTemplate.scala 357:16]
  always @(posedge clock) begin
    if (reset) begin // @[SRAMTemplate.scala 361:58]
      REG <= 1'h0; // @[SRAMTemplate.scala 361:58]
    end else begin
      REG <= _T; // @[SRAMTemplate.scala 361:58]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_0_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_0_data <= ram_io_rresp_data_0_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_1_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_1_data <= ram_io_rresp_data_1_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_2_data <= ram_io_rresp_data_2_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_3_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG) begin // @[Reg.scala 28:19]
      REG_1_3_data <= ram_io_rresp_data_3_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[SRAMTemplate.scala 361:58]
      REG_2 <= 1'h0; // @[SRAMTemplate.scala 361:58]
    end else begin
      REG_2 <= _T_2; // @[SRAMTemplate.scala 361:58]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_0_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_2) begin // @[Reg.scala 28:19]
      REG_3_0_data <= ram_io_rresp_data_0_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_1_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_2) begin // @[Reg.scala 28:19]
      REG_3_1_data <= ram_io_rresp_data_1_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_2) begin // @[Reg.scala 28:19]
      REG_3_2_data <= ram_io_rresp_data_2_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_3_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (REG_2) begin // @[Reg.scala 28:19]
      REG_3_3_data <= ram_io_rresp_data_3_data; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  REG_1_0_data = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  REG_1_1_data = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  REG_1_2_data = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  REG_1_3_data = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  REG_2 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  REG_3_0_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  REG_3_1_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  REG_3_2_data = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  REG_3_3_data = _RAND_9[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_Arbiter_4(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [2:0]  io_in_0_bits_size,
  input  [86:0] io_in_0_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [86:0] io_out_bits_user
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_addr = io_in_0_bits_addr; // @[Arbiter.scala 124:15]
  assign io_out_bits_size = io_in_0_bits_size; // @[Arbiter.scala 124:15]
  assign io_out_bits_user = io_in_0_bits_user; // @[Arbiter.scala 124:15]
endmodule
module ysyx_210000_Cache(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [86:0] io_in_req_bits_user,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output [86:0] io_in_resp_bits_user,
  input  [1:0]  io_flush,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_empty,
  input         MOUFlushICache
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [95:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire  s1_io_in_ready; // @[Cache.scala 476:18]
  wire  s1_io_in_valid; // @[Cache.scala 476:18]
  wire [31:0] s1_io_in_bits_addr; // @[Cache.scala 476:18]
  wire [2:0] s1_io_in_bits_size; // @[Cache.scala 476:18]
  wire [86:0] s1_io_in_bits_user; // @[Cache.scala 476:18]
  wire  s1_io_out_ready; // @[Cache.scala 476:18]
  wire  s1_io_out_valid; // @[Cache.scala 476:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[Cache.scala 476:18]
  wire [2:0] s1_io_out_bits_req_size; // @[Cache.scala 476:18]
  wire [86:0] s1_io_out_bits_req_user; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_req_ready; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_req_valid; // @[Cache.scala 476:18]
  wire [3:0] s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [21:0] s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 476:18]
  wire [21:0] s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 476:18]
  wire [21:0] s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 476:18]
  wire [21:0] s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 476:18]
  wire  s1_io_dataReadBus_req_ready; // @[Cache.scala 476:18]
  wire  s1_io_dataReadBus_req_valid; // @[Cache.scala 476:18]
  wire [6:0] s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 476:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 476:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 476:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 476:18]
  wire  s2_clock; // @[Cache.scala 477:18]
  wire  s2_reset; // @[Cache.scala 477:18]
  wire  s2_io_in_ready; // @[Cache.scala 477:18]
  wire  s2_io_in_valid; // @[Cache.scala 477:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[Cache.scala 477:18]
  wire [2:0] s2_io_in_bits_req_size; // @[Cache.scala 477:18]
  wire [86:0] s2_io_in_bits_req_user; // @[Cache.scala 477:18]
  wire  s2_io_out_ready; // @[Cache.scala 477:18]
  wire  s2_io_out_valid; // @[Cache.scala 477:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[Cache.scala 477:18]
  wire [2:0] s2_io_out_bits_req_size; // @[Cache.scala 477:18]
  wire [86:0] s2_io_out_bits_req_user; // @[Cache.scala 477:18]
  wire [21:0] s2_io_out_bits_metas_0_tag; // @[Cache.scala 477:18]
  wire [21:0] s2_io_out_bits_metas_1_tag; // @[Cache.scala 477:18]
  wire [21:0] s2_io_out_bits_metas_2_tag; // @[Cache.scala 477:18]
  wire [21:0] s2_io_out_bits_metas_3_tag; // @[Cache.scala 477:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[Cache.scala 477:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[Cache.scala 477:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[Cache.scala 477:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[Cache.scala 477:18]
  wire  s2_io_out_bits_hit; // @[Cache.scala 477:18]
  wire [3:0] s2_io_out_bits_waymask; // @[Cache.scala 477:18]
  wire  s2_io_out_bits_mmio; // @[Cache.scala 477:18]
  wire  s2_io_out_bits_isForwardData; // @[Cache.scala 477:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[Cache.scala 477:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[Cache.scala 477:18]
  wire [21:0] s2_io_metaReadResp_0_tag; // @[Cache.scala 477:18]
  wire  s2_io_metaReadResp_0_valid; // @[Cache.scala 477:18]
  wire [21:0] s2_io_metaReadResp_1_tag; // @[Cache.scala 477:18]
  wire  s2_io_metaReadResp_1_valid; // @[Cache.scala 477:18]
  wire [21:0] s2_io_metaReadResp_2_tag; // @[Cache.scala 477:18]
  wire  s2_io_metaReadResp_2_valid; // @[Cache.scala 477:18]
  wire [21:0] s2_io_metaReadResp_3_tag; // @[Cache.scala 477:18]
  wire  s2_io_metaReadResp_3_valid; // @[Cache.scala 477:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[Cache.scala 477:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[Cache.scala 477:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[Cache.scala 477:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[Cache.scala 477:18]
  wire  s2_io_metaWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [21:0] s2_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 477:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s2_io_dataWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [6:0] s2_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 477:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_clock; // @[Cache.scala 478:18]
  wire  s3_reset; // @[Cache.scala 478:18]
  wire  s3_io_in_ready; // @[Cache.scala 478:18]
  wire  s3_io_in_valid; // @[Cache.scala 478:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[Cache.scala 478:18]
  wire [2:0] s3_io_in_bits_req_size; // @[Cache.scala 478:18]
  wire [86:0] s3_io_in_bits_req_user; // @[Cache.scala 478:18]
  wire [21:0] s3_io_in_bits_metas_0_tag; // @[Cache.scala 478:18]
  wire [21:0] s3_io_in_bits_metas_1_tag; // @[Cache.scala 478:18]
  wire [21:0] s3_io_in_bits_metas_2_tag; // @[Cache.scala 478:18]
  wire [21:0] s3_io_in_bits_metas_3_tag; // @[Cache.scala 478:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[Cache.scala 478:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[Cache.scala 478:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[Cache.scala 478:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[Cache.scala 478:18]
  wire  s3_io_in_bits_hit; // @[Cache.scala 478:18]
  wire [3:0] s3_io_in_bits_waymask; // @[Cache.scala 478:18]
  wire  s3_io_in_bits_mmio; // @[Cache.scala 478:18]
  wire  s3_io_in_bits_isForwardData; // @[Cache.scala 478:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[Cache.scala 478:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[Cache.scala 478:18]
  wire  s3_io_out_ready; // @[Cache.scala 478:18]
  wire  s3_io_out_valid; // @[Cache.scala 478:18]
  wire [63:0] s3_io_out_bits_rdata; // @[Cache.scala 478:18]
  wire [86:0] s3_io_out_bits_user; // @[Cache.scala 478:18]
  wire  s3_io_isFinish; // @[Cache.scala 478:18]
  wire  s3_io_flush; // @[Cache.scala 478:18]
  wire  s3_io_dataReadBus_req_ready; // @[Cache.scala 478:18]
  wire  s3_io_dataReadBus_req_valid; // @[Cache.scala 478:18]
  wire [6:0] s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 478:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[Cache.scala 478:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[Cache.scala 478:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[Cache.scala 478:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[Cache.scala 478:18]
  wire  s3_io_dataWriteBus_req_valid; // @[Cache.scala 478:18]
  wire [6:0] s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 478:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 478:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 478:18]
  wire  s3_io_metaWriteBus_req_valid; // @[Cache.scala 478:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 478:18]
  wire [21:0] s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 478:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 478:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 478:18]
  wire  s3_io_mem_req_ready; // @[Cache.scala 478:18]
  wire  s3_io_mem_req_valid; // @[Cache.scala 478:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[Cache.scala 478:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[Cache.scala 478:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[Cache.scala 478:18]
  wire  s3_io_mem_resp_ready; // @[Cache.scala 478:18]
  wire  s3_io_mem_resp_valid; // @[Cache.scala 478:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[Cache.scala 478:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[Cache.scala 478:18]
  wire  s3_io_mmio_req_ready; // @[Cache.scala 478:18]
  wire  s3_io_mmio_req_valid; // @[Cache.scala 478:18]
  wire [31:0] s3_io_mmio_req_bits_addr; // @[Cache.scala 478:18]
  wire [2:0] s3_io_mmio_req_bits_size; // @[Cache.scala 478:18]
  wire  s3_io_mmio_resp_ready; // @[Cache.scala 478:18]
  wire  s3_io_mmio_resp_valid; // @[Cache.scala 478:18]
  wire [63:0] s3_io_mmio_resp_bits_rdata; // @[Cache.scala 478:18]
  wire  s3_io_cohResp_valid; // @[Cache.scala 478:18]
  wire  metaArray_clock; // @[Cache.scala 479:25]
  wire  metaArray_reset; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_req_ready; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_req_valid; // @[Cache.scala 479:25]
  wire [3:0] metaArray_io_r0_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [21:0] metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 479:25]
  wire [21:0] metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 479:25]
  wire [21:0] metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 479:25]
  wire [21:0] metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 479:25]
  wire  metaArray_io_wreq_valid; // @[Cache.scala 479:25]
  wire [3:0] metaArray_io_wreq_bits_setIdx; // @[Cache.scala 479:25]
  wire [21:0] metaArray_io_wreq_bits_data_tag; // @[Cache.scala 479:25]
  wire  metaArray_io_wreq_bits_data_dirty; // @[Cache.scala 479:25]
  wire [3:0] metaArray_io_wreq_bits_waymask; // @[Cache.scala 479:25]
  wire  dataArray_clock; // @[Cache.scala 480:25]
  wire  dataArray_reset; // @[Cache.scala 480:25]
  wire  dataArray_io_r0_req_ready; // @[Cache.scala 480:25]
  wire  dataArray_io_r0_req_valid; // @[Cache.scala 480:25]
  wire [6:0] dataArray_io_r0_req_bits_setIdx; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r0_resp_data_0_data; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r0_resp_data_1_data; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r0_resp_data_2_data; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r0_resp_data_3_data; // @[Cache.scala 480:25]
  wire  dataArray_io_r1_req_ready; // @[Cache.scala 480:25]
  wire  dataArray_io_r1_req_valid; // @[Cache.scala 480:25]
  wire [6:0] dataArray_io_r1_req_bits_setIdx; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r1_resp_data_0_data; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r1_resp_data_1_data; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r1_resp_data_2_data; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r1_resp_data_3_data; // @[Cache.scala 480:25]
  wire  dataArray_io_wreq_valid; // @[Cache.scala 480:25]
  wire [6:0] dataArray_io_wreq_bits_setIdx; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_wreq_bits_data_data; // @[Cache.scala 480:25]
  wire [3:0] dataArray_io_wreq_bits_waymask; // @[Cache.scala 480:25]
  wire  arb_io_in_0_ready; // @[Cache.scala 489:19]
  wire  arb_io_in_0_valid; // @[Cache.scala 489:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[Cache.scala 489:19]
  wire [2:0] arb_io_in_0_bits_size; // @[Cache.scala 489:19]
  wire [86:0] arb_io_in_0_bits_user; // @[Cache.scala 489:19]
  wire  arb_io_out_ready; // @[Cache.scala 489:19]
  wire  arb_io_out_valid; // @[Cache.scala 489:19]
  wire [31:0] arb_io_out_bits_addr; // @[Cache.scala 489:19]
  wire [2:0] arb_io_out_bits_size; // @[Cache.scala 489:19]
  wire [86:0] arb_io_out_bits_user; // @[Cache.scala 489:19]
  wire  _T_2 = s2_io_out_ready & s2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T_2 ? 1'h0 : REG; // @[Pipeline.scala 25:25 Pipeline.scala 25:33 Pipeline.scala 24:24]
  wire  _T_4 = s1_io_out_valid & s2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = s1_io_out_valid & s2_io_in_ready | _GEN_0; // @[Pipeline.scala 26:38 Pipeline.scala 26:46]
  reg [31:0] REG_1_req_addr; // @[Reg.scala 27:20]
  reg [2:0] REG_1_req_size; // @[Reg.scala 27:20]
  reg [86:0] REG_1_req_user; // @[Reg.scala 27:20]
  reg  REG_2; // @[Pipeline.scala 24:24]
  wire  _GEN_9 = s3_io_isFinish ? 1'h0 : REG_2; // @[Pipeline.scala 25:25 Pipeline.scala 25:33 Pipeline.scala 24:24]
  wire  _T_7 = s2_io_out_valid & s3_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_10 = s2_io_out_valid & s3_io_in_ready | _GEN_9; // @[Pipeline.scala 26:38 Pipeline.scala 26:46]
  reg [31:0] REG_3_req_addr; // @[Reg.scala 27:20]
  reg [2:0] REG_3_req_size; // @[Reg.scala 27:20]
  reg [86:0] REG_3_req_user; // @[Reg.scala 27:20]
  reg [21:0] REG_3_metas_0_tag; // @[Reg.scala 27:20]
  reg [21:0] REG_3_metas_1_tag; // @[Reg.scala 27:20]
  reg [21:0] REG_3_metas_2_tag; // @[Reg.scala 27:20]
  reg [21:0] REG_3_metas_3_tag; // @[Reg.scala 27:20]
  reg [63:0] REG_3_datas_0_data; // @[Reg.scala 27:20]
  reg [63:0] REG_3_datas_1_data; // @[Reg.scala 27:20]
  reg [63:0] REG_3_datas_2_data; // @[Reg.scala 27:20]
  reg [63:0] REG_3_datas_3_data; // @[Reg.scala 27:20]
  reg  REG_3_hit; // @[Reg.scala 27:20]
  reg [3:0] REG_3_waymask; // @[Reg.scala 27:20]
  reg  REG_3_mmio; // @[Reg.scala 27:20]
  reg  REG_3_isForwardData; // @[Reg.scala 27:20]
  reg [63:0] REG_3_forwardData_data_data; // @[Reg.scala 27:20]
  reg [3:0] REG_3_forwardData_waymask; // @[Reg.scala 27:20]
  ysyx_210000_CacheStage1 s1 ( // @[Cache.scala 476:18]
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_size(s1_io_in_bits_size),
    .io_in_bits_user(s1_io_in_bits_user),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_size(s1_io_out_bits_req_size),
    .io_out_bits_req_user(s1_io_out_bits_req_user),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data)
  );
  ysyx_210000_CacheStage2 s2 ( // @[Cache.scala 477:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_size(s2_io_in_bits_req_size),
    .io_in_bits_req_user(s2_io_in_bits_req_user),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_size(s2_io_out_bits_req_size),
    .io_out_bits_req_user(s2_io_out_bits_req_user),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask)
  );
  ysyx_210000_CacheStage3 s3 ( // @[Cache.scala 478:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_size(s3_io_in_bits_req_size),
    .io_in_bits_req_user(s3_io_in_bits_req_user),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_ready(s3_io_out_ready),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_out_bits_user(s3_io_out_bits_user),
    .io_isFinish(s3_io_isFinish),
    .io_flush(s3_io_flush),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_mmio_req_ready(s3_io_mmio_req_ready),
    .io_mmio_req_valid(s3_io_mmio_req_valid),
    .io_mmio_req_bits_addr(s3_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(s3_io_mmio_req_bits_size),
    .io_mmio_resp_ready(s3_io_mmio_resp_ready),
    .io_mmio_resp_valid(s3_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(s3_io_mmio_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid)
  );
  ysyx_210000_SRAMTemplateWithArbiter metaArray ( // @[Cache.scala 479:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r0_req_ready(metaArray_io_r0_req_ready),
    .io_r0_req_valid(metaArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(metaArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_tag(metaArray_io_r0_resp_data_0_tag),
    .io_r0_resp_data_0_valid(metaArray_io_r0_resp_data_0_valid),
    .io_r0_resp_data_0_dirty(metaArray_io_r0_resp_data_0_dirty),
    .io_r0_resp_data_1_tag(metaArray_io_r0_resp_data_1_tag),
    .io_r0_resp_data_1_valid(metaArray_io_r0_resp_data_1_valid),
    .io_r0_resp_data_1_dirty(metaArray_io_r0_resp_data_1_dirty),
    .io_r0_resp_data_2_tag(metaArray_io_r0_resp_data_2_tag),
    .io_r0_resp_data_2_valid(metaArray_io_r0_resp_data_2_valid),
    .io_r0_resp_data_2_dirty(metaArray_io_r0_resp_data_2_dirty),
    .io_r0_resp_data_3_tag(metaArray_io_r0_resp_data_3_tag),
    .io_r0_resp_data_3_valid(metaArray_io_r0_resp_data_3_valid),
    .io_r0_resp_data_3_dirty(metaArray_io_r0_resp_data_3_dirty),
    .io_wreq_valid(metaArray_io_wreq_valid),
    .io_wreq_bits_setIdx(metaArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(metaArray_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(metaArray_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(metaArray_io_wreq_bits_waymask)
  );
  ysyx_210000_SRAMTemplateWithArbiter_1 dataArray ( // @[Cache.scala 480:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r0_req_ready(dataArray_io_r0_req_ready),
    .io_r0_req_valid(dataArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(dataArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_data(dataArray_io_r0_resp_data_0_data),
    .io_r0_resp_data_1_data(dataArray_io_r0_resp_data_1_data),
    .io_r0_resp_data_2_data(dataArray_io_r0_resp_data_2_data),
    .io_r0_resp_data_3_data(dataArray_io_r0_resp_data_3_data),
    .io_r1_req_ready(dataArray_io_r1_req_ready),
    .io_r1_req_valid(dataArray_io_r1_req_valid),
    .io_r1_req_bits_setIdx(dataArray_io_r1_req_bits_setIdx),
    .io_r1_resp_data_0_data(dataArray_io_r1_resp_data_0_data),
    .io_r1_resp_data_1_data(dataArray_io_r1_resp_data_1_data),
    .io_r1_resp_data_2_data(dataArray_io_r1_resp_data_2_data),
    .io_r1_resp_data_3_data(dataArray_io_r1_resp_data_3_data),
    .io_wreq_valid(dataArray_io_wreq_valid),
    .io_wreq_bits_setIdx(dataArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(dataArray_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(dataArray_io_wreq_bits_waymask)
  );
  ysyx_210000_Arbiter_4 arb ( // @[Cache.scala 489:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_size(arb_io_in_0_bits_size),
    .io_in_0_bits_user(arb_io_in_0_bits_user),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_size(arb_io_out_bits_size),
    .io_out_bits_user(arb_io_out_bits_user)
  );
  assign io_in_req_ready = arb_io_in_0_ready; // @[Cache.scala 490:28]
  assign io_in_resp_valid = s3_io_out_valid; // @[Cache.scala 506:100]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[Cache.scala 500:14]
  assign io_in_resp_bits_user = s3_io_out_bits_user; // @[Cache.scala 500:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[Cache.scala 502:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[Cache.scala 502:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[Cache.scala 502:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[Cache.scala 502:14]
  assign io_mmio_req_valid = s3_io_mmio_req_valid; // @[Cache.scala 503:11]
  assign io_mmio_req_bits_addr = s3_io_mmio_req_bits_addr; // @[Cache.scala 503:11]
  assign io_mmio_req_bits_size = s3_io_mmio_req_bits_size; // @[Cache.scala 503:11]
  assign io_empty = ~s2_io_in_valid & ~s3_io_in_valid; // @[Cache.scala 504:31]
  assign s1_io_in_valid = arb_io_out_valid; // @[Cache.scala 492:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[Cache.scala 492:12]
  assign s1_io_in_bits_size = arb_io_out_bits_size; // @[Cache.scala 492:12]
  assign s1_io_in_bits_user = arb_io_out_bits_user; // @[Cache.scala 492:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r0_req_ready; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r0_req_ready; // @[Cache.scala 525:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r0_resp_data_0_data; // @[Cache.scala 525:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r0_resp_data_1_data; // @[Cache.scala 525:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r0_resp_data_2_data; // @[Cache.scala 525:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r0_resp_data_3_data; // @[Cache.scala 525:21]
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = REG; // @[Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = REG_1_req_addr; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_size = REG_1_req_size; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_user = REG_1_req_user; // @[Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 532:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 532:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 532:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 532:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 534:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 534:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 534:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 534:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 533:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 533:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 533:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 533:22]
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = REG_2; // @[Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = REG_3_req_addr; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_size = REG_3_req_size; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_user = REG_3_req_user; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = REG_3_metas_0_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = REG_3_metas_1_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = REG_3_metas_2_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = REG_3_metas_3_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = REG_3_datas_0_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = REG_3_datas_1_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = REG_3_datas_2_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = REG_3_datas_3_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = REG_3_hit; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = REG_3_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = REG_3_mmio; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = REG_3_isForwardData; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = REG_3_forwardData_data_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = REG_3_forwardData_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_out_ready = io_in_resp_ready; // @[Cache.scala 500:14]
  assign s3_io_flush = io_flush[1]; // @[Cache.scala 501:26]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r1_req_ready; // @[Cache.scala 526:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r1_resp_data_0_data; // @[Cache.scala 526:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r1_resp_data_1_data; // @[Cache.scala 526:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r1_resp_data_2_data; // @[Cache.scala 526:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r1_resp_data_3_data; // @[Cache.scala 526:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[Cache.scala 502:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[Cache.scala 502:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[Cache.scala 502:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[Cache.scala 502:14]
  assign s3_io_mmio_req_ready = io_mmio_req_ready; // @[Cache.scala 503:11]
  assign s3_io_mmio_resp_valid = io_mmio_resp_valid; // @[Cache.scala 503:11]
  assign s3_io_mmio_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[Cache.scala 503:11]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset | MOUFlushICache; // @[Cache.scala 486:37]
  assign metaArray_io_r0_req_valid = s1_io_metaReadBus_req_valid; // @[Cache.scala 524:21]
  assign metaArray_io_r0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 524:21]
  assign metaArray_io_wreq_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 528:18]
  assign metaArray_io_wreq_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 528:18]
  assign metaArray_io_wreq_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 528:18]
  assign metaArray_io_wreq_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 528:18]
  assign metaArray_io_wreq_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 528:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r0_req_valid = s1_io_dataReadBus_req_valid; // @[Cache.scala 525:21]
  assign dataArray_io_r0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 525:21]
  assign dataArray_io_r1_req_valid = s3_io_dataReadBus_req_valid; // @[Cache.scala 526:21]
  assign dataArray_io_r1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 526:21]
  assign dataArray_io_wreq_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 529:18]
  assign dataArray_io_wreq_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 529:18]
  assign dataArray_io_wreq_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 529:18]
  assign dataArray_io_wreq_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 529:18]
  assign arb_io_in_0_valid = io_in_req_valid; // @[Cache.scala 490:28]
  assign arb_io_in_0_bits_addr = io_in_req_bits_addr; // @[Cache.scala 490:28]
  assign arb_io_in_0_bits_size = io_in_req_bits_size; // @[Cache.scala 490:28]
  assign arb_io_in_0_bits_user = io_in_req_bits_user; // @[Cache.scala 490:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[Cache.scala 492:12]
  always @(posedge clock) begin
    if (reset) begin // @[Pipeline.scala 24:24]
      REG <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (io_flush[0]) begin // @[Pipeline.scala 27:20]
      REG <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG <= _GEN_1;
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_req_addr <= 32'h0; // @[Reg.scala 27:20]
    end else if (_T_4) begin // @[Reg.scala 28:19]
      REG_1_req_addr <= s1_io_out_bits_req_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_req_size <= 3'h0; // @[Reg.scala 27:20]
    end else if (_T_4) begin // @[Reg.scala 28:19]
      REG_1_req_size <= s1_io_out_bits_req_size; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_req_user <= 87'h0; // @[Reg.scala 27:20]
    end else if (_T_4) begin // @[Reg.scala 28:19]
      REG_1_req_user <= s1_io_out_bits_req_user; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Pipeline.scala 24:24]
      REG_2 <= 1'h0; // @[Pipeline.scala 24:24]
    end else if (io_flush[1]) begin // @[Pipeline.scala 27:20]
      REG_2 <= 1'h0; // @[Pipeline.scala 27:28]
    end else begin
      REG_2 <= _GEN_10;
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_req_addr <= 32'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_req_addr <= s2_io_out_bits_req_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_req_size <= 3'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_req_size <= s2_io_out_bits_req_size; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_req_user <= 87'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_req_user <= s2_io_out_bits_req_user; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_metas_0_tag <= 22'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_metas_0_tag <= s2_io_out_bits_metas_0_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_metas_1_tag <= 22'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_metas_1_tag <= s2_io_out_bits_metas_1_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_metas_2_tag <= 22'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_metas_2_tag <= s2_io_out_bits_metas_2_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_metas_3_tag <= 22'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_metas_3_tag <= s2_io_out_bits_metas_3_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_datas_0_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_datas_0_data <= s2_io_out_bits_datas_0_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_datas_1_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_datas_1_data <= s2_io_out_bits_datas_1_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_datas_2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_datas_2_data <= s2_io_out_bits_datas_2_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_datas_3_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_datas_3_data <= s2_io_out_bits_datas_3_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_hit <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_hit <= s2_io_out_bits_hit; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_waymask <= 4'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_waymask <= s2_io_out_bits_waymask; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_mmio <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_mmio <= s2_io_out_bits_mmio; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_isForwardData <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_isForwardData <= s2_io_out_bits_isForwardData; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_forwardData_data_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_forwardData_data_data <= s2_io_out_bits_forwardData_data_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_forwardData_waymask <= 4'h0; // @[Reg.scala 27:20]
    end else if (_T_7) begin // @[Reg.scala 28:19]
      REG_3_forwardData_waymask <= s2_io_out_bits_forwardData_waymask; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1_req_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  REG_1_req_size = _RAND_2[2:0];
  _RAND_3 = {3{`RANDOM}};
  REG_1_req_user = _RAND_3[86:0];
  _RAND_4 = {1{`RANDOM}};
  REG_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG_3_req_addr = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  REG_3_req_size = _RAND_6[2:0];
  _RAND_7 = {3{`RANDOM}};
  REG_3_req_user = _RAND_7[86:0];
  _RAND_8 = {1{`RANDOM}};
  REG_3_metas_0_tag = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  REG_3_metas_1_tag = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  REG_3_metas_2_tag = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  REG_3_metas_3_tag = _RAND_11[21:0];
  _RAND_12 = {2{`RANDOM}};
  REG_3_datas_0_data = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  REG_3_datas_1_data = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  REG_3_datas_2_data = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  REG_3_datas_3_data = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  REG_3_hit = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  REG_3_waymask = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  REG_3_mmio = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  REG_3_isForwardData = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  REG_3_forwardData_data_data = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  REG_3_forwardData_waymask = _RAND_21[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_EmbeddedTLBExec_1(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [38:0]  io_in_bits_addr,
  input  [2:0]   io_in_bits_size,
  input  [3:0]   io_in_bits_cmd,
  input  [7:0]   io_in_bits_wmask,
  input  [63:0]  io_in_bits_wdata,
  input          io_out_ready,
  output         io_out_valid,
  output [31:0]  io_out_bits_addr,
  output [2:0]   io_out_bits_size,
  output [3:0]   io_out_bits_cmd,
  output [7:0]   io_out_bits_wmask,
  output [63:0]  io_out_bits_wdata,
  input  [120:0] io_md_0,
  input  [120:0] io_md_1,
  input  [120:0] io_md_2,
  input  [120:0] io_md_3,
  output         io_mdWrite_wen,
  output [3:0]   io_mdWrite_windex,
  output [3:0]   io_mdWrite_waymask,
  output [120:0] io_mdWrite_wdata,
  input          io_mdReady,
  input          io_mem_req_ready,
  output         io_mem_req_valid,
  output [31:0]  io_mem_req_bits_addr,
  output [3:0]   io_mem_req_bits_cmd,
  output [63:0]  io_mem_req_bits_wdata,
  output         io_mem_resp_ready,
  input          io_mem_resp_valid,
  input  [63:0]  io_mem_resp_bits_rdata,
  input  [63:0]  io_satp,
  input  [1:0]   io_pf_priviledgeMode,
  input          io_pf_status_sum,
  input          io_pf_status_mxr,
  output         io_pf_loadPF,
  output         io_pf_storePF,
  output [38:0]  io_pf_addr,
  output         io_isFinish,
  input          ISAMO
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[EmbeddedTLB.scala 193:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[EmbeddedTLB.scala 193:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[EmbeddedTLB.scala 193:54]
  wire [19:0] satp_ppn = io_satp[19:0]; // @[EmbeddedTLB.scala 195:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[EmbeddedTLB.scala 195:30]
  wire [26:0] _T_43 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[EmbeddedTLB.scala 204:201]
  wire [26:0] _T_44 = {9'h1ff,io_md_0[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_45 = _T_44 & io_md_0[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_47 = _T_44 & _T_43; // @[TLB.scala 131:84]
  wire  _T_48 = _T_45 == _T_47; // @[TLB.scala 131:48]
  wire  _T_49 = io_md_0[52] & io_md_0[93:78] == satp_asid & _T_48; // @[EmbeddedTLB.scala 204:132]
  wire [26:0] _T_85 = {9'h1ff,io_md_1[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_86 = _T_85 & io_md_1[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_88 = _T_85 & _T_43; // @[TLB.scala 131:84]
  wire  _T_89 = _T_86 == _T_88; // @[TLB.scala 131:48]
  wire  _T_90 = io_md_1[52] & io_md_1[93:78] == satp_asid & _T_89; // @[EmbeddedTLB.scala 204:132]
  wire [26:0] _T_126 = {9'h1ff,io_md_2[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_127 = _T_126 & io_md_2[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_129 = _T_126 & _T_43; // @[TLB.scala 131:84]
  wire  _T_130 = _T_127 == _T_129; // @[TLB.scala 131:48]
  wire  _T_131 = io_md_2[52] & io_md_2[93:78] == satp_asid & _T_130; // @[EmbeddedTLB.scala 204:132]
  wire [26:0] _T_167 = {9'h1ff,io_md_3[77:60]}; // @[Cat.scala 30:58]
  wire [26:0] _T_168 = _T_167 & io_md_3[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_170 = _T_167 & _T_43; // @[TLB.scala 131:84]
  wire  _T_171 = _T_168 == _T_170; // @[TLB.scala 131:48]
  wire  _T_172 = io_md_3[52] & io_md_3[93:78] == satp_asid & _T_171; // @[EmbeddedTLB.scala 204:132]
  wire [3:0] hitVec = {_T_172,_T_131,_T_90,_T_49}; // @[EmbeddedTLB.scala 204:211]
  wire  _T_173 = |hitVec; // @[EmbeddedTLB.scala 205:35]
  wire  hit = io_in_valid & |hitVec; // @[EmbeddedTLB.scala 205:25]
  wire  miss = io_in_valid & ~_T_173; // @[EmbeddedTLB.scala 206:26]
  reg [63:0] REG; // @[LFSR64.scala 25:23]
  wire  hi_5 = REG[0] ^ REG[1] ^ REG[3] ^ REG[4]; // @[LFSR64.scala 26:43]
  wire [62:0] lo_1 = REG[63:1]; // @[LFSR64.scala 28:51]
  wire [63:0] _T_183 = {hi_5,lo_1}; // @[Cat.scala 30:58]
  wire [3:0] victimWaymask = 4'h1 << REG[1:0]; // @[EmbeddedTLB.scala 208:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[EmbeddedTLB.scala 209:20]
  wire [120:0] _T_190 = waymask[0] ? io_md_0 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_191 = waymask[1] ? io_md_1 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_192 = waymask[2] ? io_md_2 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_193 = waymask[3] ? io_md_3 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_194 = _T_190 | _T_191; // @[Mux.scala 27:72]
  wire [120:0] _T_195 = _T_194 | _T_192; // @[Mux.scala 27:72]
  wire [120:0] _T_196 = _T_195 | _T_193; // @[Mux.scala 27:72]
  wire [7:0] hitMeta_flag = _T_196[59:52]; // @[EmbeddedTLB.scala 215:70]
  wire [17:0] hitMeta_mask = _T_196[77:60]; // @[EmbeddedTLB.scala 215:70]
  wire [15:0] hitMeta_asid = _T_196[93:78]; // @[EmbeddedTLB.scala 215:70]
  wire [31:0] hitData_pteaddr = _T_196[31:0]; // @[EmbeddedTLB.scala 216:70]
  wire [19:0] hitData_ppn = _T_196[51:32]; // @[EmbeddedTLB.scala 216:70]
  wire  hitFlag_v = hitMeta_flag[0]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_r = hitMeta_flag[1]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_g = hitMeta_flag[5]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[EmbeddedTLB.scala 217:38]
  reg [2:0] state; // @[EmbeddedTLB.scala 247:22]
  wire  _T_294 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_241 = io_pf_priviledgeMode == 2'h0; // @[EmbeddedTLB.scala 226:62]
  wire  _T_246 = io_pf_priviledgeMode == 2'h1; // @[EmbeddedTLB.scala 226:110]
  wire  _T_248 = ~io_pf_status_sum; // @[EmbeddedTLB.scala 226:137]
  wire  hitCheck = hit & ~(io_pf_priviledgeMode == 2'h0 & ~hitFlag_u) & ~(io_pf_priviledgeMode == 2'h1 & hitFlag_u & ~
    io_pf_status_sum); // @[EmbeddedTLB.scala 226:87]
  wire  hitLoad = hitCheck & (hitFlag_r | io_pf_status_mxr & hitFlag_x); // @[EmbeddedTLB.scala 228:26]
  wire  _T_259 = ~io_in_bits_cmd[0] & ~io_in_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_261 = ~hitLoad & _T_259 & hit; // @[EmbeddedTLB.scala 241:40]
  wire  _T_262 = ~ISAMO; // @[EmbeddedTLB.scala 241:50]
  wire  _T_300 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_302 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_312 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[EmbeddedTLB.scala 255:49]
  wire [7:0] _T_303 = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,memRdata_flag_w,
    memRdata_flag_r,memRdata_flag_v}; // @[EmbeddedTLB.scala 292:44]
  reg [1:0] level; // @[EmbeddedTLB.scala 248:22]
  wire  _T_315 = level == 2'h3; // @[EmbeddedTLB.scala 297:58]
  wire  _T_316 = level == 2'h2; // @[EmbeddedTLB.scala 297:73]
  wire  _T_329 = _T_259 & _T_262; // @[EmbeddedTLB.scala 302:38]
  wire  _GEN_19 = ~_T_303[0] | ~_T_303[1] & _T_303[2] ? _T_259 & _T_262 : ~hitLoad & _T_259 & hit & ~ISAMO; // @[EmbeddedTLB.scala 298:60 EmbeddedTLB.scala 302:22 EmbeddedTLB.scala 241:12]
  wire  _T_358 = _T_303[0] & ~(_T_241 & ~_T_303[4]) & ~(_T_246 & _T_303[4] & _T_248); // @[EmbeddedTLB.scala 314:87]
  wire  _T_362 = _T_358 & (_T_303[1] | io_pf_status_mxr & _T_303[3]); // @[EmbeddedTLB.scala 316:36]
  wire  _T_363 = _T_358 & _T_303[2]; // @[EmbeddedTLB.scala 317:37]
  wire  _GEN_23 = ~_T_362 & _T_259 | ~_T_363 & io_in_bits_cmd[0] ? _T_329 : ~hitLoad & _T_259 & hit & ~ISAMO; // @[EmbeddedTLB.scala 330:80 EmbeddedTLB.scala 332:22 EmbeddedTLB.scala 241:12]
  wire  _GEN_29 = level != 2'h0 ? _GEN_23 : ~hitLoad & _T_259 & hit & ~ISAMO; // @[EmbeddedTLB.scala 313:36 EmbeddedTLB.scala 241:12]
  wire  _GEN_35 = ~(_T_303[1] | _T_303[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_19 : _GEN_29; // @[EmbeddedTLB.scala 297:82]
  wire  _GEN_54 = _T_312 ? _GEN_35 : ~hitLoad & _T_259 & hit & ~ISAMO; // @[EmbeddedTLB.scala 293:33 EmbeddedTLB.scala 241:12]
  wire  _GEN_78 = _T_302 ? _GEN_54 : ~hitLoad & _T_259 & hit & ~ISAMO; // @[Conditional.scala 39:67 EmbeddedTLB.scala 241:12]
  wire  _GEN_91 = _T_300 ? ~hitLoad & _T_259 & hit & ~ISAMO : _GEN_78; // @[Conditional.scala 39:67 EmbeddedTLB.scala 241:12]
  wire  loadPF = _T_294 ? ~hitLoad & _T_259 & hit & ~ISAMO : _GEN_91; // @[Conditional.scala 40:58 EmbeddedTLB.scala 241:12]
  wire  hitStore = hitCheck & hitFlag_w; // @[EmbeddedTLB.scala 229:27]
  wire  _T_331 = io_in_bits_cmd[0] | ISAMO; // @[EmbeddedTLB.scala 303:40]
  wire  _GEN_20 = ~_T_303[0] | ~_T_303[1] & _T_303[2] ? io_in_bits_cmd[0] | ISAMO : ~hitStore & io_in_bits_cmd[0] & hit
     | _T_261 & ISAMO; // @[EmbeddedTLB.scala 298:60 EmbeddedTLB.scala 303:23 EmbeddedTLB.scala 242:13]
  wire  _GEN_24 = ~_T_362 & _T_259 | ~_T_363 & io_in_bits_cmd[0] ? _T_331 : ~hitStore & io_in_bits_cmd[0] & hit | _T_261
     & ISAMO; // @[EmbeddedTLB.scala 330:80 EmbeddedTLB.scala 333:23 EmbeddedTLB.scala 242:13]
  wire  _GEN_30 = level != 2'h0 ? _GEN_24 : ~hitStore & io_in_bits_cmd[0] & hit | _T_261 & ISAMO; // @[EmbeddedTLB.scala 313:36 EmbeddedTLB.scala 242:13]
  wire  _GEN_36 = ~(_T_303[1] | _T_303[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_20 : _GEN_30; // @[EmbeddedTLB.scala 297:82]
  wire  _GEN_55 = _T_312 ? _GEN_36 : ~hitStore & io_in_bits_cmd[0] & hit | _T_261 & ISAMO; // @[EmbeddedTLB.scala 293:33 EmbeddedTLB.scala 242:13]
  wire  _GEN_79 = _T_302 ? _GEN_55 : ~hitStore & io_in_bits_cmd[0] & hit | _T_261 & ISAMO; // @[Conditional.scala 39:67 EmbeddedTLB.scala 242:13]
  wire  _GEN_92 = _T_300 ? ~hitStore & io_in_bits_cmd[0] & hit | _T_261 & ISAMO : _GEN_79; // @[Conditional.scala 39:67 EmbeddedTLB.scala 242:13]
  wire  storePF = _T_294 ? ~hitStore & io_in_bits_cmd[0] & hit | _T_261 & ISAMO : _GEN_92; // @[Conditional.scala 40:58 EmbeddedTLB.scala 242:13]
  wire  _T_235 = io_pf_loadPF | io_pf_storePF; // @[Bundle.scala 133:23]
  wire  hitWB = hit & (~hitFlag_a | ~hitFlag_d & io_in_bits_cmd[0]) & ~(loadPF | storePF | _T_235); // @[EmbeddedTLB.scala 221:81]
  wire [7:0] _T_238 = {io_in_bits_cmd[0],1'h1,6'h0}; // @[Cat.scala 30:58]
  wire [7:0] _T_239 = {hitFlag_d,hitFlag_a,hitFlag_g,hitFlag_u,hitFlag_x,hitFlag_w,hitFlag_r,hitFlag_v}; // @[EmbeddedTLB.scala 222:79]
  wire [7:0] hitRefillFlag = _T_238 | _T_239; // @[EmbeddedTLB.scala 222:69]
  wire [39:0] _T_240 = {10'h0,hitData_ppn,2'h0,hitRefillFlag}; // @[Cat.scala 30:58]
  reg [39:0] hitWBStore; // @[Reg.scala 27:20]
  reg  REG_1; // @[EmbeddedTLB.scala 236:26]
  reg  REG_2; // @[EmbeddedTLB.scala 237:27]
  reg [63:0] memRespStore; // @[EmbeddedTLB.scala 250:29]
  reg [17:0] missMaskStore; // @[EmbeddedTLB.scala 252:30]
  wire [19:0] memRdata_ppn = io_mem_resp_bits_rdata[29:10]; // @[EmbeddedTLB.scala 255:49]
  reg [31:0] raddr; // @[EmbeddedTLB.scala 256:22]
  wire  _T_289 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_2 = _T_289 | alreadyOutFire; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [31:0] _T_299 = {satp_ppn,vpn_vpn2,3'h0}; // @[Cat.scala 30:58]
  wire  _T_301 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [8:0] lo_5 = _T_315 ? vpn_vpn1 : vpn_vpn0; // @[EmbeddedTLB.scala 311:50]
  wire [31:0] _T_345 = {memRdata_ppn,lo_5,3'h0}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_18 = ~_T_303[0] | ~_T_303[1] & _T_303[2] ? 3'h5 : 3'h1; // @[EmbeddedTLB.scala 298:60 EmbeddedTLB.scala 299:73 EmbeddedTLB.scala 310:19]
  wire [31:0] _GEN_21 = ~_T_303[0] | ~_T_303[1] & _T_303[2] ? raddr : _T_345; // @[EmbeddedTLB.scala 298:60 EmbeddedTLB.scala 256:22 EmbeddedTLB.scala 311:19]
  wire  _T_368 = ~_T_303[6] | ~_T_303[7] & io_in_bits_cmd[0]; // @[EmbeddedTLB.scala 318:72]
  wire [63:0] _T_369 = {56'h0,io_in_bits_cmd[0],7'h40}; // @[Cat.scala 30:58]
  wire [7:0] _T_371 = {_T_303[7],_T_303[6],_T_303[5],_T_303[4],_T_303[3],_T_303[2],_T_303[1],_T_303[0]}; // @[EmbeddedTLB.scala 320:79]
  wire [7:0] _T_372 = _T_238 | _T_371; // @[EmbeddedTLB.scala 320:68]
  wire [63:0] _T_373 = io_mem_resp_bits_rdata | _T_369; // @[EmbeddedTLB.scala 321:50]
  wire [2:0] _T_394 = _T_368 ? 3'h3 : 3'h4; // @[EmbeddedTLB.scala 335:27]
  wire [2:0] _GEN_22 = ~_T_362 & _T_259 | ~_T_363 & io_in_bits_cmd[0] ? 3'h5 : _T_394; // @[EmbeddedTLB.scala 330:80 EmbeddedTLB.scala 331:21 EmbeddedTLB.scala 335:21]
  wire  _GEN_25 = ~_T_362 & _T_259 | ~_T_363 & io_in_bits_cmd[0] ? 1'h0 : 1'h1; // @[EmbeddedTLB.scala 330:80 EmbeddedTLB.scala 336:30]
  wire [17:0] _T_397 = _T_316 ? 18'h3fe00 : 18'h3ffff; // @[EmbeddedTLB.scala 339:59]
  wire [17:0] _T_398 = _T_315 ? 18'h0 : _T_397; // @[EmbeddedTLB.scala 339:26]
  wire [7:0] _GEN_26 = level != 2'h0 ? _T_372 : 8'h0; // @[EmbeddedTLB.scala 313:36 EmbeddedTLB.scala 320:26]
  wire [63:0] _GEN_27 = level != 2'h0 ? _T_373 : memRespStore; // @[EmbeddedTLB.scala 313:36 EmbeddedTLB.scala 321:24 EmbeddedTLB.scala 250:29]
  wire [2:0] _GEN_28 = level != 2'h0 ? _GEN_22 : state; // @[EmbeddedTLB.scala 313:36 EmbeddedTLB.scala 247:22]
  wire  _GEN_31 = level != 2'h0 & _GEN_25; // @[EmbeddedTLB.scala 313:36]
  wire [17:0] _GEN_32 = level != 2'h0 ? _T_398 : 18'h3ffff; // @[EmbeddedTLB.scala 313:36 EmbeddedTLB.scala 339:20]
  wire [17:0] _GEN_41 = ~(_T_303[1] | _T_303[3]) & (level == 2'h3 | level == 2'h2) ? 18'h3ffff : _GEN_32; // @[EmbeddedTLB.scala 297:82]
  wire [17:0] _GEN_60 = _T_312 ? _GEN_41 : 18'h3ffff; // @[EmbeddedTLB.scala 293:33]
  wire [17:0] _GEN_84 = _T_302 ? _GEN_60 : 18'h3ffff; // @[Conditional.scala 39:67]
  wire [17:0] _GEN_97 = _T_300 ? 18'h3ffff : _GEN_84; // @[Conditional.scala 39:67]
  wire [17:0] missMask = _T_294 ? 18'h3ffff : _GEN_97; // @[Conditional.scala 40:58]
  wire [17:0] _GEN_33 = level != 2'h0 ? missMask : missMaskStore; // @[EmbeddedTLB.scala 313:36 EmbeddedTLB.scala 340:25 EmbeddedTLB.scala 252:30]
  wire [2:0] _GEN_34 = ~(_T_303[1] | _T_303[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_18 : _GEN_28; // @[EmbeddedTLB.scala 297:82]
  wire [31:0] _GEN_37 = ~(_T_303[1] | _T_303[3]) & (level == 2'h3 | level == 2'h2) ? _GEN_21 : raddr; // @[EmbeddedTLB.scala 297:82 EmbeddedTLB.scala 256:22]
  wire [7:0] _GEN_38 = ~(_T_303[1] | _T_303[3]) & (level == 2'h3 | level == 2'h2) ? 8'h0 : _GEN_26; // @[EmbeddedTLB.scala 297:82]
  wire [63:0] _GEN_39 = ~(_T_303[1] | _T_303[3]) & (level == 2'h3 | level == 2'h2) ? memRespStore : _GEN_27; // @[EmbeddedTLB.scala 297:82 EmbeddedTLB.scala 250:29]
  wire  _GEN_40 = ~(_T_303[1] | _T_303[3]) & (level == 2'h3 | level == 2'h2) ? 1'h0 : _GEN_31; // @[EmbeddedTLB.scala 297:82]
  wire [17:0] _GEN_42 = ~(_T_303[1] | _T_303[3]) & (level == 2'h3 | level == 2'h2) ? missMaskStore : _GEN_33; // @[EmbeddedTLB.scala 297:82 EmbeddedTLB.scala 252:30]
  wire [1:0] _T_400 = level - 2'h1; // @[EmbeddedTLB.scala 342:24]
  wire [2:0] _GEN_52 = _T_312 ? _GEN_34 : state; // @[EmbeddedTLB.scala 293:33 EmbeddedTLB.scala 247:22]
  wire [31:0] _GEN_56 = _T_312 ? _GEN_37 : raddr; // @[EmbeddedTLB.scala 293:33 EmbeddedTLB.scala 256:22]
  wire [7:0] _GEN_57 = _T_312 ? _GEN_38 : 8'h0; // @[EmbeddedTLB.scala 293:33]
  wire [63:0] _GEN_58 = _T_312 ? _GEN_39 : memRespStore; // @[EmbeddedTLB.scala 293:33 EmbeddedTLB.scala 250:29]
  wire  _GEN_59 = _T_312 & _GEN_40; // @[EmbeddedTLB.scala 293:33]
  wire [17:0] _GEN_61 = _T_312 ? _GEN_42 : missMaskStore; // @[EmbeddedTLB.scala 293:33 EmbeddedTLB.scala 252:30]
  wire [1:0] _GEN_62 = _T_312 ? _T_400 : level; // @[EmbeddedTLB.scala 293:33 EmbeddedTLB.scala 342:15 EmbeddedTLB.scala 248:22]
  wire  _T_401 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_63 = _T_301 ? 3'h4 : state; // @[EmbeddedTLB.scala 350:38 EmbeddedTLB.scala 350:46 EmbeddedTLB.scala 247:22]
  wire  _T_403 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_65 = _GEN_2 ? 3'h0 : state; // @[EmbeddedTLB.scala 353:73 EmbeddedTLB.scala 354:13 EmbeddedTLB.scala 247:22]
  wire  _GEN_67 = _GEN_2 ? 1'h0 : _GEN_2; // @[EmbeddedTLB.scala 353:73 EmbeddedTLB.scala 356:22]
  wire  _T_407 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_68 = _T_407 ? 3'h0 : state; // @[Conditional.scala 39:67 EmbeddedTLB.scala 360:13 EmbeddedTLB.scala 247:22]
  wire [2:0] _GEN_69 = _T_403 ? _GEN_65 : _GEN_68; // @[Conditional.scala 39:67]
  wire  _GEN_71 = _T_403 ? _GEN_67 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_72 = _T_401 ? _GEN_63 : _GEN_69; // @[Conditional.scala 39:67]
  wire  _GEN_75 = _T_401 ? _GEN_2 : _GEN_71; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_81 = _T_302 ? _GEN_57 : 8'h0; // @[Conditional.scala 39:67]
  wire  _GEN_96 = _T_300 ? 1'h0 : _T_302 & _GEN_59; // @[Conditional.scala 39:67]
  wire  missMetaRefill = _T_294 ? 1'h0 : _GEN_96; // @[Conditional.scala 40:58]
  wire  cmd = state == 3'h3; // @[EmbeddedTLB.scala 365:23]
  wire  _T_418 = state == 3'h0; // @[EmbeddedTLB.scala 371:82]
  reg  REG_7; // @[EmbeddedTLB.scala 371:33]
  reg [3:0] REG_8; // @[EmbeddedTLB.scala 372:21]
  reg [3:0] REG_9; // @[EmbeddedTLB.scala 372:65]
  reg [26:0] hi_hi_hi; // @[EmbeddedTLB.scala 372:94]
  reg [15:0] hi_hi_lo; // @[EmbeddedTLB.scala 373:19]
  reg [17:0] hi_lo_4; // @[EmbeddedTLB.scala 373:77]
  reg [7:0] lo_hi_hi; // @[EmbeddedTLB.scala 374:19]
  reg [19:0] lo_hi_lo; // @[EmbeddedTLB.scala 374:82]
  reg [31:0] lo_lo_3; // @[EmbeddedTLB.scala 375:22]
  wire [59:0] lo_8 = {lo_hi_hi,lo_hi_lo,lo_lo_3}; // @[Cat.scala 30:58]
  wire [60:0] hi_16 = {hi_hi_hi,hi_hi_lo,hi_lo_4}; // @[Cat.scala 30:58]
  wire [31:0] _T_434 = {hitData_ppn,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_435 = {2'h3,hitMeta_mask,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_436 = _T_434 & _T_435; // @[BitUtils.scala 32:13]
  wire [31:0] _T_437 = ~_T_435; // @[BitUtils.scala 32:38]
  wire [31:0] _T_438 = io_in_bits_addr[31:0] & _T_437; // @[BitUtils.scala 32:36]
  wire [31:0] _T_439 = _T_436 | _T_438; // @[BitUtils.scala 32:25]
  wire [31:0] _T_452 = {memRespStore[29:10],12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_453 = {2'h3,missMaskStore,12'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_454 = _T_452 & _T_453; // @[BitUtils.scala 32:13]
  wire [31:0] _T_455 = ~_T_453; // @[BitUtils.scala 32:38]
  wire [31:0] _T_456 = io_in_bits_addr[31:0] & _T_455; // @[BitUtils.scala 32:36]
  wire [31:0] _T_457 = _T_454 | _T_456; // @[BitUtils.scala 32:25]
  wire  _T_459 = ~hitWB; // @[EmbeddedTLB.scala 380:45]
  wire  _T_466 = hit & ~hitWB ? ~(_T_235 | loadPF | storePF) : state == 3'h4; // @[EmbeddedTLB.scala 380:37]
  assign io_in_ready = io_out_ready & _T_418 & ~miss & _T_459 & io_mdReady & (~_T_235 & ~loadPF & ~storePF); // @[EmbeddedTLB.scala 382:86]
  assign io_out_valid = io_in_valid & _T_466; // @[EmbeddedTLB.scala 380:31]
  assign io_out_bits_addr = hit ? _T_439 : _T_457; // @[EmbeddedTLB.scala 379:26]
  assign io_out_bits_size = io_in_bits_size; // @[EmbeddedTLB.scala 378:15]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[EmbeddedTLB.scala 378:15]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[EmbeddedTLB.scala 378:15]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[EmbeddedTLB.scala 378:15]
  assign io_mdWrite_wen = REG_7; // @[TLB.scala 214:14]
  assign io_mdWrite_windex = REG_8; // @[TLB.scala 215:17]
  assign io_mdWrite_waymask = REG_9; // @[TLB.scala 216:18]
  assign io_mdWrite_wdata = {hi_16,lo_8}; // @[Cat.scala 30:58]
  assign io_mem_req_valid = state == 3'h1 | cmd; // @[EmbeddedTLB.scala 367:48]
  assign io_mem_req_bits_addr = hitWB ? hitData_pteaddr : raddr; // @[EmbeddedTLB.scala 366:35]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[EmbeddedTLB.scala 365:23]
  assign io_mem_req_bits_wdata = hitWB ? {{24'd0}, hitWBStore} : memRespStore; // @[EmbeddedTLB.scala 366:138]
  assign io_mem_resp_ready = 1'h1; // @[EmbeddedTLB.scala 368:21]
  assign io_pf_loadPF = REG_1; // @[EmbeddedTLB.scala 236:16]
  assign io_pf_storePF = REG_2; // @[EmbeddedTLB.scala 237:17]
  assign io_pf_addr = io_in_bits_addr; // @[EmbeddedTLB.scala 201:11]
  assign io_isFinish = _T_289 | _T_235; // @[EmbeddedTLB.scala 385:32]
  always @(posedge clock) begin
    if (reset) begin // @[LFSR64.scala 25:23]
      REG <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG == 64'h0) begin // @[LFSR64.scala 28:18]
      REG <= 64'h1;
    end else begin
      REG <= _T_183;
    end
    if (reset) begin // @[EmbeddedTLB.scala 247:22]
      state <= 3'h0; // @[EmbeddedTLB.scala 247:22]
    end else if (_T_294) begin // @[Conditional.scala 40:58]
      if (hitWB) begin // @[EmbeddedTLB.scala 271:32]
        state <= 3'h3; // @[EmbeddedTLB.scala 272:15]
      end else if (miss) begin // @[EmbeddedTLB.scala 275:37]
        state <= 3'h1; // @[EmbeddedTLB.scala 276:15]
      end
    end else if (_T_300) begin // @[Conditional.scala 39:67]
      if (_T_301) begin // @[EmbeddedTLB.scala 288:38]
        state <= 3'h2; // @[EmbeddedTLB.scala 288:46]
      end
    end else if (_T_302) begin // @[Conditional.scala 39:67]
      state <= _GEN_52;
    end else begin
      state <= _GEN_72;
    end
    if (reset) begin // @[EmbeddedTLB.scala 248:22]
      level <= 2'h3; // @[EmbeddedTLB.scala 248:22]
    end else if (_T_294) begin // @[Conditional.scala 40:58]
      if (!(hitWB)) begin // @[EmbeddedTLB.scala 271:32]
        if (miss) begin // @[EmbeddedTLB.scala 275:37]
          level <= 2'h3; // @[EmbeddedTLB.scala 278:15]
        end
      end
    end else if (!(_T_300)) begin // @[Conditional.scala 39:67]
      if (_T_302) begin // @[Conditional.scala 39:67]
        level <= _GEN_62;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      hitWBStore <= 40'h0; // @[Reg.scala 27:20]
    end else if (hitWB) begin // @[Reg.scala 28:19]
      hitWBStore <= _T_240; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[EmbeddedTLB.scala 236:26]
      REG_1 <= 1'h0; // @[EmbeddedTLB.scala 236:26]
    end else if (_T_294) begin // @[Conditional.scala 40:58]
      REG_1 <= ~hitLoad & _T_259 & hit & ~ISAMO; // @[EmbeddedTLB.scala 241:12]
    end else if (_T_300) begin // @[Conditional.scala 39:67]
      REG_1 <= ~hitLoad & _T_259 & hit & ~ISAMO; // @[EmbeddedTLB.scala 241:12]
    end else if (_T_302) begin // @[Conditional.scala 39:67]
      REG_1 <= _GEN_54;
    end else begin
      REG_1 <= ~hitLoad & _T_259 & hit & ~ISAMO; // @[EmbeddedTLB.scala 241:12]
    end
    if (reset) begin // @[EmbeddedTLB.scala 237:27]
      REG_2 <= 1'h0; // @[EmbeddedTLB.scala 237:27]
    end else if (_T_294) begin // @[Conditional.scala 40:58]
      REG_2 <= ~hitStore & io_in_bits_cmd[0] & hit | _T_261 & ISAMO; // @[EmbeddedTLB.scala 242:13]
    end else if (_T_300) begin // @[Conditional.scala 39:67]
      REG_2 <= ~hitStore & io_in_bits_cmd[0] & hit | _T_261 & ISAMO; // @[EmbeddedTLB.scala 242:13]
    end else if (_T_302) begin // @[Conditional.scala 39:67]
      REG_2 <= _GEN_55;
    end else begin
      REG_2 <= ~hitStore & io_in_bits_cmd[0] & hit | _T_261 & ISAMO; // @[EmbeddedTLB.scala 242:13]
    end
    if (reset) begin // @[EmbeddedTLB.scala 250:29]
      memRespStore <= 64'h0; // @[EmbeddedTLB.scala 250:29]
    end else if (!(_T_294)) begin // @[Conditional.scala 40:58]
      if (!(_T_300)) begin // @[Conditional.scala 39:67]
        if (_T_302) begin // @[Conditional.scala 39:67]
          memRespStore <= _GEN_58;
        end
      end
    end
    if (reset) begin // @[EmbeddedTLB.scala 252:30]
      missMaskStore <= 18'h0; // @[EmbeddedTLB.scala 252:30]
    end else if (!(_T_294)) begin // @[Conditional.scala 40:58]
      if (!(_T_300)) begin // @[Conditional.scala 39:67]
        if (_T_302) begin // @[Conditional.scala 39:67]
          missMaskStore <= _GEN_61;
        end
      end
    end
    if (reset) begin // @[EmbeddedTLB.scala 256:22]
      raddr <= 32'h0; // @[EmbeddedTLB.scala 256:22]
    end else if (_T_294) begin // @[Conditional.scala 40:58]
      if (!(hitWB)) begin // @[EmbeddedTLB.scala 271:32]
        if (miss) begin // @[EmbeddedTLB.scala 275:37]
          raddr <= _T_299; // @[EmbeddedTLB.scala 277:15]
        end
      end
    end else if (!(_T_300)) begin // @[Conditional.scala 39:67]
      if (_T_302) begin // @[Conditional.scala 39:67]
        raddr <= _GEN_56;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      alreadyOutFire <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_294) begin // @[Conditional.scala 40:58]
      if (hitWB) begin // @[EmbeddedTLB.scala 271:32]
        alreadyOutFire <= 1'h0; // @[EmbeddedTLB.scala 274:24]
      end else if (miss) begin // @[EmbeddedTLB.scala 275:37]
        alreadyOutFire <= 1'h0; // @[EmbeddedTLB.scala 280:24]
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else if (_T_300) begin // @[Conditional.scala 39:67]
      alreadyOutFire <= _GEN_2;
    end else if (_T_302) begin // @[Conditional.scala 39:67]
      alreadyOutFire <= _GEN_2;
    end else begin
      alreadyOutFire <= _GEN_75;
    end
    if (reset) begin // @[EmbeddedTLB.scala 371:33]
      REG_7 <= 1'h0; // @[EmbeddedTLB.scala 371:33]
    end else begin
      REG_7 <= missMetaRefill | hitWB & state == 3'h0; // @[EmbeddedTLB.scala 371:33]
    end
    if (reset) begin // @[EmbeddedTLB.scala 372:21]
      REG_8 <= 4'h0; // @[EmbeddedTLB.scala 372:21]
    end else begin
      REG_8 <= io_in_bits_addr[15:12]; // @[EmbeddedTLB.scala 372:21]
    end
    if (reset) begin // @[EmbeddedTLB.scala 372:65]
      REG_9 <= 4'h0; // @[EmbeddedTLB.scala 372:65]
    end else if (hit) begin // @[EmbeddedTLB.scala 209:20]
      REG_9 <= hitVec;
    end else begin
      REG_9 <= victimWaymask;
    end
    if (reset) begin // @[EmbeddedTLB.scala 372:94]
      hi_hi_hi <= 27'h0; // @[EmbeddedTLB.scala 372:94]
    end else begin
      hi_hi_hi <= _T_43; // @[EmbeddedTLB.scala 372:94]
    end
    if (reset) begin // @[EmbeddedTLB.scala 373:19]
      hi_hi_lo <= 16'h0; // @[EmbeddedTLB.scala 373:19]
    end else if (hitWB) begin // @[EmbeddedTLB.scala 373:23]
      hi_hi_lo <= hitMeta_asid;
    end else begin
      hi_hi_lo <= satp_asid;
    end
    if (reset) begin // @[EmbeddedTLB.scala 373:77]
      hi_lo_4 <= 18'h0; // @[EmbeddedTLB.scala 373:77]
    end else if (hitWB) begin // @[EmbeddedTLB.scala 373:81]
      hi_lo_4 <= hitMeta_mask;
    end else if (_T_294) begin // @[Conditional.scala 40:58]
      hi_lo_4 <= 18'h3ffff;
    end else if (_T_300) begin // @[Conditional.scala 39:67]
      hi_lo_4 <= 18'h3ffff;
    end else begin
      hi_lo_4 <= _GEN_84;
    end
    if (reset) begin // @[EmbeddedTLB.scala 374:19]
      lo_hi_hi <= 8'h0; // @[EmbeddedTLB.scala 374:19]
    end else if (hitWB) begin // @[EmbeddedTLB.scala 374:23]
      lo_hi_hi <= hitRefillFlag;
    end else if (_T_294) begin // @[Conditional.scala 40:58]
      lo_hi_hi <= 8'h0;
    end else if (_T_300) begin // @[Conditional.scala 39:67]
      lo_hi_hi <= 8'h0;
    end else begin
      lo_hi_hi <= _GEN_81;
    end
    if (reset) begin // @[EmbeddedTLB.scala 374:82]
      lo_hi_lo <= 20'h0; // @[EmbeddedTLB.scala 374:82]
    end else if (hitWB) begin // @[EmbeddedTLB.scala 374:86]
      lo_hi_lo <= hitData_ppn;
    end else begin
      lo_hi_lo <= memRdata_ppn;
    end
    if (reset) begin // @[EmbeddedTLB.scala 375:22]
      lo_lo_3 <= 32'h0; // @[EmbeddedTLB.scala 375:22]
    end else if (hitWB) begin // @[EmbeddedTLB.scala 366:35]
      lo_lo_3 <= hitData_pteaddr;
    end else begin
      lo_lo_3 <= raddr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  REG = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  level = _RAND_2[1:0];
  _RAND_3 = {2{`RANDOM}};
  hitWBStore = _RAND_3[39:0];
  _RAND_4 = {1{`RANDOM}};
  REG_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG_2 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  memRespStore = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  missMaskStore = _RAND_7[17:0];
  _RAND_8 = {1{`RANDOM}};
  raddr = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  alreadyOutFire = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  REG_7 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG_8 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  REG_9 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  hi_hi_hi = _RAND_13[26:0];
  _RAND_14 = {1{`RANDOM}};
  hi_hi_lo = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  hi_lo_4 = _RAND_15[17:0];
  _RAND_16 = {1{`RANDOM}};
  lo_hi_hi = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  lo_hi_lo = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  lo_lo_3 = _RAND_18[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_EmbeddedTLBEmpty_1(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata
);
  assign io_in_ready = io_out_ready; // @[EmbeddedTLB.scala 403:10]
  assign io_out_valid = io_in_valid; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_size = io_in_bits_size; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[EmbeddedTLB.scala 403:10]
endmodule
module ysyx_210000_EmbeddedTLBMD_1(
  input          clock,
  input          reset,
  output [120:0] io_tlbmd_0,
  output [120:0] io_tlbmd_1,
  output [120:0] io_tlbmd_2,
  output [120:0] io_tlbmd_3,
  input          io_write_wen,
  input  [3:0]   io_write_windex,
  input  [3:0]   io_write_waymask,
  input  [120:0] io_write_wdata,
  input  [3:0]   io_rindex,
  output         io_ready
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [120:0] tlbmd_0 [0:15]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_0_MPORT_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_0_MPORT_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_0_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_0_MPORT_1_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0_MPORT_1_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0_MPORT_1_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_1 [0:15]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_1_MPORT_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_1_MPORT_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_1_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_1_MPORT_1_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1_MPORT_1_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1_MPORT_1_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_2 [0:15]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_2_MPORT_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_2_MPORT_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_2_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_2_MPORT_1_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2_MPORT_1_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2_MPORT_1_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_3 [0:15]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_3_MPORT_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_3_MPORT_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_3_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_3_MPORT_1_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3_MPORT_1_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3_MPORT_1_en; // @[EmbeddedTLB.scala 38:18]
  reg  resetState; // @[EmbeddedTLB.scala 42:27]
  reg [3:0] resetSet; // @[Counter.scala 60:40]
  wire  _T = resetSet == 4'hf; // @[Counter.scala 72:24]
  wire [3:0] _T_2 = resetSet + 4'h1; // @[Counter.scala 76:24]
  wire  resetFinish = resetState & _T; // @[Counter.scala 118:17 Counter.scala 118:24]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[EmbeddedTLB.scala 44:22 EmbeddedTLB.scala 44:35 EmbeddedTLB.scala 42:27]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[EmbeddedTLB.scala 53:20]
  assign tlbmd_0_MPORT_addr = io_rindex;
  assign tlbmd_0_MPORT_data = tlbmd_0[tlbmd_0_MPORT_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_0_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_0_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_0_MPORT_1_mask = waymask[0];
  assign tlbmd_0_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_1_MPORT_addr = io_rindex;
  assign tlbmd_1_MPORT_data = tlbmd_1[tlbmd_1_MPORT_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_1_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_1_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_1_MPORT_1_mask = waymask[1];
  assign tlbmd_1_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_2_MPORT_addr = io_rindex;
  assign tlbmd_2_MPORT_data = tlbmd_2[tlbmd_2_MPORT_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_2_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_2_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_2_MPORT_1_mask = waymask[2];
  assign tlbmd_2_MPORT_1_en = resetState | io_write_wen;
  assign tlbmd_3_MPORT_addr = io_rindex;
  assign tlbmd_3_MPORT_data = tlbmd_3[tlbmd_3_MPORT_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_3_MPORT_1_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_3_MPORT_1_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_3_MPORT_1_mask = waymask[3];
  assign tlbmd_3_MPORT_1_en = resetState | io_write_wen;
  assign io_tlbmd_0 = tlbmd_0_MPORT_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_1 = tlbmd_1_MPORT_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_2 = tlbmd_2_MPORT_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_3 = tlbmd_3_MPORT_data; // @[EmbeddedTLB.scala 39:12]
  assign io_ready = ~resetState; // @[EmbeddedTLB.scala 59:15]
  always @(posedge clock) begin
    if(tlbmd_0_MPORT_1_en & tlbmd_0_MPORT_1_mask) begin
      tlbmd_0[tlbmd_0_MPORT_1_addr] <= tlbmd_0_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_1_MPORT_1_en & tlbmd_1_MPORT_1_mask) begin
      tlbmd_1[tlbmd_1_MPORT_1_addr] <= tlbmd_1_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_2_MPORT_1_en & tlbmd_2_MPORT_1_mask) begin
      tlbmd_2[tlbmd_2_MPORT_1_addr] <= tlbmd_2_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_3_MPORT_1_en & tlbmd_3_MPORT_1_mask) begin
      tlbmd_3[tlbmd_3_MPORT_1_addr] <= tlbmd_3_MPORT_1_data; // @[EmbeddedTLB.scala 38:18]
    end
    resetState <= reset | _GEN_2; // @[EmbeddedTLB.scala 42:27 EmbeddedTLB.scala 42:27]
    if (reset) begin // @[Counter.scala 60:40]
      resetSet <= 4'h0; // @[Counter.scala 60:40]
    end else if (resetState) begin // @[Counter.scala 118:17]
      resetSet <= _T_2; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[120:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  resetSet = _RAND_5[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_EmbeddedTLB_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  input         io_mem_resp_valid,
  input  [63:0] io_mem_resp_bits_rdata,
  input  [1:0]  io_csrMMU_priviledgeMode,
  input         io_csrMMU_status_sum,
  input         io_csrMMU_status_mxr,
  output        io_csrMMU_loadPF,
  output        io_csrMMU_storePF,
  output [38:0] io_csrMMU_addr,
  output        _T_28_0,
  input  [63:0] CSRSATP,
  input         amoReq,
  output        vmEnable_0,
  output        _T_27_0,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_reset; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_in_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_in_valid; // @[EmbeddedTLB.scala 80:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [2:0] tlbExec_io_in_bits_size; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_in_bits_cmd; // @[EmbeddedTLB.scala 80:23]
  wire [7:0] tlbExec_io_in_bits_wmask; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_in_bits_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_out_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_out_valid; // @[EmbeddedTLB.scala 80:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [2:0] tlbExec_io_out_bits_size; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_out_bits_cmd; // @[EmbeddedTLB.scala 80:23]
  wire [7:0] tlbExec_io_out_bits_wmask; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_out_bits_wdata; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_0; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_1; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_2; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_3; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mdWrite_windex; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mdReady; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_req_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 80:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_resp_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_resp_valid; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_satp; // @[EmbeddedTLB.scala 80:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_status_sum; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_status_mxr; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 80:23]
  wire [38:0] tlbExec_io_pf_addr; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_isFinish; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_ISAMO; // @[EmbeddedTLB.scala 80:23]
  wire  tlbEmpty_io_in_ready; // @[EmbeddedTLB.scala 81:24]
  wire  tlbEmpty_io_in_valid; // @[EmbeddedTLB.scala 81:24]
  wire [31:0] tlbEmpty_io_in_bits_addr; // @[EmbeddedTLB.scala 81:24]
  wire [2:0] tlbEmpty_io_in_bits_size; // @[EmbeddedTLB.scala 81:24]
  wire [3:0] tlbEmpty_io_in_bits_cmd; // @[EmbeddedTLB.scala 81:24]
  wire [7:0] tlbEmpty_io_in_bits_wmask; // @[EmbeddedTLB.scala 81:24]
  wire [63:0] tlbEmpty_io_in_bits_wdata; // @[EmbeddedTLB.scala 81:24]
  wire  tlbEmpty_io_out_ready; // @[EmbeddedTLB.scala 81:24]
  wire  tlbEmpty_io_out_valid; // @[EmbeddedTLB.scala 81:24]
  wire [31:0] tlbEmpty_io_out_bits_addr; // @[EmbeddedTLB.scala 81:24]
  wire [2:0] tlbEmpty_io_out_bits_size; // @[EmbeddedTLB.scala 81:24]
  wire [3:0] tlbEmpty_io_out_bits_cmd; // @[EmbeddedTLB.scala 81:24]
  wire [7:0] tlbEmpty_io_out_bits_wmask; // @[EmbeddedTLB.scala 81:24]
  wire [63:0] tlbEmpty_io_out_bits_wdata; // @[EmbeddedTLB.scala 81:24]
  wire  mdTLB_clock; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_reset; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_0; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_1; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_2; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_3; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_io_write_wen; // @[EmbeddedTLB.scala 82:21]
  wire [3:0] mdTLB_io_write_windex; // @[EmbeddedTLB.scala 82:21]
  wire [3:0] mdTLB_io_write_waymask; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_write_wdata; // @[EmbeddedTLB.scala 82:21]
  wire [3:0] mdTLB_io_rindex; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_io_ready; // @[EmbeddedTLB.scala 82:21]
  reg [120:0] REG__0; // @[Reg.scala 27:20]
  reg [120:0] REG__1; // @[Reg.scala 27:20]
  reg [120:0] REG__2; // @[Reg.scala 27:20]
  reg [120:0] REG__3; // @[Reg.scala 27:20]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[EmbeddedTLB.scala 114:26]
  wire  vmEnable = CSRSATP[63:60] == 4'h8 & io_csrMMU_priviledgeMode < 2'h3; // @[EmbeddedTLB.scala 102:57]
  reg  REG_1; // @[EmbeddedTLB.scala 105:24]
  wire  _GEN_4 = tlbExec_io_isFinish ? 1'h0 : REG_1; // @[EmbeddedTLB.scala 106:25 EmbeddedTLB.scala 106:33 EmbeddedTLB.scala 105:24]
  wire  _GEN_5 = mdUpdate & vmEnable | _GEN_4; // @[EmbeddedTLB.scala 107:50 EmbeddedTLB.scala 107:58]
  reg [38:0] REG_2_addr; // @[Reg.scala 27:20]
  reg [2:0] REG_2_size; // @[Reg.scala 27:20]
  reg [3:0] REG_2_cmd; // @[Reg.scala 27:20]
  reg [7:0] REG_2_wmask; // @[Reg.scala 27:20]
  reg [63:0] REG_2_wdata; // @[Reg.scala 27:20]
  wire  _T_15 = tlbEmpty_io_out_ready & tlbEmpty_io_out_valid; // @[Decoupled.scala 40:37]
  reg  REG_3; // @[Pipeline.scala 24:24]
  wire  _GEN_12 = _T_15 ? 1'h0 : REG_3; // @[Pipeline.scala 25:25 Pipeline.scala 25:33 Pipeline.scala 24:24]
  wire  _T_16 = tlbExec_io_out_valid & tlbEmpty_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_13 = tlbExec_io_out_valid & tlbEmpty_io_in_ready | _GEN_12; // @[Pipeline.scala 26:38 Pipeline.scala 26:46]
  reg [31:0] REG_4_addr; // @[Reg.scala 27:20]
  reg [2:0] REG_4_size; // @[Reg.scala 27:20]
  reg [3:0] REG_4_cmd; // @[Reg.scala 27:20]
  reg [7:0] REG_4_wmask; // @[Reg.scala 27:20]
  reg [63:0] REG_4_wdata; // @[Reg.scala 27:20]
  wire  _T_21 = tlbExec_io_out_valid & ~tlbExec_io_out_ready; // @[EmbeddedTLB.scala 142:81]
  reg  REG_5; // @[Reg.scala 27:20]
  wire  _GEN_29 = _T_21 | REG_5; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _T_22 = tlbExec_io_out_ready & tlbExec_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_26 = tlbExec_io_pf_loadPF | tlbExec_io_pf_storePF; // @[Bundle.scala 133:23]
  wire  _T_27 = tlbExec_io_out_valid & ~REG_5 | _T_26; // @[EmbeddedTLB.scala 144:65]
  wire  _T_28 = io_csrMMU_loadPF | io_csrMMU_storePF; // @[Bundle.scala 133:23]
  ysyx_210000_EmbeddedTLBExec_1 tlbExec ( // @[EmbeddedTLB.scala 80:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_size(tlbExec_io_in_bits_size),
    .io_in_bits_cmd(tlbExec_io_in_bits_cmd),
    .io_in_bits_wmask(tlbExec_io_in_bits_wmask),
    .io_in_bits_wdata(tlbExec_io_in_bits_wdata),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_size(tlbExec_io_out_bits_size),
    .io_out_bits_cmd(tlbExec_io_out_bits_cmd),
    .io_out_bits_wmask(tlbExec_io_out_bits_wmask),
    .io_out_bits_wdata(tlbExec_io_out_bits_wdata),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_windex(tlbExec_io_mdWrite_windex),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_status_sum(tlbExec_io_pf_status_sum),
    .io_pf_status_mxr(tlbExec_io_pf_status_mxr),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_pf_addr(tlbExec_io_pf_addr),
    .io_isFinish(tlbExec_io_isFinish),
    .ISAMO(tlbExec_ISAMO)
  );
  ysyx_210000_EmbeddedTLBEmpty_1 tlbEmpty ( // @[EmbeddedTLB.scala 81:24]
    .io_in_ready(tlbEmpty_io_in_ready),
    .io_in_valid(tlbEmpty_io_in_valid),
    .io_in_bits_addr(tlbEmpty_io_in_bits_addr),
    .io_in_bits_size(tlbEmpty_io_in_bits_size),
    .io_in_bits_cmd(tlbEmpty_io_in_bits_cmd),
    .io_in_bits_wmask(tlbEmpty_io_in_bits_wmask),
    .io_in_bits_wdata(tlbEmpty_io_in_bits_wdata),
    .io_out_ready(tlbEmpty_io_out_ready),
    .io_out_valid(tlbEmpty_io_out_valid),
    .io_out_bits_addr(tlbEmpty_io_out_bits_addr),
    .io_out_bits_size(tlbEmpty_io_out_bits_size),
    .io_out_bits_cmd(tlbEmpty_io_out_bits_cmd),
    .io_out_bits_wmask(tlbEmpty_io_out_bits_wmask),
    .io_out_bits_wdata(tlbEmpty_io_out_bits_wdata)
  );
  ysyx_210000_EmbeddedTLBMD_1 mdTLB ( // @[EmbeddedTLB.scala 82:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_windex(mdTLB_io_write_windex),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_rindex(mdTLB_io_rindex),
    .io_ready(mdTLB_io_ready)
  );
  assign io_in_req_ready = ~vmEnable ? io_out_req_ready : tlbExec_io_in_ready; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 127:21 EmbeddedTLB.scala 110:16]
  assign io_in_resp_valid = io_out_resp_valid; // @[EmbeddedTLB.scala 138:15]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 138:15]
  assign io_out_req_valid = ~vmEnable ? io_in_req_valid : tlbEmpty_io_out_valid; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 126:22 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_addr = ~vmEnable ? io_in_req_bits_addr[31:0] : tlbEmpty_io_out_bits_addr; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 128:26 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_size = ~vmEnable ? io_in_req_bits_size : tlbEmpty_io_out_bits_size; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 129:26 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_cmd = ~vmEnable ? io_in_req_bits_cmd : tlbEmpty_io_out_bits_cmd; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 130:25 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_wmask = ~vmEnable ? io_in_req_bits_wmask : tlbEmpty_io_out_bits_wmask; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 131:27 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_wdata = ~vmEnable ? io_in_req_bits_wdata : tlbEmpty_io_out_bits_wdata; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 132:27 EmbeddedTLB.scala 135:41]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 87:18]
  assign io_csrMMU_loadPF = tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 88:17]
  assign io_csrMMU_storePF = tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 88:17]
  assign io_csrMMU_addr = tlbExec_io_pf_addr; // @[EmbeddedTLB.scala 88:17]
  assign _T_28_0 = _T_28;
  assign vmEnable_0 = vmEnable;
  assign _T_27_0 = _T_27;
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = REG_1; // @[EmbeddedTLB.scala 112:17]
  assign tlbExec_io_in_bits_addr = REG_2_addr; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_size = REG_2_size; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_cmd = REG_2_cmd; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_wmask = REG_2_wmask; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_wdata = REG_2_wdata; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_out_ready = ~vmEnable | tlbEmpty_io_in_ready; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 124:26 Pipeline.scala 29:16]
  assign tlbExec_io_md_0 = REG__0; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_1 = REG__1; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_2 = REG__2; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_3 = REG__3; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[EmbeddedTLB.scala 90:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_satp = CSRSATP; // @[EmbeddedTLB.scala 86:19]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 88:17]
  assign tlbExec_io_pf_status_sum = io_csrMMU_status_sum; // @[EmbeddedTLB.scala 88:17]
  assign tlbExec_io_pf_status_mxr = io_csrMMU_status_mxr; // @[EmbeddedTLB.scala 88:17]
  assign tlbExec_ISAMO = amoReq;
  assign tlbEmpty_io_in_valid = REG_3; // @[Pipeline.scala 31:17]
  assign tlbEmpty_io_in_bits_addr = REG_4_addr; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_size = REG_4_size; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_cmd = REG_4_cmd; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wmask = REG_4_wmask; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wdata = REG_4_wdata; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_out_ready = ~vmEnable | io_out_req_ready; // @[EmbeddedTLB.scala 123:19 EmbeddedTLB.scala 125:52 EmbeddedTLB.scala 135:41]
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[EmbeddedTLB.scala 99:31]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_windex = tlbExec_io_mdWrite_windex; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_rindex = io_in_req_bits_addr[15:12]; // @[TLB.scala 200:19]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      REG__0 <= 121'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG__0 <= mdTLB_io_tlbmd_0; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG__1 <= 121'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG__1 <= mdTLB_io_tlbmd_1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG__2 <= 121'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG__2 <= mdTLB_io_tlbmd_2; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG__3 <= 121'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG__3 <= mdTLB_io_tlbmd_3; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[EmbeddedTLB.scala 105:24]
      REG_1 <= 1'h0; // @[EmbeddedTLB.scala 105:24]
    end else begin
      REG_1 <= _GEN_5;
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_2_addr <= 39'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG_2_addr <= io_in_req_bits_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_2_size <= 3'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG_2_size <= io_in_req_bits_size; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_2_cmd <= 4'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG_2_cmd <= io_in_req_bits_cmd; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_2_wmask <= 8'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG_2_wmask <= io_in_req_bits_wmask; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_2_wdata <= 64'h0; // @[Reg.scala 27:20]
    end else if (mdUpdate) begin // @[Reg.scala 28:19]
      REG_2_wdata <= io_in_req_bits_wdata; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Pipeline.scala 24:24]
      REG_3 <= 1'h0; // @[Pipeline.scala 24:24]
    end else begin
      REG_3 <= _GEN_13;
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_4_addr <= 32'h0; // @[Reg.scala 27:20]
    end else if (_T_16) begin // @[Reg.scala 28:19]
      REG_4_addr <= tlbExec_io_out_bits_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_4_size <= 3'h0; // @[Reg.scala 27:20]
    end else if (_T_16) begin // @[Reg.scala 28:19]
      REG_4_size <= tlbExec_io_out_bits_size; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_4_cmd <= 4'h0; // @[Reg.scala 27:20]
    end else if (_T_16) begin // @[Reg.scala 28:19]
      REG_4_cmd <= tlbExec_io_out_bits_cmd; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_4_wmask <= 8'h0; // @[Reg.scala 27:20]
    end else if (_T_16) begin // @[Reg.scala 28:19]
      REG_4_wmask <= tlbExec_io_out_bits_wmask; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_4_wdata <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_16) begin // @[Reg.scala 28:19]
      REG_4_wdata <= tlbExec_io_out_bits_wdata; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_5 <= 1'h0; // @[Reg.scala 27:20]
    end else if (REG_5 & _T_22) begin // @[EmbeddedTLB.scala 143:53]
      REG_5 <= 1'h0; // @[EmbeddedTLB.scala 143:72]
    end else begin
      REG_5 <= _GEN_29;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  REG__0 = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  REG__1 = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  REG__2 = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  REG__3 = _RAND_3[120:0];
  _RAND_4 = {1{`RANDOM}};
  REG_1 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  REG_2_addr = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  REG_2_size = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  REG_2_cmd = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  REG_2_wmask = _RAND_8[7:0];
  _RAND_9 = {2{`RANDOM}};
  REG_2_wdata = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  REG_3 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG_4_addr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  REG_4_size = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  REG_4_cmd = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  REG_4_wmask = _RAND_14[7:0];
  _RAND_15 = {2{`RANDOM}};
  REG_4_wdata = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  REG_5 = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_CacheStage1_1(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  input         io_metaReadBus_req_ready,
  output        io_metaReadBus_req_valid,
  output [3:0]  io_metaReadBus_req_bits_setIdx,
  input  [21:0] io_metaReadBus_resp_data_0_tag,
  input         io_metaReadBus_resp_data_0_valid,
  input         io_metaReadBus_resp_data_0_dirty,
  input  [21:0] io_metaReadBus_resp_data_1_tag,
  input         io_metaReadBus_resp_data_1_valid,
  input         io_metaReadBus_resp_data_1_dirty,
  input  [21:0] io_metaReadBus_resp_data_2_tag,
  input         io_metaReadBus_resp_data_2_valid,
  input         io_metaReadBus_resp_data_2_dirty,
  input  [21:0] io_metaReadBus_resp_data_3_tag,
  input         io_metaReadBus_resp_data_3_valid,
  input         io_metaReadBus_resp_data_3_dirty,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [6:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data
);
  wire  _T_20 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = (~io_in_valid | _T_20) & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 134:78]
  assign io_out_valid = io_in_valid & io_metaReadBus_req_ready & io_dataReadBus_req_ready; // @[Cache.scala 133:59]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[Cache.scala 132:19]
  assign io_out_bits_req_size = io_in_bits_size; // @[Cache.scala 132:19]
  assign io_out_bits_req_cmd = io_in_bits_cmd; // @[Cache.scala 132:19]
  assign io_out_bits_req_wmask = io_in_bits_wmask; // @[Cache.scala 132:19]
  assign io_out_bits_req_wdata = io_in_bits_wdata; // @[Cache.scala 132:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 128:34]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[9:6]; // @[Cache.scala 79:45]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[Cache.scala 128:34]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[9:6],io_in_bits_addr[5:3]}; // @[Cat.scala 30:58]
endmodule
module ysyx_210000_CacheStage2_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  output [21:0] io_out_bits_metas_0_tag,
  output        io_out_bits_metas_0_dirty,
  output [21:0] io_out_bits_metas_1_tag,
  output        io_out_bits_metas_1_dirty,
  output [21:0] io_out_bits_metas_2_tag,
  output        io_out_bits_metas_2_dirty,
  output [21:0] io_out_bits_metas_3_tag,
  output        io_out_bits_metas_3_dirty,
  output [63:0] io_out_bits_datas_0_data,
  output [63:0] io_out_bits_datas_1_data,
  output [63:0] io_out_bits_datas_2_data,
  output [63:0] io_out_bits_datas_3_data,
  output        io_out_bits_hit,
  output [3:0]  io_out_bits_waymask,
  output        io_out_bits_mmio,
  output        io_out_bits_isForwardData,
  output [63:0] io_out_bits_forwardData_data_data,
  output [3:0]  io_out_bits_forwardData_waymask,
  input  [21:0] io_metaReadResp_0_tag,
  input         io_metaReadResp_0_valid,
  input         io_metaReadResp_0_dirty,
  input  [21:0] io_metaReadResp_1_tag,
  input         io_metaReadResp_1_valid,
  input         io_metaReadResp_1_dirty,
  input  [21:0] io_metaReadResp_2_tag,
  input         io_metaReadResp_2_valid,
  input         io_metaReadResp_2_dirty,
  input  [21:0] io_metaReadResp_3_tag,
  input         io_metaReadResp_3_valid,
  input         io_metaReadResp_3_dirty,
  input  [63:0] io_dataReadResp_0_data,
  input  [63:0] io_dataReadResp_1_data,
  input  [63:0] io_dataReadResp_2_data,
  input  [63:0] io_dataReadResp_3_data,
  input         io_metaWriteBus_req_valid,
  input  [3:0]  io_metaWriteBus_req_bits_setIdx,
  input  [21:0] io_metaWriteBus_req_bits_data_tag,
  input         io_metaWriteBus_req_bits_data_dirty,
  input  [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_dataWriteBus_req_valid,
  input  [6:0]  io_dataWriteBus_req_bits_setIdx,
  input  [63:0] io_dataWriteBus_req_bits_data_data,
  input  [3:0]  io_dataWriteBus_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 162:31]
  wire [3:0] addr_index = io_in_bits_req_addr[9:6]; // @[Cache.scala 162:31]
  wire [21:0] addr_tag = io_in_bits_req_addr[31:10]; // @[Cache.scala 162:31]
  wire  isForwardMeta = io_in_valid & io_metaWriteBus_req_valid & io_metaWriteBus_req_bits_setIdx == addr_index; // @[Cache.scala 164:64]
  reg  isForwardMetaReg; // @[Cache.scala 165:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[Cache.scala 166:24 Cache.scala 166:43 Cache.scala 165:33]
  wire  _T_10 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_11 = ~io_in_valid; // @[Cache.scala 167:25]
  wire  _T_12 = _T_10 | ~io_in_valid; // @[Cache.scala 167:22]
  reg [21:0] forwardMetaReg_data_tag; // @[Reg.scala 27:20]
  reg  forwardMetaReg_data_valid; // @[Reg.scala 27:20]
  reg  forwardMetaReg_data_dirty; // @[Reg.scala 27:20]
  reg [3:0] forwardMetaReg_waymask; // @[Reg.scala 27:20]
  wire [3:0] _GEN_2 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _GEN_3 = isForwardMeta ? io_metaWriteBus_req_bits_data_dirty : forwardMetaReg_data_dirty; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _GEN_4 = isForwardMeta | forwardMetaReg_data_valid; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire [21:0] _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[Cache.scala 171:42]
  wire  forwardWaymask_0 = _GEN_2[0]; // @[Cache.scala 173:61]
  wire  forwardWaymask_1 = _GEN_2[1]; // @[Cache.scala 173:61]
  wire  forwardWaymask_2 = _GEN_2[2]; // @[Cache.scala 173:61]
  wire  forwardWaymask_3 = _GEN_2[3]; // @[Cache.scala 173:61]
  wire [21:0] metaWay_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 175:22]
  wire  metaWay_0_valid = pickForwardMeta & forwardWaymask_0 ? _GEN_4 : io_metaReadResp_0_valid; // @[Cache.scala 175:22]
  wire [21:0] metaWay_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 175:22]
  wire  metaWay_1_valid = pickForwardMeta & forwardWaymask_1 ? _GEN_4 : io_metaReadResp_1_valid; // @[Cache.scala 175:22]
  wire [21:0] metaWay_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 175:22]
  wire  metaWay_2_valid = pickForwardMeta & forwardWaymask_2 ? _GEN_4 : io_metaReadResp_2_valid; // @[Cache.scala 175:22]
  wire [21:0] metaWay_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 175:22]
  wire  metaWay_3_valid = pickForwardMeta & forwardWaymask_3 ? _GEN_4 : io_metaReadResp_3_valid; // @[Cache.scala 175:22]
  wire  _T_23 = metaWay_0_valid & metaWay_0_tag == addr_tag & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_26 = metaWay_1_valid & metaWay_1_tag == addr_tag & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_29 = metaWay_2_valid & metaWay_2_tag == addr_tag & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_32 = metaWay_3_valid & metaWay_3_tag == addr_tag & io_in_valid; // @[Cache.scala 178:73]
  wire [3:0] hitVec = {_T_32,_T_29,_T_26,_T_23}; // @[Cache.scala 178:90]
  reg [63:0] REG; // @[LFSR64.scala 25:23]
  wire  hi_1 = REG[0] ^ REG[1] ^ REG[3] ^ REG[4]; // @[LFSR64.scala 26:43]
  wire [62:0] lo_1 = REG[63:1]; // @[LFSR64.scala 28:51]
  wire [63:0] _T_40 = {hi_1,lo_1}; // @[Cat.scala 30:58]
  wire [3:0] victimWaymask = 4'h1 << REG[1:0]; // @[Cache.scala 179:42]
  wire  _T_43 = ~metaWay_0_valid; // @[Cache.scala 181:45]
  wire  _T_44 = ~metaWay_1_valid; // @[Cache.scala 181:45]
  wire  _T_45 = ~metaWay_2_valid; // @[Cache.scala 181:45]
  wire  _T_46 = ~metaWay_3_valid; // @[Cache.scala 181:45]
  wire [3:0] invalidVec = {_T_46,_T_45,_T_44,_T_43}; // @[Cache.scala 181:56]
  wire  hasInvalidWay = |invalidVec; // @[Cache.scala 182:34]
  wire [1:0] _T_50 = invalidVec >= 4'h2 ? 2'h2 : 2'h1; // @[Cache.scala 185:8]
  wire [2:0] _T_51 = invalidVec >= 4'h4 ? 3'h4 : {{1'd0}, _T_50}; // @[Cache.scala 184:8]
  wire [3:0] refillInvalidWaymask = invalidVec >= 4'h8 ? 4'h8 : {{1'd0}, _T_51}; // @[Cache.scala 183:33]
  wire [3:0] _T_52 = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[Cache.scala 188:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _T_52; // @[Cache.scala 188:20]
  wire [1:0] _T_57 = waymask[0] + waymask[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_59 = waymask[2] + waymask[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_61 = _T_57 + _T_59; // @[Bitwise.scala 47:55]
  wire  _T_63 = _T_61 > 3'h1; // @[Cache.scala 189:26]
  wire  _T_127 = io_in_bits_req_addr < 32'h10000000; // @[NutCore.scala 115:32]
  wire  _T_131 = io_in_bits_req_addr >= 32'h10000000 & io_in_bits_req_addr < 32'h80000000; // @[NutCore.scala 115:24]
  wire [6:0] _T_141 = {addr_index,addr_wordIndex}; // @[Cat.scala 30:58]
  wire  _T_143 = io_dataWriteBus_req_valid & io_dataWriteBus_req_bits_setIdx == _T_141; // @[Cache.scala 205:13]
  wire  isForwardData = io_in_valid & _T_143; // @[Cache.scala 204:35]
  reg  isForwardDataReg; // @[Cache.scala 207:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[Cache.scala 208:24 Cache.scala 208:43 Cache.scala 207:33]
  reg [63:0] forwardDataReg_data_data; // @[Reg.scala 27:20]
  reg [3:0] forwardDataReg_waymask; // @[Reg.scala 27:20]
  wire  _T_150 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = _T_11 | _T_150; // @[Cache.scala 216:31]
  assign io_out_valid = io_in_valid; // @[Cache.scala 215:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[Cache.scala 214:19]
  assign io_out_bits_req_size = io_in_bits_req_size; // @[Cache.scala 214:19]
  assign io_out_bits_req_cmd = io_in_bits_req_cmd; // @[Cache.scala 214:19]
  assign io_out_bits_req_wmask = io_in_bits_req_wmask; // @[Cache.scala 214:19]
  assign io_out_bits_req_wdata = io_in_bits_req_wdata; // @[Cache.scala 214:19]
  assign io_out_bits_metas_0_tag = pickForwardMeta & forwardWaymask_0 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 175:22]
  assign io_out_bits_metas_0_dirty = pickForwardMeta & forwardWaymask_0 ? _GEN_3 : io_metaReadResp_0_dirty; // @[Cache.scala 175:22]
  assign io_out_bits_metas_1_tag = pickForwardMeta & forwardWaymask_1 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 175:22]
  assign io_out_bits_metas_1_dirty = pickForwardMeta & forwardWaymask_1 ? _GEN_3 : io_metaReadResp_1_dirty; // @[Cache.scala 175:22]
  assign io_out_bits_metas_2_tag = pickForwardMeta & forwardWaymask_2 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 175:22]
  assign io_out_bits_metas_2_dirty = pickForwardMeta & forwardWaymask_2 ? _GEN_3 : io_metaReadResp_2_dirty; // @[Cache.scala 175:22]
  assign io_out_bits_metas_3_tag = pickForwardMeta & forwardWaymask_3 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 175:22]
  assign io_out_bits_metas_3_dirty = pickForwardMeta & forwardWaymask_3 ? _GEN_3 : io_metaReadResp_3_dirty; // @[Cache.scala 175:22]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[Cache.scala 201:21]
  assign io_out_bits_hit = io_in_valid & |hitVec; // @[Cache.scala 199:34]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _T_52; // @[Cache.scala 188:20]
  assign io_out_bits_mmio = _T_127 | _T_131; // @[NutCore.scala 116:15]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[Cache.scala 211:49]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data :
    forwardDataReg_data_data; // @[Cache.scala 212:33]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[Cache.scala 212:33]
  always @(posedge clock) begin
    if (reset) begin // @[Cache.scala 165:33]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 165:33]
    end else if (_T_10 | ~io_in_valid) begin // @[Cache.scala 167:39]
      isForwardMetaReg <= 1'h0; // @[Cache.scala 167:58]
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (reset) begin // @[Reg.scala 27:20]
      forwardMetaReg_data_tag <= 22'h0; // @[Reg.scala 27:20]
    end else if (isForwardMeta) begin // @[Reg.scala 28:19]
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      forwardMetaReg_data_valid <= 1'h0; // @[Reg.scala 27:20]
    end else begin
      forwardMetaReg_data_valid <= _GEN_4;
    end
    if (reset) begin // @[Reg.scala 27:20]
      forwardMetaReg_data_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (isForwardMeta) begin // @[Reg.scala 28:19]
      forwardMetaReg_data_dirty <= io_metaWriteBus_req_bits_data_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      forwardMetaReg_waymask <= 4'h0; // @[Reg.scala 27:20]
    end else if (isForwardMeta) begin // @[Reg.scala 28:19]
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[LFSR64.scala 25:23]
      REG <= 64'h1234567887654321; // @[LFSR64.scala 25:23]
    end else if (REG == 64'h0) begin // @[LFSR64.scala 28:18]
      REG <= 64'h1;
    end else begin
      REG <= _T_40;
    end
    if (reset) begin // @[Cache.scala 207:33]
      isForwardDataReg <= 1'h0; // @[Cache.scala 207:33]
    end else if (_T_12) begin // @[Cache.scala 209:39]
      isForwardDataReg <= 1'h0; // @[Cache.scala 209:58]
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (reset) begin // @[Reg.scala 27:20]
      forwardDataReg_data_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (isForwardData) begin // @[Reg.scala 28:19]
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      forwardDataReg_waymask <= 4'h0; // @[Reg.scala 27:20]
    end else if (isForwardData) begin // @[Reg.scala 28:19]
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask; // @[Reg.scala 28:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_in_valid & _T_63) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:196 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[Cache.scala 196:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_valid & _T_63) | reset)) begin
          $fatal; // @[Cache.scala 196:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_data_dirty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_4[3:0];
  _RAND_5 = {2{`RANDOM}};
  REG = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  isForwardDataReg = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_8[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_CacheStage3_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input  [21:0] io_in_bits_metas_0_tag,
  input         io_in_bits_metas_0_dirty,
  input  [21:0] io_in_bits_metas_1_tag,
  input         io_in_bits_metas_1_dirty,
  input  [21:0] io_in_bits_metas_2_tag,
  input         io_in_bits_metas_2_dirty,
  input  [21:0] io_in_bits_metas_3_tag,
  input         io_in_bits_metas_3_dirty,
  input  [63:0] io_in_bits_datas_0_data,
  input  [63:0] io_in_bits_datas_1_data,
  input  [63:0] io_in_bits_datas_2_data,
  input  [63:0] io_in_bits_datas_3_data,
  input         io_in_bits_hit,
  input  [3:0]  io_in_bits_waymask,
  input         io_in_bits_mmio,
  input         io_in_bits_isForwardData,
  input  [63:0] io_in_bits_forwardData_data_data,
  input  [3:0]  io_in_bits_forwardData_waymask,
  input         io_out_ready,
  output        io_out_valid,
  output [3:0]  io_out_bits_cmd,
  output [63:0] io_out_bits_rdata,
  output        io_isFinish,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [6:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  output        io_dataWriteBus_req_valid,
  output [6:0]  io_dataWriteBus_req_bits_setIdx,
  output [63:0] io_dataWriteBus_req_bits_data_data,
  output [3:0]  io_dataWriteBus_req_bits_waymask,
  output        io_metaWriteBus_req_valid,
  output [3:0]  io_metaWriteBus_req_bits_setIdx,
  output [21:0] io_metaWriteBus_req_bits_data_tag,
  output        io_metaWriteBus_req_bits_data_dirty,
  output [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  output        io_mem_resp_ready,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  output        io_mmio_resp_ready,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_cohResp_valid,
  output [3:0]  io_cohResp_bits_cmd,
  output [63:0] io_cohResp_bits_rdata,
  output        io_dataReadRespToL1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 241:28]
  wire [21:0] metaWriteArb_io_in_0_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_0_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_valid; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 241:28]
  wire [21:0] metaWriteArb_io_in_1_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_valid; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 241:28]
  wire [21:0] metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[Cache.scala 241:28]
  wire  dataWriteArb_io_in_0_valid; // @[Cache.scala 242:28]
  wire [6:0] dataWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_in_1_valid; // @[Cache.scala 242:28]
  wire [6:0] dataWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_out_valid; // @[Cache.scala 242:28]
  wire [6:0] dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[Cache.scala 242:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 245:31]
  wire [3:0] addr_index = io_in_bits_req_addr[9:6]; // @[Cache.scala 245:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[Cache.scala 246:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[Cache.scala 247:25]
  wire  miss = io_in_valid & ~io_in_bits_hit; // @[Cache.scala 248:26]
  wire  _T_6 = io_in_bits_req_cmd == 4'h8; // @[SimpleBus.scala 79:23]
  wire  probe = io_in_valid & _T_6; // @[Cache.scala 249:39]
  wire  _T_7 = io_in_bits_req_cmd == 4'h2; // @[SimpleBus.scala 76:27]
  wire  hitReadBurst = hit & _T_7; // @[Cache.scala 250:26]
  wire  meta_dirty = io_in_bits_waymask[0] & io_in_bits_metas_0_dirty | io_in_bits_waymask[1] & io_in_bits_metas_1_dirty
     | io_in_bits_waymask[2] & io_in_bits_metas_2_dirty | io_in_bits_waymask[3] & io_in_bits_metas_3_dirty; // @[Mux.scala 27:72]
  wire [21:0] _T_26 = io_in_bits_waymask[0] ? io_in_bits_metas_0_tag : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_27 = io_in_bits_waymask[1] ? io_in_bits_metas_1_tag : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_28 = io_in_bits_waymask[2] ? io_in_bits_metas_2_tag : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_29 = io_in_bits_waymask[3] ? io_in_bits_metas_3_tag : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_30 = _T_26 | _T_27; // @[Mux.scala 27:72]
  wire [21:0] _T_31 = _T_30 | _T_28; // @[Mux.scala 27:72]
  wire [21:0] meta_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  wire  useForwardData = io_in_bits_isForwardData & io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[Cache.scala 260:49]
  wire [63:0] _T_43 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_44 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_47 = _T_43 | _T_44; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = _T_47 | _T_45; // @[Mux.scala 27:72]
  wire [63:0] _T_49 = _T_48 | _T_46; // @[Mux.scala 27:72]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _T_49; // @[Cache.scala 262:21]
  wire [7:0] lo_lo_lo = io_in_bits_req_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lo_lo_hi = io_in_bits_req_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lo_hi_lo = io_in_bits_req_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lo_hi_hi = io_in_bits_req_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_lo_lo = io_in_bits_req_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_lo_hi = io_in_bits_req_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_hi_lo = io_in_bits_req_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_hi_hi = io_in_bits_req_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_69 = {hi_hi_hi,hi_hi_lo,hi_lo_hi,hi_lo_lo,lo_hi_hi,lo_hi_lo,lo_lo_hi,lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] wordMask = io_in_bits_req_cmd[0] ? _T_69 : 64'h0; // @[Cache.scala 263:21]
  reg [2:0] value; // @[Counter.scala 60:40]
  wire  _T_70 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_71 = io_in_bits_req_cmd == 4'h3; // @[Cache.scala 266:34]
  wire  _T_72 = io_in_bits_req_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_73 = io_in_bits_req_cmd == 4'h3 | _T_72; // @[Cache.scala 266:62]
  wire [2:0] _value_T_1 = value + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_0 = _T_70 & (io_in_bits_req_cmd == 4'h3 | _T_72) ? _value_T_1 : value; // @[Cache.scala 266:85 Counter.scala 76:15 Counter.scala 60:40]
  wire  hitWrite = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 270:22]
  wire [63:0] _T_77 = io_in_bits_req_wdata & wordMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_78 = ~wordMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_79 = dataRead & _T_78; // @[BitUtils.scala 32:36]
  wire [2:0] lo_1 = _T_73 ? value : addr_wordIndex; // @[Cache.scala 273:51]
  wire  metaHitWriteBus_req_valid = hitWrite & ~meta_dirty; // @[Cache.scala 276:22]
  reg [3:0] state; // @[Cache.scala 281:22]
  reg [2:0] value_1; // @[Counter.scala 60:40]
  reg [2:0] value_2; // @[Counter.scala 60:40]
  reg [1:0] state2; // @[Cache.scala 291:23]
  wire  _T_95 = state == 4'h3; // @[Cache.scala 293:39]
  wire  _T_96 = state == 4'h8; // @[Cache.scala 293:66]
  wire [2:0] lo_2 = _T_96 ? value_1 : value_2; // @[Cache.scala 294:33]
  wire  _T_102 = state2 == 2'h1; // @[Cache.scala 295:105]
  reg [63:0] dataWay_0_data; // @[Reg.scala 27:20]
  reg [63:0] dataWay_1_data; // @[Reg.scala 27:20]
  reg [63:0] dataWay_2_data; // @[Reg.scala 27:20]
  reg [63:0] dataWay_3_data; // @[Reg.scala 27:20]
  wire [63:0] _T_107 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_108 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_109 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_110 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_111 = _T_107 | _T_108; // @[Mux.scala 27:72]
  wire [63:0] _T_112 = _T_111 | _T_109; // @[Mux.scala 27:72]
  wire  _T_114 = 2'h0 == state2; // @[Conditional.scala 37:30]
  wire  _T_115 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_116 = 2'h1 == state2; // @[Conditional.scala 37:30]
  wire  _T_117 = 2'h2 == state2; // @[Conditional.scala 37:30]
  wire  _T_118 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_121 = hitReadBurst & io_out_ready; // @[Cache.scala 301:83]
  wire [1:0] _GEN_8 = _T_118 | io_cohResp_valid | hitReadBurst & io_out_ready ? 2'h0 : state2; // @[Cache.scala 301:100 Cache.scala 301:109 Cache.scala 291:23]
  wire [28:0] hi_1 = io_in_bits_req_addr[31:3]; // @[Cache.scala 305:44]
  wire [31:0] raddr = {hi_1,3'h0}; // @[Cat.scala 30:58]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[Cat.scala 30:58]
  wire  _T_123 = state == 4'h1; // @[Cache.scala 309:23]
  wire [2:0] _T_125 = value_2 == 3'h7 ? 3'h7 : 3'h3; // @[Cache.scala 310:8]
  wire [2:0] cmd = state == 4'h1 ? 3'h2 : _T_125; // @[Cache.scala 309:16]
  wire  _T_131 = state2 == 2'h2; // @[Cache.scala 316:89]
  reg  afterFirstRead; // @[Cache.scala 323:31]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_12 = _T_70 | alreadyOutFire; // @[Reg.scala 28:19 Reg.scala 28:23 Reg.scala 27:20]
  wire  _T_137 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_139 = state == 4'h2; // @[Cache.scala 325:70]
  wire  readingFirst = ~afterFirstRead & _T_137 & state == 4'h2; // @[Cache.scala 325:60]
  wire  _T_142 = mmio ? state == 4'h6 : readingFirst; // @[Cache.scala 328:39]
  reg [63:0] inRdataRegDemand; // @[Reg.scala 27:20]
  wire  _T_143 = state == 4'h0; // @[Cache.scala 331:31]
  wire  _T_147 = _T_96 & _T_131; // @[Cache.scala 332:46]
  wire  _T_151 = _T_96 & io_cohResp_valid; // @[Cache.scala 334:49]
  reg [2:0] REG; // @[Counter.scala 60:40]
  wire  _T_152 = REG == 3'h7; // @[Counter.scala 72:24]
  wire [2:0] _T_154 = REG + 3'h1; // @[Counter.scala 76:24]
  wire  releaseLast = _T_151 & _T_152; // @[Counter.scala 118:17 Counter.scala 118:24]
  wire [2:0] _T_156 = releaseLast ? 3'h6 : 3'h0; // @[Cache.scala 335:54]
  wire [3:0] _T_157 = hit ? 4'hc : 4'h8; // @[Cache.scala 336:8]
  wire  respToL1Fire = _T_121 & _T_131; // @[Cache.scala 338:51]
  wire  _T_167 = (_T_143 | _T_147) & hitReadBurst & io_out_ready; // @[Cache.scala 339:112]
  reg [2:0] REG_1; // @[Counter.scala 60:40]
  wire  _T_168 = REG_1 == 3'h7; // @[Counter.scala 72:24]
  wire [2:0] _T_170 = REG_1 + 3'h1; // @[Counter.scala 76:24]
  wire  respToL1Last = _T_167 & _T_168; // @[Counter.scala 118:17 Counter.scala 118:24]
  wire  _T_171 = 4'h0 == state; // @[Conditional.scala 37:30]
  wire [3:0] _T_173 = hit ? 4'h8 : 4'h0; // @[Cache.scala 348:23]
  wire [2:0] _value_T_4 = addr_wordIndex + 3'h1; // @[Cache.scala 353:93]
  wire [2:0] _value_T_5 = addr_wordIndex == 3'h7 ? 3'h0 : _value_T_4; // @[Cache.scala 353:33]
  wire [3:0] _T_180 = meta_dirty ? 4'h3 : 4'h1; // @[Cache.scala 355:42]
  wire [3:0] _T_181 = mmio ? 4'h5 : _T_180; // @[Cache.scala 355:21]
  wire [3:0] _GEN_20 = miss | mmio ? _T_181 : state; // @[Cache.scala 354:49 Cache.scala 355:15 Cache.scala 281:22]
  wire  _T_182 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_183 = io_mmio_req_ready & io_mmio_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_184 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire  _T_185 = io_mmio_resp_ready & io_mmio_resp_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_26 = _T_185 ? 4'h7 : state; // @[Cache.scala 360:50 Cache.scala 360:58 Cache.scala 281:22]
  wire  _T_186 = 4'h8 == state; // @[Conditional.scala 37:30]
  wire [2:0] _value_T_7 = value_1 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_27 = io_cohResp_valid | respToL1Fire ? _value_T_7 : value_1; // @[Cache.scala 363:48 Counter.scala 76:15 Counter.scala 60:40]
  wire [3:0] _GEN_28 = probe & io_cohResp_valid & releaseLast | respToL1Fire & respToL1Last ? 4'h0 : state; // @[Cache.scala 364:88 Cache.scala 364:96 Cache.scala 281:22]
  wire  _T_195 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_29 = _T_118 ? 4'h2 : state; // @[Cache.scala 367:50 Cache.scala 368:13 Cache.scala 281:22]
  wire [2:0] _GEN_30 = _T_118 ? addr_wordIndex : value_1; // @[Cache.scala 367:50 Cache.scala 369:25 Counter.scala 60:40]
  wire  _T_197 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_31 = _T_71 ? 3'h0 : _GEN_0; // @[Cache.scala 376:52 Cache.scala 376:75]
  wire  _T_201 = io_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [3:0] _GEN_32 = _T_201 ? 4'h7 : state; // @[Cache.scala 377:46 Cache.scala 377:54 Cache.scala 281:22]
  wire  _GEN_33 = _T_137 | afterFirstRead; // @[Cache.scala 373:33 Cache.scala 374:24 Cache.scala 323:31]
  wire [2:0] _GEN_34 = _T_137 ? _value_T_7 : value_1; // @[Cache.scala 373:33 Counter.scala 76:15 Counter.scala 60:40]
  wire [2:0] _GEN_35 = _T_137 ? _GEN_31 : _GEN_0; // @[Cache.scala 373:33]
  wire [3:0] _GEN_36 = _T_137 ? _GEN_32 : state; // @[Cache.scala 373:33 Cache.scala 281:22]
  wire  _T_202 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _value_T_11 = value_2 + 3'h1; // @[Counter.scala 76:24]
  wire [2:0] _GEN_37 = _T_118 ? _value_T_11 : value_2; // @[Cache.scala 382:32 Counter.scala 76:15 Counter.scala 60:40]
  wire  _T_205 = io_mem_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire [3:0] _GEN_38 = _T_205 & _T_118 ? 4'h4 : state; // @[Cache.scala 383:65 Cache.scala 383:73 Cache.scala 281:22]
  wire  _T_208 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_39 = _T_137 ? 4'h1 : state; // @[Cache.scala 386:53 Cache.scala 386:61 Cache.scala 281:22]
  wire  _T_210 = 4'h7 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_40 = _GEN_12 ? 4'h0 : state; // @[Cache.scala 387:76 Cache.scala 387:84 Cache.scala 281:22]
  wire [3:0] _GEN_41 = _T_210 ? _GEN_40 : state; // @[Conditional.scala 39:67 Cache.scala 281:22]
  wire [3:0] _GEN_42 = _T_208 ? _GEN_39 : _GEN_41; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_43 = _T_202 ? _GEN_37 : value_2; // @[Conditional.scala 39:67 Counter.scala 60:40]
  wire [3:0] _GEN_44 = _T_202 ? _GEN_38 : _GEN_42; // @[Conditional.scala 39:67]
  wire  _GEN_45 = _T_197 ? _GEN_33 : afterFirstRead; // @[Conditional.scala 39:67 Cache.scala 323:31]
  wire [2:0] _GEN_46 = _T_197 ? _GEN_34 : value_1; // @[Conditional.scala 39:67 Counter.scala 60:40]
  wire [2:0] _GEN_47 = _T_197 ? _GEN_35 : _GEN_0; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_48 = _T_197 ? _GEN_36 : _GEN_44; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_49 = _T_197 ? value_2 : _GEN_43; // @[Conditional.scala 39:67 Counter.scala 60:40]
  wire [3:0] _GEN_50 = _T_195 ? _GEN_29 : _GEN_48; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_51 = _T_195 ? _GEN_30 : _GEN_46; // @[Conditional.scala 39:67]
  wire  _GEN_52 = _T_195 ? afterFirstRead : _GEN_45; // @[Conditional.scala 39:67 Cache.scala 323:31]
  wire [2:0] _GEN_53 = _T_195 ? _GEN_0 : _GEN_47; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_54 = _T_195 ? value_2 : _GEN_49; // @[Conditional.scala 39:67 Counter.scala 60:40]
  wire [2:0] _GEN_55 = _T_186 ? _GEN_27 : _GEN_51; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_56 = _T_186 ? _GEN_28 : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_186 ? afterFirstRead : _GEN_52; // @[Conditional.scala 39:67 Cache.scala 323:31]
  wire [2:0] _GEN_58 = _T_186 ? _GEN_0 : _GEN_53; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_59 = _T_186 ? value_2 : _GEN_54; // @[Conditional.scala 39:67 Counter.scala 60:40]
  wire [63:0] _T_214 = readingFirst ? wordMask : 64'h0; // @[Cache.scala 390:67]
  wire [63:0] _T_215 = io_in_bits_req_wdata & _T_214; // @[BitUtils.scala 32:13]
  wire [63:0] _T_216 = ~_T_214; // @[BitUtils.scala 32:38]
  wire [63:0] _T_217 = io_mem_resp_bits_rdata & _T_216; // @[BitUtils.scala 32:36]
  wire  dataRefillWriteBus_req_valid = _T_139 & _T_137; // @[Cache.scala 392:39]
  wire  metaRefillWriteBus_req_valid = dataRefillWriteBus_req_valid & _T_201; // @[Cache.scala 400:61]
  wire  _T_239 = ~io_in_bits_req_cmd[0] & ~io_in_bits_req_cmd[3]; // @[SimpleBus.scala 73:26]
  wire [2:0] _T_241 = io_in_bits_req_cmd[0] ? 3'h5 : 3'h0; // @[Cache.scala 428:79]
  wire [2:0] _T_242 = _T_239 ? 3'h6 : _T_241; // @[Cache.scala 428:27]
  wire  _T_247 = state == 4'h7; // @[Cache.scala 434:48]
  wire  _T_266 = io_in_bits_req_cmd[0] | mmio ? _T_247 : afterFirstRead & ~alreadyOutFire; // @[Cache.scala 435:45]
  wire  _T_268 = probe ? 1'h0 : hit | _T_266; // @[Cache.scala 435:8]
  wire  _T_275 = miss ? _T_143 : _T_96 & releaseLast; // @[Cache.scala 442:53]
  wire  _T_284 = hit | io_in_bits_req_cmd[0] ? _T_70 : _T_247 & _GEN_12; // @[Cache.scala 443:8]
  ysyx_210000_Arbiter metaWriteArb ( // @[Cache.scala 241:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_dirty(metaWriteArb_io_in_0_bits_data_dirty),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  ysyx_210000_Arbiter_1 dataWriteArb ( // @[Cache.scala 242:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = io_out_ready & (_T_143 & ~hitReadBurst) & ~miss & ~probe; // @[Cache.scala 446:79]
  assign io_out_valid = io_in_valid & _T_268; // @[Cache.scala 433:31]
  assign io_out_bits_cmd = {{1'd0}, _T_242}; // @[Cache.scala 428:27]
  assign io_out_bits_rdata = hit ? dataRead : inRdataRegDemand; // @[Cache.scala 427:29]
  assign io_isFinish = probe ? io_cohResp_valid & _T_275 : _T_284; // @[Cache.scala 442:21]
  assign io_dataReadBus_req_valid = (state == 4'h3 | state == 4'h8) & state2 == 2'h0; // @[Cache.scala 293:81]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,lo_2}; // @[Cat.scala 30:58]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[Cache.scala 397:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 397:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[Cache.scala 397:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[Cache.scala 397:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[Cache.scala 407:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 407:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 407:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 407:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[Cache.scala 407:23]
  assign io_mem_req_valid = _T_123 | _T_95 & state2 == 2'h2; // @[Cache.scala 316:48]
  assign io_mem_req_bits_addr = _T_123 ? raddr : waddr; // @[Cache.scala 311:35]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[Cache.scala 309:16]
  assign io_mem_req_bits_wdata = _T_112 | _T_110; // @[Mux.scala 27:72]
  assign io_mem_resp_ready = 1'h1; // @[Cache.scala 315:21]
  assign io_mmio_req_valid = state == 4'h5; // @[Cache.scala 321:31]
  assign io_mmio_req_bits_addr = io_in_bits_req_addr; // @[Cache.scala 319:20]
  assign io_mmio_req_bits_size = io_in_bits_req_size; // @[Cache.scala 319:20]
  assign io_mmio_req_bits_cmd = io_in_bits_req_cmd; // @[Cache.scala 319:20]
  assign io_mmio_req_bits_wmask = io_in_bits_req_wmask; // @[Cache.scala 319:20]
  assign io_mmio_req_bits_wdata = io_in_bits_req_wdata; // @[Cache.scala 319:20]
  assign io_mmio_resp_ready = 1'h1; // @[Cache.scala 320:22]
  assign io_cohResp_valid = state == 4'h0 & probe | _T_147; // @[Cache.scala 331:53]
  assign io_cohResp_bits_cmd = _T_96 ? {{1'd0}, _T_156} : _T_157; // @[Cache.scala 335:29]
  assign io_cohResp_bits_rdata = _T_112 | _T_110; // @[Mux.scala 27:72]
  assign io_dataReadRespToL1 = hitReadBurst & (_T_143 & io_out_ready | _T_147); // @[Cache.scala 447:39]
  assign metaWriteArb_io_in_0_valid = hitWrite & ~meta_dirty; // @[Cache.scala 276:22]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[9:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_0_bits_data_tag = _T_31 | _T_29; // @[Mux.scala 27:72]
  assign metaWriteArb_io_in_0_bits_data_dirty = 1'h1; // @[Cache.scala 277:16 Cache.scala 97:16]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 275:29 SRAMTemplate.scala 90:24]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_req_valid & _T_201; // @[Cache.scala 400:61]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[9:6]; // @[Cache.scala 79:45]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:10]; // @[Cache.scala 245:31]
  assign metaWriteArb_io_in_1_bits_data_dirty = io_in_bits_req_cmd[0]; // @[SimpleBus.scala 74:22]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 399:32 SRAMTemplate.scala 90:24]
  assign dataWriteArb_io_in_0_valid = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 270:22]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,lo_1}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_0_bits_data_data = _T_77 | _T_79; // @[BitUtils.scala 32:25]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 271:29 SRAMTemplate.scala 90:24]
  assign dataWriteArb_io_in_1_valid = _T_139 & _T_137; // @[Cache.scala 392:39]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,value_1}; // @[Cat.scala 30:58]
  assign dataWriteArb_io_in_1_bits_data_data = _T_215 | _T_217; // @[BitUtils.scala 32:25]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 391:32 SRAMTemplate.scala 90:24]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 60:40]
      value <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_171) begin // @[Conditional.scala 40:58]
      value <= _GEN_0;
    end else if (_T_182) begin // @[Conditional.scala 39:67]
      value <= _GEN_0;
    end else if (_T_184) begin // @[Conditional.scala 39:67]
      value <= _GEN_0;
    end else begin
      value <= _GEN_58;
    end
    if (reset) begin // @[Cache.scala 281:22]
      state <= 4'h0; // @[Cache.scala 281:22]
    end else if (_T_171) begin // @[Conditional.scala 40:58]
      if (probe) begin // @[Cache.scala 346:20]
        if (io_cohResp_valid) begin // @[Cache.scala 347:34]
          state <= _T_173; // @[Cache.scala 348:17]
        end
      end else if (_T_121) begin // @[Cache.scala 351:50]
        state <= 4'h8; // @[Cache.scala 352:15]
      end else begin
        state <= _GEN_20;
      end
    end else if (_T_182) begin // @[Conditional.scala 39:67]
      if (_T_183) begin // @[Cache.scala 359:48]
        state <= 4'h6; // @[Cache.scala 359:56]
      end
    end else if (_T_184) begin // @[Conditional.scala 39:67]
      state <= _GEN_26;
    end else begin
      state <= _GEN_56;
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_171) begin // @[Conditional.scala 40:58]
      if (probe) begin // @[Cache.scala 346:20]
        if (io_cohResp_valid) begin // @[Cache.scala 347:34]
          value_1 <= addr_wordIndex; // @[Cache.scala 349:29]
        end
      end else if (_T_121) begin // @[Cache.scala 351:50]
        value_1 <= _value_T_5; // @[Cache.scala 353:27]
      end
    end else if (!(_T_182)) begin // @[Conditional.scala 39:67]
      if (!(_T_184)) begin // @[Conditional.scala 39:67]
        value_1 <= _GEN_55;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_2 <= 3'h0; // @[Counter.scala 60:40]
    end else if (!(_T_171)) begin // @[Conditional.scala 40:58]
      if (!(_T_182)) begin // @[Conditional.scala 39:67]
        if (!(_T_184)) begin // @[Conditional.scala 39:67]
          value_2 <= _GEN_59;
        end
      end
    end
    if (reset) begin // @[Cache.scala 291:23]
      state2 <= 2'h0; // @[Cache.scala 291:23]
    end else if (_T_114) begin // @[Conditional.scala 40:58]
      if (_T_115) begin // @[Cache.scala 299:53]
        state2 <= 2'h1; // @[Cache.scala 299:62]
      end
    end else if (_T_116) begin // @[Conditional.scala 39:67]
      state2 <= 2'h2; // @[Cache.scala 300:35]
    end else if (_T_117) begin // @[Conditional.scala 39:67]
      state2 <= _GEN_8;
    end
    if (reset) begin // @[Reg.scala 27:20]
      dataWay_0_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_102) begin // @[Reg.scala 28:19]
      dataWay_0_data <= io_dataReadBus_resp_data_0_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      dataWay_1_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_102) begin // @[Reg.scala 28:19]
      dataWay_1_data <= io_dataReadBus_resp_data_1_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      dataWay_2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_102) begin // @[Reg.scala 28:19]
      dataWay_2_data <= io_dataReadBus_resp_data_2_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      dataWay_3_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_102) begin // @[Reg.scala 28:19]
      dataWay_3_data <= io_dataReadBus_resp_data_3_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Cache.scala 323:31]
      afterFirstRead <= 1'h0; // @[Cache.scala 323:31]
    end else if (_T_171) begin // @[Conditional.scala 40:58]
      afterFirstRead <= 1'h0; // @[Cache.scala 343:22]
    end else if (!(_T_182)) begin // @[Conditional.scala 39:67]
      if (!(_T_184)) begin // @[Conditional.scala 39:67]
        afterFirstRead <= _GEN_57;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      alreadyOutFire <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_171) begin // @[Conditional.scala 40:58]
      alreadyOutFire <= 1'h0; // @[Cache.scala 344:22]
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (reset) begin // @[Reg.scala 27:20]
      inRdataRegDemand <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_142) begin // @[Reg.scala 28:19]
      if (mmio) begin // @[Cache.scala 326:39]
        inRdataRegDemand <= io_mmio_resp_bits_rdata;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      REG <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_151) begin // @[Counter.scala 118:17]
      REG <= _T_154; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      REG_1 <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_167) begin // @[Counter.scala 118:17]
      REG_1 <= _T_170; // @[Counter.scala 76:15]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:252 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"
            ); // @[Cache.scala 252:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(mmio & hit) | reset)) begin
          $fatal; // @[Cache.scala 252:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(metaHitWriteBus_req_valid & metaRefillWriteBus_req_valid) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:449 assert(!(metaHitWriteBus.req.valid && metaRefillWriteBus.req.valid))\n"
            ); // @[Cache.scala 449:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(metaHitWriteBus_req_valid & metaRefillWriteBus_req_valid) | reset)) begin
          $fatal; // @[Cache.scala 449:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(hitWrite & dataRefillWriteBus_req_valid) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Cache.scala:450 assert(!(dataHitWriteBus.req.valid && dataRefillWriteBus.req.valid))\n"
            ); // @[Cache.scala 450:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(hitWrite & dataRefillWriteBus_req_valid) | reset)) begin
          $fatal; // @[Cache.scala 450:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  REG = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  REG_1 = _RAND_13[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_Arbiter_9(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [2:0]  io_in_1_bits_size,
  input  [3:0]  io_in_1_bits_cmd,
  input  [7:0]  io_in_1_bits_wmask,
  input  [63:0] io_in_1_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:19]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:19]
  assign io_out_valid = ~grant_1 | io_in_1_valid; // @[Arbiter.scala 135:31]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  assign io_out_bits_size = io_in_0_valid ? 3'h3 : io_in_1_bits_size; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  assign io_out_bits_cmd = io_in_0_valid ? 4'h8 : io_in_1_bits_cmd; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  assign io_out_bits_wmask = io_in_0_valid ? 8'hff : io_in_1_bits_wmask; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
  assign io_out_bits_wdata = io_in_0_valid ? io_in_0_bits_wdata : io_in_1_bits_wdata; // @[Arbiter.scala 126:27 Arbiter.scala 128:19 Arbiter.scala 124:15]
endmodule
module ysyx_210000_Cache_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  output        io_out_coh_req_ready,
  input         io_out_coh_req_valid,
  input  [31:0] io_out_coh_req_bits_addr,
  input  [63:0] io_out_coh_req_bits_wdata,
  output        io_out_coh_resp_valid,
  output [3:0]  io_out_coh_resp_bits_cmd,
  output [63:0] io_out_coh_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
`endif // RANDOMIZE_REG_INIT
  wire  s1_io_in_ready; // @[Cache.scala 476:18]
  wire  s1_io_in_valid; // @[Cache.scala 476:18]
  wire [31:0] s1_io_in_bits_addr; // @[Cache.scala 476:18]
  wire [2:0] s1_io_in_bits_size; // @[Cache.scala 476:18]
  wire [3:0] s1_io_in_bits_cmd; // @[Cache.scala 476:18]
  wire [7:0] s1_io_in_bits_wmask; // @[Cache.scala 476:18]
  wire [63:0] s1_io_in_bits_wdata; // @[Cache.scala 476:18]
  wire  s1_io_out_ready; // @[Cache.scala 476:18]
  wire  s1_io_out_valid; // @[Cache.scala 476:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[Cache.scala 476:18]
  wire [2:0] s1_io_out_bits_req_size; // @[Cache.scala 476:18]
  wire [3:0] s1_io_out_bits_req_cmd; // @[Cache.scala 476:18]
  wire [7:0] s1_io_out_bits_req_wmask; // @[Cache.scala 476:18]
  wire [63:0] s1_io_out_bits_req_wdata; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_req_ready; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_req_valid; // @[Cache.scala 476:18]
  wire [3:0] s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [21:0] s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 476:18]
  wire [21:0] s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 476:18]
  wire [21:0] s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 476:18]
  wire [21:0] s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 476:18]
  wire  s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 476:18]
  wire  s1_io_dataReadBus_req_ready; // @[Cache.scala 476:18]
  wire  s1_io_dataReadBus_req_valid; // @[Cache.scala 476:18]
  wire [6:0] s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 476:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 476:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 476:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 476:18]
  wire  s2_clock; // @[Cache.scala 477:18]
  wire  s2_reset; // @[Cache.scala 477:18]
  wire  s2_io_in_ready; // @[Cache.scala 477:18]
  wire  s2_io_in_valid; // @[Cache.scala 477:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[Cache.scala 477:18]
  wire [2:0] s2_io_in_bits_req_size; // @[Cache.scala 477:18]
  wire [3:0] s2_io_in_bits_req_cmd; // @[Cache.scala 477:18]
  wire [7:0] s2_io_in_bits_req_wmask; // @[Cache.scala 477:18]
  wire [63:0] s2_io_in_bits_req_wdata; // @[Cache.scala 477:18]
  wire  s2_io_out_ready; // @[Cache.scala 477:18]
  wire  s2_io_out_valid; // @[Cache.scala 477:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[Cache.scala 477:18]
  wire [2:0] s2_io_out_bits_req_size; // @[Cache.scala 477:18]
  wire [3:0] s2_io_out_bits_req_cmd; // @[Cache.scala 477:18]
  wire [7:0] s2_io_out_bits_req_wmask; // @[Cache.scala 477:18]
  wire [63:0] s2_io_out_bits_req_wdata; // @[Cache.scala 477:18]
  wire [21:0] s2_io_out_bits_metas_0_tag; // @[Cache.scala 477:18]
  wire  s2_io_out_bits_metas_0_dirty; // @[Cache.scala 477:18]
  wire [21:0] s2_io_out_bits_metas_1_tag; // @[Cache.scala 477:18]
  wire  s2_io_out_bits_metas_1_dirty; // @[Cache.scala 477:18]
  wire [21:0] s2_io_out_bits_metas_2_tag; // @[Cache.scala 477:18]
  wire  s2_io_out_bits_metas_2_dirty; // @[Cache.scala 477:18]
  wire [21:0] s2_io_out_bits_metas_3_tag; // @[Cache.scala 477:18]
  wire  s2_io_out_bits_metas_3_dirty; // @[Cache.scala 477:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[Cache.scala 477:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[Cache.scala 477:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[Cache.scala 477:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[Cache.scala 477:18]
  wire  s2_io_out_bits_hit; // @[Cache.scala 477:18]
  wire [3:0] s2_io_out_bits_waymask; // @[Cache.scala 477:18]
  wire  s2_io_out_bits_mmio; // @[Cache.scala 477:18]
  wire  s2_io_out_bits_isForwardData; // @[Cache.scala 477:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[Cache.scala 477:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[Cache.scala 477:18]
  wire [21:0] s2_io_metaReadResp_0_tag; // @[Cache.scala 477:18]
  wire  s2_io_metaReadResp_0_valid; // @[Cache.scala 477:18]
  wire  s2_io_metaReadResp_0_dirty; // @[Cache.scala 477:18]
  wire [21:0] s2_io_metaReadResp_1_tag; // @[Cache.scala 477:18]
  wire  s2_io_metaReadResp_1_valid; // @[Cache.scala 477:18]
  wire  s2_io_metaReadResp_1_dirty; // @[Cache.scala 477:18]
  wire [21:0] s2_io_metaReadResp_2_tag; // @[Cache.scala 477:18]
  wire  s2_io_metaReadResp_2_valid; // @[Cache.scala 477:18]
  wire  s2_io_metaReadResp_2_dirty; // @[Cache.scala 477:18]
  wire [21:0] s2_io_metaReadResp_3_tag; // @[Cache.scala 477:18]
  wire  s2_io_metaReadResp_3_valid; // @[Cache.scala 477:18]
  wire  s2_io_metaReadResp_3_dirty; // @[Cache.scala 477:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[Cache.scala 477:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[Cache.scala 477:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[Cache.scala 477:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[Cache.scala 477:18]
  wire  s2_io_metaWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [21:0] s2_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 477:18]
  wire  s2_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 477:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s2_io_dataWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [6:0] s2_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 477:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_clock; // @[Cache.scala 478:18]
  wire  s3_reset; // @[Cache.scala 478:18]
  wire  s3_io_in_ready; // @[Cache.scala 478:18]
  wire  s3_io_in_valid; // @[Cache.scala 478:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[Cache.scala 478:18]
  wire [2:0] s3_io_in_bits_req_size; // @[Cache.scala 478:18]
  wire [3:0] s3_io_in_bits_req_cmd; // @[Cache.scala 478:18]
  wire [7:0] s3_io_in_bits_req_wmask; // @[Cache.scala 478:18]
  wire [63:0] s3_io_in_bits_req_wdata; // @[Cache.scala 478:18]
  wire [21:0] s3_io_in_bits_metas_0_tag; // @[Cache.scala 478:18]
  wire  s3_io_in_bits_metas_0_dirty; // @[Cache.scala 478:18]
  wire [21:0] s3_io_in_bits_metas_1_tag; // @[Cache.scala 478:18]
  wire  s3_io_in_bits_metas_1_dirty; // @[Cache.scala 478:18]
  wire [21:0] s3_io_in_bits_metas_2_tag; // @[Cache.scala 478:18]
  wire  s3_io_in_bits_metas_2_dirty; // @[Cache.scala 478:18]
  wire [21:0] s3_io_in_bits_metas_3_tag; // @[Cache.scala 478:18]
  wire  s3_io_in_bits_metas_3_dirty; // @[Cache.scala 478:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[Cache.scala 478:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[Cache.scala 478:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[Cache.scala 478:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[Cache.scala 478:18]
  wire  s3_io_in_bits_hit; // @[Cache.scala 478:18]
  wire [3:0] s3_io_in_bits_waymask; // @[Cache.scala 478:18]
  wire  s3_io_in_bits_mmio; // @[Cache.scala 478:18]
  wire  s3_io_in_bits_isForwardData; // @[Cache.scala 478:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[Cache.scala 478:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[Cache.scala 478:18]
  wire  s3_io_out_ready; // @[Cache.scala 478:18]
  wire  s3_io_out_valid; // @[Cache.scala 478:18]
  wire [3:0] s3_io_out_bits_cmd; // @[Cache.scala 478:18]
  wire [63:0] s3_io_out_bits_rdata; // @[Cache.scala 478:18]
  wire  s3_io_isFinish; // @[Cache.scala 478:18]
  wire  s3_io_dataReadBus_req_ready; // @[Cache.scala 478:18]
  wire  s3_io_dataReadBus_req_valid; // @[Cache.scala 478:18]
  wire [6:0] s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 478:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[Cache.scala 478:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[Cache.scala 478:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[Cache.scala 478:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[Cache.scala 478:18]
  wire  s3_io_dataWriteBus_req_valid; // @[Cache.scala 478:18]
  wire [6:0] s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 478:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 478:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 478:18]
  wire  s3_io_metaWriteBus_req_valid; // @[Cache.scala 478:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 478:18]
  wire [21:0] s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 478:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 478:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 478:18]
  wire  s3_io_mem_req_ready; // @[Cache.scala 478:18]
  wire  s3_io_mem_req_valid; // @[Cache.scala 478:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[Cache.scala 478:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[Cache.scala 478:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[Cache.scala 478:18]
  wire  s3_io_mem_resp_ready; // @[Cache.scala 478:18]
  wire  s3_io_mem_resp_valid; // @[Cache.scala 478:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[Cache.scala 478:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[Cache.scala 478:18]
  wire  s3_io_mmio_req_ready; // @[Cache.scala 478:18]
  wire  s3_io_mmio_req_valid; // @[Cache.scala 478:18]
  wire [31:0] s3_io_mmio_req_bits_addr; // @[Cache.scala 478:18]
  wire [2:0] s3_io_mmio_req_bits_size; // @[Cache.scala 478:18]
  wire [3:0] s3_io_mmio_req_bits_cmd; // @[Cache.scala 478:18]
  wire [7:0] s3_io_mmio_req_bits_wmask; // @[Cache.scala 478:18]
  wire [63:0] s3_io_mmio_req_bits_wdata; // @[Cache.scala 478:18]
  wire  s3_io_mmio_resp_ready; // @[Cache.scala 478:18]
  wire  s3_io_mmio_resp_valid; // @[Cache.scala 478:18]
  wire [63:0] s3_io_mmio_resp_bits_rdata; // @[Cache.scala 478:18]
  wire  s3_io_cohResp_valid; // @[Cache.scala 478:18]
  wire [3:0] s3_io_cohResp_bits_cmd; // @[Cache.scala 478:18]
  wire [63:0] s3_io_cohResp_bits_rdata; // @[Cache.scala 478:18]
  wire  s3_io_dataReadRespToL1; // @[Cache.scala 478:18]
  wire  metaArray_clock; // @[Cache.scala 479:25]
  wire  metaArray_reset; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_req_ready; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_req_valid; // @[Cache.scala 479:25]
  wire [3:0] metaArray_io_r0_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [21:0] metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 479:25]
  wire [21:0] metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 479:25]
  wire [21:0] metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 479:25]
  wire [21:0] metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 479:25]
  wire  metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 479:25]
  wire  metaArray_io_wreq_valid; // @[Cache.scala 479:25]
  wire [3:0] metaArray_io_wreq_bits_setIdx; // @[Cache.scala 479:25]
  wire [21:0] metaArray_io_wreq_bits_data_tag; // @[Cache.scala 479:25]
  wire  metaArray_io_wreq_bits_data_dirty; // @[Cache.scala 479:25]
  wire [3:0] metaArray_io_wreq_bits_waymask; // @[Cache.scala 479:25]
  wire  dataArray_clock; // @[Cache.scala 480:25]
  wire  dataArray_reset; // @[Cache.scala 480:25]
  wire  dataArray_io_r0_req_ready; // @[Cache.scala 480:25]
  wire  dataArray_io_r0_req_valid; // @[Cache.scala 480:25]
  wire [6:0] dataArray_io_r0_req_bits_setIdx; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r0_resp_data_0_data; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r0_resp_data_1_data; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r0_resp_data_2_data; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r0_resp_data_3_data; // @[Cache.scala 480:25]
  wire  dataArray_io_r1_req_ready; // @[Cache.scala 480:25]
  wire  dataArray_io_r1_req_valid; // @[Cache.scala 480:25]
  wire [6:0] dataArray_io_r1_req_bits_setIdx; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r1_resp_data_0_data; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r1_resp_data_1_data; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r1_resp_data_2_data; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_r1_resp_data_3_data; // @[Cache.scala 480:25]
  wire  dataArray_io_wreq_valid; // @[Cache.scala 480:25]
  wire [6:0] dataArray_io_wreq_bits_setIdx; // @[Cache.scala 480:25]
  wire [63:0] dataArray_io_wreq_bits_data_data; // @[Cache.scala 480:25]
  wire [3:0] dataArray_io_wreq_bits_waymask; // @[Cache.scala 480:25]
  wire  arb_io_in_0_ready; // @[Cache.scala 489:19]
  wire  arb_io_in_0_valid; // @[Cache.scala 489:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[Cache.scala 489:19]
  wire [63:0] arb_io_in_0_bits_wdata; // @[Cache.scala 489:19]
  wire  arb_io_in_1_ready; // @[Cache.scala 489:19]
  wire  arb_io_in_1_valid; // @[Cache.scala 489:19]
  wire [31:0] arb_io_in_1_bits_addr; // @[Cache.scala 489:19]
  wire [2:0] arb_io_in_1_bits_size; // @[Cache.scala 489:19]
  wire [3:0] arb_io_in_1_bits_cmd; // @[Cache.scala 489:19]
  wire [7:0] arb_io_in_1_bits_wmask; // @[Cache.scala 489:19]
  wire [63:0] arb_io_in_1_bits_wdata; // @[Cache.scala 489:19]
  wire  arb_io_out_ready; // @[Cache.scala 489:19]
  wire  arb_io_out_valid; // @[Cache.scala 489:19]
  wire [31:0] arb_io_out_bits_addr; // @[Cache.scala 489:19]
  wire [2:0] arb_io_out_bits_size; // @[Cache.scala 489:19]
  wire [3:0] arb_io_out_bits_cmd; // @[Cache.scala 489:19]
  wire [7:0] arb_io_out_bits_wmask; // @[Cache.scala 489:19]
  wire [63:0] arb_io_out_bits_wdata; // @[Cache.scala 489:19]
  wire  _T = s2_io_out_ready & s2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : REG; // @[Pipeline.scala 25:25 Pipeline.scala 25:33 Pipeline.scala 24:24]
  wire  _T_2 = s1_io_out_valid & s2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = s1_io_out_valid & s2_io_in_ready | _GEN_0; // @[Pipeline.scala 26:38 Pipeline.scala 26:46]
  reg [31:0] REG_1_req_addr; // @[Reg.scala 27:20]
  reg [2:0] REG_1_req_size; // @[Reg.scala 27:20]
  reg [3:0] REG_1_req_cmd; // @[Reg.scala 27:20]
  reg [7:0] REG_1_req_wmask; // @[Reg.scala 27:20]
  reg [63:0] REG_1_req_wdata; // @[Reg.scala 27:20]
  reg  REG_2; // @[Pipeline.scala 24:24]
  wire  _GEN_8 = s3_io_isFinish ? 1'h0 : REG_2; // @[Pipeline.scala 25:25 Pipeline.scala 25:33 Pipeline.scala 24:24]
  wire  _T_5 = s2_io_out_valid & s3_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_9 = s2_io_out_valid & s3_io_in_ready | _GEN_8; // @[Pipeline.scala 26:38 Pipeline.scala 26:46]
  reg [31:0] REG_3_req_addr; // @[Reg.scala 27:20]
  reg [2:0] REG_3_req_size; // @[Reg.scala 27:20]
  reg [3:0] REG_3_req_cmd; // @[Reg.scala 27:20]
  reg [7:0] REG_3_req_wmask; // @[Reg.scala 27:20]
  reg [63:0] REG_3_req_wdata; // @[Reg.scala 27:20]
  reg [21:0] REG_3_metas_0_tag; // @[Reg.scala 27:20]
  reg  REG_3_metas_0_dirty; // @[Reg.scala 27:20]
  reg [21:0] REG_3_metas_1_tag; // @[Reg.scala 27:20]
  reg  REG_3_metas_1_dirty; // @[Reg.scala 27:20]
  reg [21:0] REG_3_metas_2_tag; // @[Reg.scala 27:20]
  reg  REG_3_metas_2_dirty; // @[Reg.scala 27:20]
  reg [21:0] REG_3_metas_3_tag; // @[Reg.scala 27:20]
  reg  REG_3_metas_3_dirty; // @[Reg.scala 27:20]
  reg [63:0] REG_3_datas_0_data; // @[Reg.scala 27:20]
  reg [63:0] REG_3_datas_1_data; // @[Reg.scala 27:20]
  reg [63:0] REG_3_datas_2_data; // @[Reg.scala 27:20]
  reg [63:0] REG_3_datas_3_data; // @[Reg.scala 27:20]
  reg  REG_3_hit; // @[Reg.scala 27:20]
  reg [3:0] REG_3_waymask; // @[Reg.scala 27:20]
  reg  REG_3_mmio; // @[Reg.scala 27:20]
  reg  REG_3_isForwardData; // @[Reg.scala 27:20]
  reg [63:0] REG_3_forwardData_data_data; // @[Reg.scala 27:20]
  reg [3:0] REG_3_forwardData_waymask; // @[Reg.scala 27:20]
  wire  _T_11 = s3_io_out_bits_cmd == 4'h4; // @[SimpleBus.scala 95:26]
  ysyx_210000_CacheStage1_1 s1 ( // @[Cache.scala 476:18]
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_size(s1_io_in_bits_size),
    .io_in_bits_cmd(s1_io_in_bits_cmd),
    .io_in_bits_wmask(s1_io_in_bits_wmask),
    .io_in_bits_wdata(s1_io_in_bits_wdata),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_size(s1_io_out_bits_req_size),
    .io_out_bits_req_cmd(s1_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s1_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s1_io_out_bits_req_wdata),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_0_dirty(s1_io_metaReadBus_resp_data_0_dirty),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_1_dirty(s1_io_metaReadBus_resp_data_1_dirty),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_2_dirty(s1_io_metaReadBus_resp_data_2_dirty),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_metaReadBus_resp_data_3_dirty(s1_io_metaReadBus_resp_data_3_dirty),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data)
  );
  ysyx_210000_CacheStage2_1 s2 ( // @[Cache.scala 477:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_size(s2_io_in_bits_req_size),
    .io_in_bits_req_cmd(s2_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s2_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s2_io_in_bits_req_wdata),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_size(s2_io_out_bits_req_size),
    .io_out_bits_req_cmd(s2_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s2_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s2_io_out_bits_req_wdata),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_0_dirty(s2_io_out_bits_metas_0_dirty),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_1_dirty(s2_io_out_bits_metas_1_dirty),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_2_dirty(s2_io_out_bits_metas_2_dirty),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_metas_3_dirty(s2_io_out_bits_metas_3_dirty),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_0_dirty(s2_io_metaReadResp_0_dirty),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_1_dirty(s2_io_metaReadResp_1_dirty),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_2_dirty(s2_io_metaReadResp_2_dirty),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_metaReadResp_3_dirty(s2_io_metaReadResp_3_dirty),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s2_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask)
  );
  ysyx_210000_CacheStage3_1 s3 ( // @[Cache.scala 478:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_size(s3_io_in_bits_req_size),
    .io_in_bits_req_cmd(s3_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s3_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s3_io_in_bits_req_wdata),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_0_dirty(s3_io_in_bits_metas_0_dirty),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_1_dirty(s3_io_in_bits_metas_1_dirty),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_2_dirty(s3_io_in_bits_metas_2_dirty),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_metas_3_dirty(s3_io_in_bits_metas_3_dirty),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_ready(s3_io_out_ready),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_cmd(s3_io_out_bits_cmd),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_isFinish(s3_io_isFinish),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_mmio_req_ready(s3_io_mmio_req_ready),
    .io_mmio_req_valid(s3_io_mmio_req_valid),
    .io_mmio_req_bits_addr(s3_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(s3_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(s3_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(s3_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(s3_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(s3_io_mmio_resp_ready),
    .io_mmio_resp_valid(s3_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(s3_io_mmio_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid),
    .io_cohResp_bits_cmd(s3_io_cohResp_bits_cmd),
    .io_cohResp_bits_rdata(s3_io_cohResp_bits_rdata),
    .io_dataReadRespToL1(s3_io_dataReadRespToL1)
  );
  ysyx_210000_SRAMTemplateWithArbiter metaArray ( // @[Cache.scala 479:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r0_req_ready(metaArray_io_r0_req_ready),
    .io_r0_req_valid(metaArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(metaArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_tag(metaArray_io_r0_resp_data_0_tag),
    .io_r0_resp_data_0_valid(metaArray_io_r0_resp_data_0_valid),
    .io_r0_resp_data_0_dirty(metaArray_io_r0_resp_data_0_dirty),
    .io_r0_resp_data_1_tag(metaArray_io_r0_resp_data_1_tag),
    .io_r0_resp_data_1_valid(metaArray_io_r0_resp_data_1_valid),
    .io_r0_resp_data_1_dirty(metaArray_io_r0_resp_data_1_dirty),
    .io_r0_resp_data_2_tag(metaArray_io_r0_resp_data_2_tag),
    .io_r0_resp_data_2_valid(metaArray_io_r0_resp_data_2_valid),
    .io_r0_resp_data_2_dirty(metaArray_io_r0_resp_data_2_dirty),
    .io_r0_resp_data_3_tag(metaArray_io_r0_resp_data_3_tag),
    .io_r0_resp_data_3_valid(metaArray_io_r0_resp_data_3_valid),
    .io_r0_resp_data_3_dirty(metaArray_io_r0_resp_data_3_dirty),
    .io_wreq_valid(metaArray_io_wreq_valid),
    .io_wreq_bits_setIdx(metaArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(metaArray_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(metaArray_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(metaArray_io_wreq_bits_waymask)
  );
  ysyx_210000_SRAMTemplateWithArbiter_1 dataArray ( // @[Cache.scala 480:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r0_req_ready(dataArray_io_r0_req_ready),
    .io_r0_req_valid(dataArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(dataArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_data(dataArray_io_r0_resp_data_0_data),
    .io_r0_resp_data_1_data(dataArray_io_r0_resp_data_1_data),
    .io_r0_resp_data_2_data(dataArray_io_r0_resp_data_2_data),
    .io_r0_resp_data_3_data(dataArray_io_r0_resp_data_3_data),
    .io_r1_req_ready(dataArray_io_r1_req_ready),
    .io_r1_req_valid(dataArray_io_r1_req_valid),
    .io_r1_req_bits_setIdx(dataArray_io_r1_req_bits_setIdx),
    .io_r1_resp_data_0_data(dataArray_io_r1_resp_data_0_data),
    .io_r1_resp_data_1_data(dataArray_io_r1_resp_data_1_data),
    .io_r1_resp_data_2_data(dataArray_io_r1_resp_data_2_data),
    .io_r1_resp_data_3_data(dataArray_io_r1_resp_data_3_data),
    .io_wreq_valid(dataArray_io_wreq_valid),
    .io_wreq_bits_setIdx(dataArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(dataArray_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(dataArray_io_wreq_bits_waymask)
  );
  ysyx_210000_Arbiter_9 arb ( // @[Cache.scala 489:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_wdata(arb_io_in_0_bits_wdata),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_size(arb_io_in_1_bits_size),
    .io_in_1_bits_cmd(arb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(arb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(arb_io_in_1_bits_wdata),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_size(arb_io_out_bits_size),
    .io_out_bits_cmd(arb_io_out_bits_cmd),
    .io_out_bits_wmask(arb_io_out_bits_wmask),
    .io_out_bits_wdata(arb_io_out_bits_wdata)
  );
  assign io_in_req_ready = arb_io_in_1_ready; // @[Cache.scala 490:28]
  assign io_in_resp_valid = s3_io_out_valid & _T_11 ? 1'h0 : s3_io_out_valid | s3_io_dataReadRespToL1; // @[Cache.scala 506:26]
  assign io_in_resp_bits_cmd = s3_io_out_bits_cmd; // @[Cache.scala 500:14]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[Cache.scala 500:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[Cache.scala 502:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[Cache.scala 502:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[Cache.scala 502:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[Cache.scala 502:14]
  assign io_out_coh_req_ready = arb_io_in_0_ready; // @[Cache.scala 515:26]
  assign io_out_coh_resp_valid = s3_io_cohResp_valid; // @[Cache.scala 516:21]
  assign io_out_coh_resp_bits_cmd = s3_io_cohResp_bits_cmd; // @[Cache.scala 516:21]
  assign io_out_coh_resp_bits_rdata = s3_io_cohResp_bits_rdata; // @[Cache.scala 516:21]
  assign io_mmio_req_valid = s3_io_mmio_req_valid; // @[Cache.scala 503:11]
  assign io_mmio_req_bits_addr = s3_io_mmio_req_bits_addr; // @[Cache.scala 503:11]
  assign io_mmio_req_bits_size = s3_io_mmio_req_bits_size; // @[Cache.scala 503:11]
  assign io_mmio_req_bits_cmd = s3_io_mmio_req_bits_cmd; // @[Cache.scala 503:11]
  assign io_mmio_req_bits_wmask = s3_io_mmio_req_bits_wmask; // @[Cache.scala 503:11]
  assign io_mmio_req_bits_wdata = s3_io_mmio_req_bits_wdata; // @[Cache.scala 503:11]
  assign s1_io_in_valid = arb_io_out_valid; // @[Cache.scala 492:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[Cache.scala 492:12]
  assign s1_io_in_bits_size = arb_io_out_bits_size; // @[Cache.scala 492:12]
  assign s1_io_in_bits_cmd = arb_io_out_bits_cmd; // @[Cache.scala 492:12]
  assign s1_io_in_bits_wmask = arb_io_out_bits_wmask; // @[Cache.scala 492:12]
  assign s1_io_in_bits_wdata = arb_io_out_bits_wdata; // @[Cache.scala 492:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r0_req_ready; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_0_dirty = metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_1_dirty = metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_2_dirty = metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 524:21]
  assign s1_io_metaReadBus_resp_data_3_dirty = metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r0_req_ready; // @[Cache.scala 525:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r0_resp_data_0_data; // @[Cache.scala 525:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r0_resp_data_1_data; // @[Cache.scala 525:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r0_resp_data_2_data; // @[Cache.scala 525:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r0_resp_data_3_data; // @[Cache.scala 525:21]
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = REG; // @[Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = REG_1_req_addr; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_size = REG_1_req_size; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_cmd = REG_1_req_cmd; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wmask = REG_1_req_wmask; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wdata = REG_1_req_wdata; // @[Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_0_dirty = s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_1_dirty = s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_2_dirty = s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 531:22]
  assign s2_io_metaReadResp_3_dirty = s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 532:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 532:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 532:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 532:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 534:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 534:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 534:22]
  assign s2_io_metaWriteBus_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 534:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 534:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 533:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 533:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 533:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 533:22]
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = REG_2; // @[Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = REG_3_req_addr; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_size = REG_3_req_size; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_cmd = REG_3_req_cmd; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wmask = REG_3_req_wmask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wdata = REG_3_req_wdata; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = REG_3_metas_0_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_dirty = REG_3_metas_0_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = REG_3_metas_1_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_dirty = REG_3_metas_1_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = REG_3_metas_2_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_dirty = REG_3_metas_2_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = REG_3_metas_3_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_dirty = REG_3_metas_3_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = REG_3_datas_0_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = REG_3_datas_1_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = REG_3_datas_2_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = REG_3_datas_3_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = REG_3_hit; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = REG_3_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = REG_3_mmio; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = REG_3_isForwardData; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = REG_3_forwardData_data_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = REG_3_forwardData_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_out_ready = io_in_resp_ready; // @[Cache.scala 500:14]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r1_req_ready; // @[Cache.scala 526:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r1_resp_data_0_data; // @[Cache.scala 526:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r1_resp_data_1_data; // @[Cache.scala 526:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r1_resp_data_2_data; // @[Cache.scala 526:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r1_resp_data_3_data; // @[Cache.scala 526:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[Cache.scala 502:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[Cache.scala 502:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[Cache.scala 502:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[Cache.scala 502:14]
  assign s3_io_mmio_req_ready = io_mmio_req_ready; // @[Cache.scala 503:11]
  assign s3_io_mmio_resp_valid = io_mmio_resp_valid; // @[Cache.scala 503:11]
  assign s3_io_mmio_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[Cache.scala 503:11]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r0_req_valid = s1_io_metaReadBus_req_valid; // @[Cache.scala 524:21]
  assign metaArray_io_r0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 524:21]
  assign metaArray_io_wreq_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 528:18]
  assign metaArray_io_wreq_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 528:18]
  assign metaArray_io_wreq_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 528:18]
  assign metaArray_io_wreq_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 528:18]
  assign metaArray_io_wreq_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 528:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r0_req_valid = s1_io_dataReadBus_req_valid; // @[Cache.scala 525:21]
  assign dataArray_io_r0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 525:21]
  assign dataArray_io_r1_req_valid = s3_io_dataReadBus_req_valid; // @[Cache.scala 526:21]
  assign dataArray_io_r1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 526:21]
  assign dataArray_io_wreq_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 529:18]
  assign dataArray_io_wreq_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 529:18]
  assign dataArray_io_wreq_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 529:18]
  assign dataArray_io_wreq_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 529:18]
  assign arb_io_in_0_valid = io_out_coh_req_valid; // @[Cache.scala 514:24]
  assign arb_io_in_0_bits_addr = io_out_coh_req_bits_addr; // @[Cache.scala 511:19 SimpleBus.scala 64:15]
  assign arb_io_in_0_bits_wdata = io_out_coh_req_bits_wdata; // @[Cache.scala 511:19 SimpleBus.scala 67:16]
  assign arb_io_in_1_valid = io_in_req_valid; // @[Cache.scala 490:28]
  assign arb_io_in_1_bits_addr = io_in_req_bits_addr; // @[Cache.scala 490:28]
  assign arb_io_in_1_bits_size = io_in_req_bits_size; // @[Cache.scala 490:28]
  assign arb_io_in_1_bits_cmd = io_in_req_bits_cmd; // @[Cache.scala 490:28]
  assign arb_io_in_1_bits_wmask = io_in_req_bits_wmask; // @[Cache.scala 490:28]
  assign arb_io_in_1_bits_wdata = io_in_req_bits_wdata; // @[Cache.scala 490:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[Cache.scala 492:12]
  always @(posedge clock) begin
    if (reset) begin // @[Pipeline.scala 24:24]
      REG <= 1'h0; // @[Pipeline.scala 24:24]
    end else begin
      REG <= _GEN_1;
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_req_addr <= 32'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_req_addr <= s1_io_out_bits_req_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_req_size <= 3'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_req_size <= s1_io_out_bits_req_size; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_req_cmd <= 4'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_req_cmd <= s1_io_out_bits_req_cmd; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_req_wmask <= 8'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_req_wmask <= s1_io_out_bits_req_wmask; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_1_req_wdata <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      REG_1_req_wdata <= s1_io_out_bits_req_wdata; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Pipeline.scala 24:24]
      REG_2 <= 1'h0; // @[Pipeline.scala 24:24]
    end else begin
      REG_2 <= _GEN_9;
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_req_addr <= 32'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_req_addr <= s2_io_out_bits_req_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_req_size <= 3'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_req_size <= s2_io_out_bits_req_size; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_req_cmd <= 4'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_req_cmd <= s2_io_out_bits_req_cmd; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_req_wmask <= 8'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_req_wmask <= s2_io_out_bits_req_wmask; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_req_wdata <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_req_wdata <= s2_io_out_bits_req_wdata; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_metas_0_tag <= 22'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_metas_0_tag <= s2_io_out_bits_metas_0_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_metas_0_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_metas_0_dirty <= s2_io_out_bits_metas_0_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_metas_1_tag <= 22'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_metas_1_tag <= s2_io_out_bits_metas_1_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_metas_1_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_metas_1_dirty <= s2_io_out_bits_metas_1_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_metas_2_tag <= 22'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_metas_2_tag <= s2_io_out_bits_metas_2_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_metas_2_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_metas_2_dirty <= s2_io_out_bits_metas_2_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_metas_3_tag <= 22'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_metas_3_tag <= s2_io_out_bits_metas_3_tag; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_metas_3_dirty <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_metas_3_dirty <= s2_io_out_bits_metas_3_dirty; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_datas_0_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_datas_0_data <= s2_io_out_bits_datas_0_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_datas_1_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_datas_1_data <= s2_io_out_bits_datas_1_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_datas_2_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_datas_2_data <= s2_io_out_bits_datas_2_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_datas_3_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_datas_3_data <= s2_io_out_bits_datas_3_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_hit <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_hit <= s2_io_out_bits_hit; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_waymask <= 4'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_waymask <= s2_io_out_bits_waymask; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_mmio <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_mmio <= s2_io_out_bits_mmio; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_isForwardData <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_isForwardData <= s2_io_out_bits_isForwardData; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_forwardData_data_data <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_forwardData_data_data <= s2_io_out_bits_forwardData_data_data; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      REG_3_forwardData_waymask <= 4'h0; // @[Reg.scala 27:20]
    end else if (_T_5) begin // @[Reg.scala 28:19]
      REG_3_forwardData_waymask <= s2_io_out_bits_forwardData_waymask; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1_req_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  REG_1_req_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  REG_1_req_cmd = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  REG_1_req_wmask = _RAND_4[7:0];
  _RAND_5 = {2{`RANDOM}};
  REG_1_req_wdata = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  REG_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  REG_3_req_addr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  REG_3_req_size = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  REG_3_req_cmd = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  REG_3_req_wmask = _RAND_10[7:0];
  _RAND_11 = {2{`RANDOM}};
  REG_3_req_wdata = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  REG_3_metas_0_tag = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  REG_3_metas_0_dirty = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  REG_3_metas_1_tag = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  REG_3_metas_1_dirty = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  REG_3_metas_2_tag = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  REG_3_metas_2_dirty = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  REG_3_metas_3_tag = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  REG_3_metas_3_dirty = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  REG_3_datas_0_data = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  REG_3_datas_1_data = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  REG_3_datas_2_data = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  REG_3_datas_3_data = _RAND_23[63:0];
  _RAND_24 = {1{`RANDOM}};
  REG_3_hit = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  REG_3_waymask = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  REG_3_mmio = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  REG_3_isForwardData = _RAND_27[0:0];
  _RAND_28 = {2{`RANDOM}};
  REG_3_forwardData_data_data = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  REG_3_forwardData_waymask = _RAND_29[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_NutCore(
  input         clock,
  input         reset,
  input         io_imem_mem_req_ready,
  output        io_imem_mem_req_valid,
  output [31:0] io_imem_mem_req_bits_addr,
  output [3:0]  io_imem_mem_req_bits_cmd,
  output [63:0] io_imem_mem_req_bits_wdata,
  input         io_imem_mem_resp_valid,
  input  [3:0]  io_imem_mem_resp_bits_cmd,
  input  [63:0] io_imem_mem_resp_bits_rdata,
  input         io_dmem_mem_req_ready,
  output        io_dmem_mem_req_valid,
  output [31:0] io_dmem_mem_req_bits_addr,
  output [3:0]  io_dmem_mem_req_bits_cmd,
  output [63:0] io_dmem_mem_req_bits_wdata,
  input         io_dmem_mem_resp_valid,
  input  [3:0]  io_dmem_mem_resp_bits_cmd,
  input  [63:0] io_dmem_mem_resp_bits_rdata,
  output        io_dmem_coh_req_ready,
  input         io_dmem_coh_req_valid,
  input  [31:0] io_dmem_coh_req_bits_addr,
  input  [63:0] io_dmem_coh_req_bits_wdata,
  output        io_dmem_coh_resp_valid,
  output [3:0]  io_dmem_coh_resp_bits_cmd,
  output [63:0] io_dmem_coh_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  output        io_mmio_resp_ready,
  input         io_mmio_resp_valid,
  input  [3:0]  io_mmio_resp_bits_cmd,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_frontend_req_ready,
  input         io_frontend_req_valid,
  input  [31:0] io_frontend_req_bits_addr,
  input  [2:0]  io_frontend_req_bits_size,
  input  [3:0]  io_frontend_req_bits_cmd,
  input  [7:0]  io_frontend_req_bits_wmask,
  input  [63:0] io_frontend_req_bits_wdata,
  input         io_frontend_resp_ready,
  output        io_frontend_resp_valid,
  output [3:0]  io_frontend_resp_bits_cmd,
  output [63:0] io_frontend_resp_bits_rdata,
  input         io_extra_mtip,
  input         io_extra_meip_0,
  input         io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
`endif // RANDOMIZE_REG_INIT
  wire  frontend_clock; // @[NutCore.scala 215:34]
  wire  frontend_reset; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_ready; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_valid; // @[NutCore.scala 215:34]
  wire [63:0] frontend_io_out_0_bits_cf_instr; // @[NutCore.scala 215:34]
  wire [38:0] frontend_io_out_0_bits_cf_pc; // @[NutCore.scala 215:34]
  wire [38:0] frontend_io_out_0_bits_cf_pnpc; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_1; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_2; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_12; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_intrVec_0; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_intrVec_1; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_intrVec_2; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_intrVec_3; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_intrVec_4; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_intrVec_5; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_intrVec_6; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_intrVec_7; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_intrVec_8; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_intrVec_9; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_intrVec_10; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_intrVec_11; // @[NutCore.scala 215:34]
  wire [3:0] frontend_io_out_0_bits_cf_brIdx; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_cf_crossPageIPFFix; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_ctrl_src1Type; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_ctrl_src2Type; // @[NutCore.scala 215:34]
  wire [2:0] frontend_io_out_0_bits_ctrl_fuType; // @[NutCore.scala 215:34]
  wire [6:0] frontend_io_out_0_bits_ctrl_fuOpType; // @[NutCore.scala 215:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc1; // @[NutCore.scala 215:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc2; // @[NutCore.scala 215:34]
  wire  frontend_io_out_0_bits_ctrl_rfWen; // @[NutCore.scala 215:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfDest; // @[NutCore.scala 215:34]
  wire [63:0] frontend_io_out_0_bits_data_imm; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_ready; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_valid; // @[NutCore.scala 215:34]
  wire [63:0] frontend_io_out_1_bits_cf_instr; // @[NutCore.scala 215:34]
  wire [38:0] frontend_io_out_1_bits_cf_pc; // @[NutCore.scala 215:34]
  wire [38:0] frontend_io_out_1_bits_cf_pnpc; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_exceptionVec_1; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_exceptionVec_2; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_exceptionVec_12; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_intrVec_0; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_intrVec_1; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_intrVec_2; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_intrVec_3; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_intrVec_4; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_intrVec_5; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_intrVec_6; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_intrVec_7; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_intrVec_8; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_intrVec_9; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_intrVec_10; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_intrVec_11; // @[NutCore.scala 215:34]
  wire [3:0] frontend_io_out_1_bits_cf_brIdx; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_cf_crossPageIPFFix; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_ctrl_src1Type; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_ctrl_src2Type; // @[NutCore.scala 215:34]
  wire [2:0] frontend_io_out_1_bits_ctrl_fuType; // @[NutCore.scala 215:34]
  wire [6:0] frontend_io_out_1_bits_ctrl_fuOpType; // @[NutCore.scala 215:34]
  wire [4:0] frontend_io_out_1_bits_ctrl_rfSrc1; // @[NutCore.scala 215:34]
  wire [4:0] frontend_io_out_1_bits_ctrl_rfSrc2; // @[NutCore.scala 215:34]
  wire  frontend_io_out_1_bits_ctrl_rfWen; // @[NutCore.scala 215:34]
  wire [4:0] frontend_io_out_1_bits_ctrl_rfDest; // @[NutCore.scala 215:34]
  wire [63:0] frontend_io_out_1_bits_data_imm; // @[NutCore.scala 215:34]
  wire  frontend_io_imem_req_ready; // @[NutCore.scala 215:34]
  wire  frontend_io_imem_req_valid; // @[NutCore.scala 215:34]
  wire [38:0] frontend_io_imem_req_bits_addr; // @[NutCore.scala 215:34]
  wire [86:0] frontend_io_imem_req_bits_user; // @[NutCore.scala 215:34]
  wire  frontend_io_imem_resp_ready; // @[NutCore.scala 215:34]
  wire  frontend_io_imem_resp_valid; // @[NutCore.scala 215:34]
  wire [63:0] frontend_io_imem_resp_bits_rdata; // @[NutCore.scala 215:34]
  wire [86:0] frontend_io_imem_resp_bits_user; // @[NutCore.scala 215:34]
  wire [3:0] frontend_io_flushVec; // @[NutCore.scala 215:34]
  wire  frontend_io_ipf; // @[NutCore.scala 215:34]
  wire [38:0] frontend_io_redirect_target; // @[NutCore.scala 215:34]
  wire  frontend_io_redirect_valid; // @[NutCore.scala 215:34]
  wire  frontend_flushICache; // @[NutCore.scala 215:34]
  wire  frontend_REG_6_valid; // @[NutCore.scala 215:34]
  wire [38:0] frontend_REG_6_pc; // @[NutCore.scala 215:34]
  wire  frontend_REG_6_isMissPredict; // @[NutCore.scala 215:34]
  wire [38:0] frontend_REG_6_actualTarget; // @[NutCore.scala 215:34]
  wire  frontend_REG_6_actualTaken; // @[NutCore.scala 215:34]
  wire [6:0] frontend_REG_6_fuOpType; // @[NutCore.scala 215:34]
  wire [1:0] frontend_REG_6_btbType; // @[NutCore.scala 215:34]
  wire  frontend_REG_6_isRVC; // @[NutCore.scala 215:34]
  wire  frontend_vmEnable; // @[NutCore.scala 215:34]
  wire [11:0] frontend_intrVec; // @[NutCore.scala 215:34]
  wire  frontend_flushTLB; // @[NutCore.scala 215:34]
  wire  Backend_inorder_clock; // @[NutCore.scala 257:25]
  wire  Backend_inorder_reset; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_ready; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_valid; // @[NutCore.scala 257:25]
  wire [63:0] Backend_inorder_io_in_0_bits_cf_instr; // @[NutCore.scala 257:25]
  wire [38:0] Backend_inorder_io_in_0_bits_cf_pc; // @[NutCore.scala 257:25]
  wire [38:0] Backend_inorder_io_in_0_bits_cf_pnpc; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_exceptionVec_1; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_exceptionVec_2; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_exceptionVec_12; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_0; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_1; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_2; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_3; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_4; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_5; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_6; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_7; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_8; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_9; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_10; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_11; // @[NutCore.scala 257:25]
  wire [3:0] Backend_inorder_io_in_0_bits_cf_brIdx; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_cf_crossPageIPFFix; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_ctrl_src1Type; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_ctrl_src2Type; // @[NutCore.scala 257:25]
  wire [2:0] Backend_inorder_io_in_0_bits_ctrl_fuType; // @[NutCore.scala 257:25]
  wire [6:0] Backend_inorder_io_in_0_bits_ctrl_fuOpType; // @[NutCore.scala 257:25]
  wire [4:0] Backend_inorder_io_in_0_bits_ctrl_rfSrc1; // @[NutCore.scala 257:25]
  wire [4:0] Backend_inorder_io_in_0_bits_ctrl_rfSrc2; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_in_0_bits_ctrl_rfWen; // @[NutCore.scala 257:25]
  wire [4:0] Backend_inorder_io_in_0_bits_ctrl_rfDest; // @[NutCore.scala 257:25]
  wire [63:0] Backend_inorder_io_in_0_bits_data_imm; // @[NutCore.scala 257:25]
  wire [1:0] Backend_inorder_io_flush; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_dmem_req_ready; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_dmem_req_valid; // @[NutCore.scala 257:25]
  wire [38:0] Backend_inorder_io_dmem_req_bits_addr; // @[NutCore.scala 257:25]
  wire [2:0] Backend_inorder_io_dmem_req_bits_size; // @[NutCore.scala 257:25]
  wire [3:0] Backend_inorder_io_dmem_req_bits_cmd; // @[NutCore.scala 257:25]
  wire [7:0] Backend_inorder_io_dmem_req_bits_wmask; // @[NutCore.scala 257:25]
  wire [63:0] Backend_inorder_io_dmem_req_bits_wdata; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_dmem_resp_valid; // @[NutCore.scala 257:25]
  wire [63:0] Backend_inorder_io_dmem_resp_bits_rdata; // @[NutCore.scala 257:25]
  wire [1:0] Backend_inorder_io_memMMU_imem_priviledgeMode; // @[NutCore.scala 257:25]
  wire [1:0] Backend_inorder_io_memMMU_dmem_priviledgeMode; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_memMMU_dmem_status_sum; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_memMMU_dmem_status_mxr; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_memMMU_dmem_loadPF; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_memMMU_dmem_storePF; // @[NutCore.scala 257:25]
  wire [38:0] Backend_inorder_io_memMMU_dmem_addr; // @[NutCore.scala 257:25]
  wire [38:0] Backend_inorder_io_redirect_target; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_redirect_valid; // @[NutCore.scala 257:25]
  wire  Backend_inorder__T_28; // @[NutCore.scala 257:25]
  wire  Backend_inorder_flushICache; // @[NutCore.scala 257:25]
  wire [63:0] Backend_inorder_satp; // @[NutCore.scala 257:25]
  wire  Backend_inorder_REG_6_valid; // @[NutCore.scala 257:25]
  wire [38:0] Backend_inorder_REG_6_pc; // @[NutCore.scala 257:25]
  wire  Backend_inorder_REG_6_isMissPredict; // @[NutCore.scala 257:25]
  wire [38:0] Backend_inorder_REG_6_actualTarget; // @[NutCore.scala 257:25]
  wire  Backend_inorder_REG_6_actualTaken; // @[NutCore.scala 257:25]
  wire [6:0] Backend_inorder_REG_6_fuOpType; // @[NutCore.scala 257:25]
  wire [1:0] Backend_inorder_REG_6_btbType; // @[NutCore.scala 257:25]
  wire  Backend_inorder_REG_6_isRVC; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_extra_mtip; // @[NutCore.scala 257:25]
  wire  Backend_inorder_amoReq; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_extra_meip_0; // @[NutCore.scala 257:25]
  wire  Backend_inorder_vmEnable; // @[NutCore.scala 257:25]
  wire [11:0] Backend_inorder_intrVec; // @[NutCore.scala 257:25]
  wire  Backend_inorder__T_27; // @[NutCore.scala 257:25]
  wire  Backend_inorder_io_extra_msip; // @[NutCore.scala 257:25]
  wire  Backend_inorder_flushTLB; // @[NutCore.scala 257:25]
  wire  SimpleBusCrossbarNto1_clock; // @[NutCore.scala 261:26]
  wire  SimpleBusCrossbarNto1_reset; // @[NutCore.scala 261:26]
  wire  SimpleBusCrossbarNto1_io_in_0_req_ready; // @[NutCore.scala 261:26]
  wire  SimpleBusCrossbarNto1_io_in_0_req_valid; // @[NutCore.scala 261:26]
  wire [31:0] SimpleBusCrossbarNto1_io_in_0_req_bits_addr; // @[NutCore.scala 261:26]
  wire [2:0] SimpleBusCrossbarNto1_io_in_0_req_bits_size; // @[NutCore.scala 261:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_0_req_bits_cmd; // @[NutCore.scala 261:26]
  wire [7:0] SimpleBusCrossbarNto1_io_in_0_req_bits_wmask; // @[NutCore.scala 261:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_0_req_bits_wdata; // @[NutCore.scala 261:26]
  wire  SimpleBusCrossbarNto1_io_in_0_resp_ready; // @[NutCore.scala 261:26]
  wire  SimpleBusCrossbarNto1_io_in_0_resp_valid; // @[NutCore.scala 261:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_0_resp_bits_cmd; // @[NutCore.scala 261:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata; // @[NutCore.scala 261:26]
  wire  SimpleBusCrossbarNto1_io_in_1_req_ready; // @[NutCore.scala 261:26]
  wire  SimpleBusCrossbarNto1_io_in_1_req_valid; // @[NutCore.scala 261:26]
  wire [31:0] SimpleBusCrossbarNto1_io_in_1_req_bits_addr; // @[NutCore.scala 261:26]
  wire [2:0] SimpleBusCrossbarNto1_io_in_1_req_bits_size; // @[NutCore.scala 261:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_1_req_bits_cmd; // @[NutCore.scala 261:26]
  wire [7:0] SimpleBusCrossbarNto1_io_in_1_req_bits_wmask; // @[NutCore.scala 261:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_1_req_bits_wdata; // @[NutCore.scala 261:26]
  wire  SimpleBusCrossbarNto1_io_in_1_resp_ready; // @[NutCore.scala 261:26]
  wire  SimpleBusCrossbarNto1_io_in_1_resp_valid; // @[NutCore.scala 261:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_1_resp_bits_cmd; // @[NutCore.scala 261:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata; // @[NutCore.scala 261:26]
  wire  SimpleBusCrossbarNto1_io_out_req_ready; // @[NutCore.scala 261:26]
  wire  SimpleBusCrossbarNto1_io_out_req_valid; // @[NutCore.scala 261:26]
  wire [31:0] SimpleBusCrossbarNto1_io_out_req_bits_addr; // @[NutCore.scala 261:26]
  wire [2:0] SimpleBusCrossbarNto1_io_out_req_bits_size; // @[NutCore.scala 261:26]
  wire [3:0] SimpleBusCrossbarNto1_io_out_req_bits_cmd; // @[NutCore.scala 261:26]
  wire [7:0] SimpleBusCrossbarNto1_io_out_req_bits_wmask; // @[NutCore.scala 261:26]
  wire [63:0] SimpleBusCrossbarNto1_io_out_req_bits_wdata; // @[NutCore.scala 261:26]
  wire  SimpleBusCrossbarNto1_io_out_resp_ready; // @[NutCore.scala 261:26]
  wire  SimpleBusCrossbarNto1_io_out_resp_valid; // @[NutCore.scala 261:26]
  wire [3:0] SimpleBusCrossbarNto1_io_out_resp_bits_cmd; // @[NutCore.scala 261:26]
  wire [63:0] SimpleBusCrossbarNto1_io_out_resp_bits_rdata; // @[NutCore.scala 261:26]
  wire  SimpleBusCrossbarNto1_1_clock; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_reset; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_in_0_req_ready; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_in_0_req_valid; // @[NutCore.scala 262:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_addr; // @[NutCore.scala 262:26]
  wire [2:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_size; // @[NutCore.scala 262:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_cmd; // @[NutCore.scala 262:26]
  wire [7:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_wmask; // @[NutCore.scala 262:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_wdata; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_in_0_resp_valid; // @[NutCore.scala 262:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_0_resp_bits_rdata; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_in_1_req_ready; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_in_1_req_valid; // @[NutCore.scala 262:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_1_req_bits_addr; // @[NutCore.scala 262:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_1_req_bits_cmd; // @[NutCore.scala 262:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_1_req_bits_wdata; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_in_1_resp_valid; // @[NutCore.scala 262:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_1_resp_bits_rdata; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_in_2_req_ready; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_in_2_req_valid; // @[NutCore.scala 262:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_2_req_bits_addr; // @[NutCore.scala 262:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_2_req_bits_cmd; // @[NutCore.scala 262:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_2_req_bits_wdata; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_in_2_resp_valid; // @[NutCore.scala 262:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_2_resp_bits_rdata; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_req_ready; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_req_valid; // @[NutCore.scala 262:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_addr; // @[NutCore.scala 262:26]
  wire [2:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_size; // @[NutCore.scala 262:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_cmd; // @[NutCore.scala 262:26]
  wire [7:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_wmask; // @[NutCore.scala 262:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_wdata; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_resp_ready; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_resp_valid; // @[NutCore.scala 262:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_3_resp_bits_cmd; // @[NutCore.scala 262:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_3_resp_bits_rdata; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_out_req_ready; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_out_req_valid; // @[NutCore.scala 262:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_out_req_bits_addr; // @[NutCore.scala 262:26]
  wire [2:0] SimpleBusCrossbarNto1_1_io_out_req_bits_size; // @[NutCore.scala 262:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_out_req_bits_cmd; // @[NutCore.scala 262:26]
  wire [7:0] SimpleBusCrossbarNto1_1_io_out_req_bits_wmask; // @[NutCore.scala 262:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_out_req_bits_wdata; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_out_resp_ready; // @[NutCore.scala 262:26]
  wire  SimpleBusCrossbarNto1_1_io_out_resp_valid; // @[NutCore.scala 262:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_out_resp_bits_cmd; // @[NutCore.scala 262:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_out_resp_bits_rdata; // @[NutCore.scala 262:26]
  wire  MMIOBridge_clock; // @[NutCore.scala 264:28]
  wire  MMIOBridge_reset; // @[NutCore.scala 264:28]
  wire  MMIOBridge_io_in_req_ready; // @[NutCore.scala 264:28]
  wire  MMIOBridge_io_in_req_valid; // @[NutCore.scala 264:28]
  wire [31:0] MMIOBridge_io_in_req_bits_addr; // @[NutCore.scala 264:28]
  wire [2:0] MMIOBridge_io_in_req_bits_size; // @[NutCore.scala 264:28]
  wire  MMIOBridge_io_in_resp_valid; // @[NutCore.scala 264:28]
  wire [63:0] MMIOBridge_io_in_resp_bits_rdata; // @[NutCore.scala 264:28]
  wire  MMIOBridge_io_out_req_ready; // @[NutCore.scala 264:28]
  wire  MMIOBridge_io_out_req_valid; // @[NutCore.scala 264:28]
  wire [31:0] MMIOBridge_io_out_req_bits_addr; // @[NutCore.scala 264:28]
  wire [2:0] MMIOBridge_io_out_req_bits_size; // @[NutCore.scala 264:28]
  wire  MMIOBridge_io_out_resp_ready; // @[NutCore.scala 264:28]
  wire  MMIOBridge_io_out_resp_valid; // @[NutCore.scala 264:28]
  wire [63:0] MMIOBridge_io_out_resp_bits_rdata; // @[NutCore.scala 264:28]
  wire  EmbeddedTLB_clock; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_reset; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_in_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_in_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [38:0] EmbeddedTLB_io_in_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [86:0] EmbeddedTLB_io_in_req_bits_user; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_in_resp_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_in_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire [86:0] EmbeddedTLB_io_in_resp_bits_user; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_out_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_out_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [31:0] EmbeddedTLB_io_out_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [2:0] EmbeddedTLB_io_out_req_bits_size; // @[EmbeddedTLB.scala 427:23]
  wire [86:0] EmbeddedTLB_io_out_req_bits_user; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_out_resp_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_out_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire [86:0] EmbeddedTLB_io_out_resp_bits_user; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_mem_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_mem_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [31:0] EmbeddedTLB_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_mem_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_flush; // @[EmbeddedTLB.scala 427:23]
  wire [1:0] EmbeddedTLB_io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_cacheEmpty; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_ipf; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_CSRSATP; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_MOUFlushTLB; // @[EmbeddedTLB.scala 427:23]
  wire  Cache_clock; // @[Cache.scala 679:35]
  wire  Cache_reset; // @[Cache.scala 679:35]
  wire  Cache_io_in_req_ready; // @[Cache.scala 679:35]
  wire  Cache_io_in_req_valid; // @[Cache.scala 679:35]
  wire [31:0] Cache_io_in_req_bits_addr; // @[Cache.scala 679:35]
  wire [2:0] Cache_io_in_req_bits_size; // @[Cache.scala 679:35]
  wire [86:0] Cache_io_in_req_bits_user; // @[Cache.scala 679:35]
  wire  Cache_io_in_resp_ready; // @[Cache.scala 679:35]
  wire  Cache_io_in_resp_valid; // @[Cache.scala 679:35]
  wire [63:0] Cache_io_in_resp_bits_rdata; // @[Cache.scala 679:35]
  wire [86:0] Cache_io_in_resp_bits_user; // @[Cache.scala 679:35]
  wire [1:0] Cache_io_flush; // @[Cache.scala 679:35]
  wire  Cache_io_out_mem_req_ready; // @[Cache.scala 679:35]
  wire  Cache_io_out_mem_req_valid; // @[Cache.scala 679:35]
  wire [31:0] Cache_io_out_mem_req_bits_addr; // @[Cache.scala 679:35]
  wire [3:0] Cache_io_out_mem_req_bits_cmd; // @[Cache.scala 679:35]
  wire [63:0] Cache_io_out_mem_req_bits_wdata; // @[Cache.scala 679:35]
  wire  Cache_io_out_mem_resp_valid; // @[Cache.scala 679:35]
  wire [3:0] Cache_io_out_mem_resp_bits_cmd; // @[Cache.scala 679:35]
  wire [63:0] Cache_io_out_mem_resp_bits_rdata; // @[Cache.scala 679:35]
  wire  Cache_io_mmio_req_ready; // @[Cache.scala 679:35]
  wire  Cache_io_mmio_req_valid; // @[Cache.scala 679:35]
  wire [31:0] Cache_io_mmio_req_bits_addr; // @[Cache.scala 679:35]
  wire [2:0] Cache_io_mmio_req_bits_size; // @[Cache.scala 679:35]
  wire  Cache_io_mmio_resp_valid; // @[Cache.scala 679:35]
  wire [63:0] Cache_io_mmio_resp_bits_rdata; // @[Cache.scala 679:35]
  wire  Cache_io_empty; // @[Cache.scala 679:35]
  wire  Cache_MOUFlushICache; // @[Cache.scala 679:35]
  wire  EmbeddedTLB_1_clock; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_reset; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_in_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_in_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [38:0] EmbeddedTLB_1_io_in_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [2:0] EmbeddedTLB_1_io_in_req_bits_size; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_1_io_in_req_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [7:0] EmbeddedTLB_1_io_in_req_bits_wmask; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_in_req_bits_wdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_in_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_out_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_out_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [31:0] EmbeddedTLB_1_io_out_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [2:0] EmbeddedTLB_1_io_out_req_bits_size; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_1_io_out_req_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [7:0] EmbeddedTLB_1_io_out_req_bits_wmask; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_out_req_bits_wdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_out_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_mem_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_mem_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [31:0] EmbeddedTLB_1_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_1_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_mem_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire [1:0] EmbeddedTLB_1_io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_csrMMU_status_sum; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_csrMMU_status_mxr; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_csrMMU_loadPF; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_csrMMU_storePF; // @[EmbeddedTLB.scala 427:23]
  wire [38:0] EmbeddedTLB_1_io_csrMMU_addr; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1__T_28_0; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_CSRSATP; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_amoReq; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_vmEnable_0; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1__T_27_0; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_MOUFlushTLB; // @[EmbeddedTLB.scala 427:23]
  wire  Cache_1_clock; // @[Cache.scala 679:35]
  wire  Cache_1_reset; // @[Cache.scala 679:35]
  wire  Cache_1_io_in_req_ready; // @[Cache.scala 679:35]
  wire  Cache_1_io_in_req_valid; // @[Cache.scala 679:35]
  wire [31:0] Cache_1_io_in_req_bits_addr; // @[Cache.scala 679:35]
  wire [2:0] Cache_1_io_in_req_bits_size; // @[Cache.scala 679:35]
  wire [3:0] Cache_1_io_in_req_bits_cmd; // @[Cache.scala 679:35]
  wire [7:0] Cache_1_io_in_req_bits_wmask; // @[Cache.scala 679:35]
  wire [63:0] Cache_1_io_in_req_bits_wdata; // @[Cache.scala 679:35]
  wire  Cache_1_io_in_resp_ready; // @[Cache.scala 679:35]
  wire  Cache_1_io_in_resp_valid; // @[Cache.scala 679:35]
  wire [3:0] Cache_1_io_in_resp_bits_cmd; // @[Cache.scala 679:35]
  wire [63:0] Cache_1_io_in_resp_bits_rdata; // @[Cache.scala 679:35]
  wire  Cache_1_io_out_mem_req_ready; // @[Cache.scala 679:35]
  wire  Cache_1_io_out_mem_req_valid; // @[Cache.scala 679:35]
  wire [31:0] Cache_1_io_out_mem_req_bits_addr; // @[Cache.scala 679:35]
  wire [3:0] Cache_1_io_out_mem_req_bits_cmd; // @[Cache.scala 679:35]
  wire [63:0] Cache_1_io_out_mem_req_bits_wdata; // @[Cache.scala 679:35]
  wire  Cache_1_io_out_mem_resp_valid; // @[Cache.scala 679:35]
  wire [3:0] Cache_1_io_out_mem_resp_bits_cmd; // @[Cache.scala 679:35]
  wire [63:0] Cache_1_io_out_mem_resp_bits_rdata; // @[Cache.scala 679:35]
  wire  Cache_1_io_out_coh_req_ready; // @[Cache.scala 679:35]
  wire  Cache_1_io_out_coh_req_valid; // @[Cache.scala 679:35]
  wire [31:0] Cache_1_io_out_coh_req_bits_addr; // @[Cache.scala 679:35]
  wire [63:0] Cache_1_io_out_coh_req_bits_wdata; // @[Cache.scala 679:35]
  wire  Cache_1_io_out_coh_resp_valid; // @[Cache.scala 679:35]
  wire [3:0] Cache_1_io_out_coh_resp_bits_cmd; // @[Cache.scala 679:35]
  wire [63:0] Cache_1_io_out_coh_resp_bits_rdata; // @[Cache.scala 679:35]
  wire  Cache_1_io_mmio_req_ready; // @[Cache.scala 679:35]
  wire  Cache_1_io_mmio_req_valid; // @[Cache.scala 679:35]
  wire [31:0] Cache_1_io_mmio_req_bits_addr; // @[Cache.scala 679:35]
  wire [2:0] Cache_1_io_mmio_req_bits_size; // @[Cache.scala 679:35]
  wire [3:0] Cache_1_io_mmio_req_bits_cmd; // @[Cache.scala 679:35]
  wire [7:0] Cache_1_io_mmio_req_bits_wmask; // @[Cache.scala 679:35]
  wire [63:0] Cache_1_io_mmio_req_bits_wdata; // @[Cache.scala 679:35]
  wire  Cache_1_io_mmio_resp_valid; // @[Cache.scala 679:35]
  wire [63:0] Cache_1_io_mmio_resp_bits_rdata; // @[Cache.scala 679:35]
  reg [63:0] REG__0_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__0_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__0_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__0_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__0_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg  REG__0_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__0_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__0_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__0_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__0_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__0_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  REG__0_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__0_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__0_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__1_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__1_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__1_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__1_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__1_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg  REG__1_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__1_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__1_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__1_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__1_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__1_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  REG__1_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__1_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__1_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__2_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__2_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__2_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__2_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__2_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg  REG__2_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__2_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__2_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__2_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__2_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__2_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  REG__2_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__2_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__2_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__3_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__3_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] REG__3_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] REG__3_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  REG__3_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg  REG__3_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  REG__3_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] REG__3_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] REG__3_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__3_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__3_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  REG__3_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] REG__3_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg [63:0] REG__3_data_imm; // @[PipelineVector.scala 29:29]
  reg [1:0] REG_1; // @[PipelineVector.scala 30:33]
  reg [1:0] REG_2; // @[PipelineVector.scala 31:33]
  wire [1:0] _T_3 = REG_1 + 2'h1; // @[PipelineVector.scala 33:63]
  wire [1:0] _T_6 = REG_1 + 2'h2; // @[PipelineVector.scala 33:63]
  wire  _T_9 = _T_3 != REG_2 & _T_6 != REG_2; // @[PipelineVector.scala 33:124]
  wire  _WIRE_5_0 = frontend_io_out_0_valid; // @[PipelineVector.scala 36:27 PipelineVector.scala 37:20]
  wire  _WIRE_5_1 = frontend_io_out_1_valid; // @[PipelineVector.scala 36:27 PipelineVector.scala 38:20]
  wire [1:0] _T_10 = _WIRE_5_0 + _WIRE_5_1; // @[PipelineVector.scala 40:46]
  wire  _T_11 = _T_10 >= 2'h1; // @[PipelineVector.scala 41:53]
  wire  _T_12 = _T_10 >= 2'h2; // @[PipelineVector.scala 41:53]
  wire  _T_13 = frontend_io_out_0_ready & frontend_io_out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_14 = frontend_io_out_1_ready & frontend_io_out_1_valid; // @[Decoupled.scala 40:37]
  wire  _T_15 = _T_13 | _T_14; // @[PipelineVector.scala 43:26]
  wire [2:0] _T_16 = {{1'd0}, REG_1}; // @[PipelineVector.scala 45:45]
  wire [63:0] _T_18_cf_instr = _WIRE_5_0 ? frontend_io_out_0_bits_cf_instr : frontend_io_out_1_bits_cf_instr; // @[PipelineVector.scala 45:69]
  wire [38:0] _T_18_cf_pc = _WIRE_5_0 ? frontend_io_out_0_bits_cf_pc : frontend_io_out_1_bits_cf_pc; // @[PipelineVector.scala 45:69]
  wire [38:0] _T_18_cf_pnpc = _WIRE_5_0 ? frontend_io_out_0_bits_cf_pnpc : frontend_io_out_1_bits_cf_pnpc; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_exceptionVec_1 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_exceptionVec_1 :
    frontend_io_out_1_bits_cf_exceptionVec_1; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_exceptionVec_2 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_exceptionVec_2 :
    frontend_io_out_1_bits_cf_exceptionVec_2; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_exceptionVec_12 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_exceptionVec_12 :
    frontend_io_out_1_bits_cf_exceptionVec_12; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_0 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_0 : frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_1 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_1 : frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_2 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_2 : frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_3 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_3 : frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_4 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_4 : frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_5 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_5 : frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_6 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_6 : frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_7 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_7 : frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_8 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_8 : frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_9 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_9 : frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_10 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_10 : frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_intrVec_11 = _WIRE_5_0 ? frontend_io_out_0_bits_cf_intrVec_11 : frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 45:69]
  wire [3:0] _T_18_cf_brIdx = _WIRE_5_0 ? frontend_io_out_0_bits_cf_brIdx : frontend_io_out_1_bits_cf_brIdx; // @[PipelineVector.scala 45:69]
  wire  _T_18_cf_crossPageIPFFix = _WIRE_5_0 ? frontend_io_out_0_bits_cf_crossPageIPFFix :
    frontend_io_out_1_bits_cf_crossPageIPFFix; // @[PipelineVector.scala 45:69]
  wire  _T_18_ctrl_src1Type = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_src1Type : frontend_io_out_1_bits_ctrl_src1Type; // @[PipelineVector.scala 45:69]
  wire  _T_18_ctrl_src2Type = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_src2Type : frontend_io_out_1_bits_ctrl_src2Type; // @[PipelineVector.scala 45:69]
  wire [2:0] _T_18_ctrl_fuType = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_fuType : frontend_io_out_1_bits_ctrl_fuType; // @[PipelineVector.scala 45:69]
  wire [6:0] _T_18_ctrl_fuOpType = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_fuOpType :
    frontend_io_out_1_bits_ctrl_fuOpType; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_18_ctrl_rfSrc1 = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_rfSrc1 : frontend_io_out_1_bits_ctrl_rfSrc1; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_18_ctrl_rfSrc2 = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_rfSrc2 : frontend_io_out_1_bits_ctrl_rfSrc2; // @[PipelineVector.scala 45:69]
  wire  _T_18_ctrl_rfWen = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_rfWen : frontend_io_out_1_bits_ctrl_rfWen; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_18_ctrl_rfDest = _WIRE_5_0 ? frontend_io_out_0_bits_ctrl_rfDest : frontend_io_out_1_bits_ctrl_rfDest; // @[PipelineVector.scala 45:69]
  wire [63:0] _T_18_data_imm = _WIRE_5_0 ? frontend_io_out_0_bits_data_imm : frontend_io_out_1_bits_data_imm; // @[PipelineVector.scala 45:69]
  wire [63:0] _GEN_4 = 2'h0 == _T_16[1:0] ? _T_18_data_imm : REG__0_data_imm; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [63:0] _GEN_5 = 2'h1 == _T_16[1:0] ? _T_18_data_imm : REG__1_data_imm; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [63:0] _GEN_6 = 2'h2 == _T_16[1:0] ? _T_18_data_imm : REG__2_data_imm; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [63:0] _GEN_7 = 2'h3 == _T_16[1:0] ? _T_18_data_imm : REG__3_data_imm; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [4:0] _GEN_48 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_rfDest : REG__0_ctrl_rfDest; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [4:0] _GEN_49 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_rfDest : REG__1_ctrl_rfDest; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [4:0] _GEN_50 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_rfDest : REG__2_ctrl_rfDest; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [4:0] _GEN_51 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_rfDest : REG__3_ctrl_rfDest; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_52 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_rfWen : REG__0_ctrl_rfWen; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_53 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_rfWen : REG__1_ctrl_rfWen; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_54 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_rfWen : REG__2_ctrl_rfWen; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_55 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_rfWen : REG__3_ctrl_rfWen; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [4:0] _GEN_56 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_rfSrc2 : REG__0_ctrl_rfSrc2; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [4:0] _GEN_57 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_rfSrc2 : REG__1_ctrl_rfSrc2; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [4:0] _GEN_58 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_rfSrc2 : REG__2_ctrl_rfSrc2; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [4:0] _GEN_59 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_rfSrc2 : REG__3_ctrl_rfSrc2; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [4:0] _GEN_60 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_rfSrc1 : REG__0_ctrl_rfSrc1; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [4:0] _GEN_61 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_rfSrc1 : REG__1_ctrl_rfSrc1; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [4:0] _GEN_62 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_rfSrc1 : REG__2_ctrl_rfSrc1; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [4:0] _GEN_63 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_rfSrc1 : REG__3_ctrl_rfSrc1; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [6:0] _GEN_64 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_fuOpType : REG__0_ctrl_fuOpType; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [6:0] _GEN_65 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_fuOpType : REG__1_ctrl_fuOpType; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [6:0] _GEN_66 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_fuOpType : REG__2_ctrl_fuOpType; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [6:0] _GEN_67 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_fuOpType : REG__3_ctrl_fuOpType; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [2:0] _GEN_68 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_fuType : REG__0_ctrl_fuType; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [2:0] _GEN_69 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_fuType : REG__1_ctrl_fuType; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [2:0] _GEN_70 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_fuType : REG__2_ctrl_fuType; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [2:0] _GEN_71 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_fuType : REG__3_ctrl_fuType; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_72 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_src2Type : REG__0_ctrl_src2Type; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_73 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_src2Type : REG__1_ctrl_src2Type; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_74 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_src2Type : REG__2_ctrl_src2Type; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_75 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_src2Type : REG__3_ctrl_src2Type; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_76 = 2'h0 == _T_16[1:0] ? _T_18_ctrl_src1Type : REG__0_ctrl_src1Type; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_77 = 2'h1 == _T_16[1:0] ? _T_18_ctrl_src1Type : REG__1_ctrl_src1Type; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_78 = 2'h2 == _T_16[1:0] ? _T_18_ctrl_src1Type : REG__2_ctrl_src1Type; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_79 = 2'h3 == _T_16[1:0] ? _T_18_ctrl_src1Type : REG__3_ctrl_src1Type; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_80 = 2'h0 == _T_16[1:0] ? _T_18_cf_crossPageIPFFix : REG__0_cf_crossPageIPFFix; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_81 = 2'h1 == _T_16[1:0] ? _T_18_cf_crossPageIPFFix : REG__1_cf_crossPageIPFFix; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_82 = 2'h2 == _T_16[1:0] ? _T_18_cf_crossPageIPFFix : REG__2_cf_crossPageIPFFix; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_83 = 2'h3 == _T_16[1:0] ? _T_18_cf_crossPageIPFFix : REG__3_cf_crossPageIPFFix; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [3:0] _GEN_88 = 2'h0 == _T_16[1:0] ? _T_18_cf_brIdx : REG__0_cf_brIdx; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [3:0] _GEN_89 = 2'h1 == _T_16[1:0] ? _T_18_cf_brIdx : REG__1_cf_brIdx; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [3:0] _GEN_90 = 2'h2 == _T_16[1:0] ? _T_18_cf_brIdx : REG__2_cf_brIdx; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [3:0] _GEN_91 = 2'h3 == _T_16[1:0] ? _T_18_cf_brIdx : REG__3_cf_brIdx; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_92 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_0 : REG__0_cf_intrVec_0; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_93 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_0 : REG__1_cf_intrVec_0; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_94 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_0 : REG__2_cf_intrVec_0; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_95 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_0 : REG__3_cf_intrVec_0; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_96 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_1 : REG__0_cf_intrVec_1; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_97 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_1 : REG__1_cf_intrVec_1; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_98 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_1 : REG__2_cf_intrVec_1; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_99 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_1 : REG__3_cf_intrVec_1; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_100 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_2 : REG__0_cf_intrVec_2; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_101 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_2 : REG__1_cf_intrVec_2; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_102 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_2 : REG__2_cf_intrVec_2; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_103 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_2 : REG__3_cf_intrVec_2; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_104 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_3 : REG__0_cf_intrVec_3; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_105 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_3 : REG__1_cf_intrVec_3; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_106 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_3 : REG__2_cf_intrVec_3; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_107 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_3 : REG__3_cf_intrVec_3; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_108 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_4 : REG__0_cf_intrVec_4; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_109 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_4 : REG__1_cf_intrVec_4; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_110 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_4 : REG__2_cf_intrVec_4; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_111 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_4 : REG__3_cf_intrVec_4; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_112 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_5 : REG__0_cf_intrVec_5; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_113 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_5 : REG__1_cf_intrVec_5; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_114 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_5 : REG__2_cf_intrVec_5; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_115 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_5 : REG__3_cf_intrVec_5; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_116 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_6 : REG__0_cf_intrVec_6; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_117 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_6 : REG__1_cf_intrVec_6; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_118 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_6 : REG__2_cf_intrVec_6; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_119 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_6 : REG__3_cf_intrVec_6; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_120 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_7 : REG__0_cf_intrVec_7; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_121 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_7 : REG__1_cf_intrVec_7; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_122 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_7 : REG__2_cf_intrVec_7; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_123 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_7 : REG__3_cf_intrVec_7; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_124 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_8 : REG__0_cf_intrVec_8; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_125 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_8 : REG__1_cf_intrVec_8; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_126 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_8 : REG__2_cf_intrVec_8; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_127 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_8 : REG__3_cf_intrVec_8; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_128 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_9 : REG__0_cf_intrVec_9; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_129 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_9 : REG__1_cf_intrVec_9; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_130 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_9 : REG__2_cf_intrVec_9; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_131 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_9 : REG__3_cf_intrVec_9; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_132 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_10 : REG__0_cf_intrVec_10; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_133 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_10 : REG__1_cf_intrVec_10; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_134 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_10 : REG__2_cf_intrVec_10; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_135 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_10 : REG__3_cf_intrVec_10; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_136 = 2'h0 == _T_16[1:0] ? _T_18_cf_intrVec_11 : REG__0_cf_intrVec_11; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_137 = 2'h1 == _T_16[1:0] ? _T_18_cf_intrVec_11 : REG__1_cf_intrVec_11; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_138 = 2'h2 == _T_16[1:0] ? _T_18_cf_intrVec_11 : REG__2_cf_intrVec_11; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_139 = 2'h3 == _T_16[1:0] ? _T_18_cf_intrVec_11 : REG__3_cf_intrVec_11; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_144 = 2'h0 == _T_16[1:0] ? _T_18_cf_exceptionVec_1 : REG__0_cf_exceptionVec_1; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_145 = 2'h1 == _T_16[1:0] ? _T_18_cf_exceptionVec_1 : REG__1_cf_exceptionVec_1; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_146 = 2'h2 == _T_16[1:0] ? _T_18_cf_exceptionVec_1 : REG__2_cf_exceptionVec_1; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_147 = 2'h3 == _T_16[1:0] ? _T_18_cf_exceptionVec_1 : REG__3_cf_exceptionVec_1; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_148 = 2'h0 == _T_16[1:0] ? _T_18_cf_exceptionVec_2 : REG__0_cf_exceptionVec_2; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_149 = 2'h1 == _T_16[1:0] ? _T_18_cf_exceptionVec_2 : REG__1_cf_exceptionVec_2; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_150 = 2'h2 == _T_16[1:0] ? _T_18_cf_exceptionVec_2 : REG__2_cf_exceptionVec_2; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_151 = 2'h3 == _T_16[1:0] ? _T_18_cf_exceptionVec_2 : REG__3_cf_exceptionVec_2; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_188 = 2'h0 == _T_16[1:0] ? _T_18_cf_exceptionVec_12 : REG__0_cf_exceptionVec_12; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_189 = 2'h1 == _T_16[1:0] ? _T_18_cf_exceptionVec_12 : REG__1_cf_exceptionVec_12; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_190 = 2'h2 == _T_16[1:0] ? _T_18_cf_exceptionVec_12 : REG__2_cf_exceptionVec_12; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire  _GEN_191 = 2'h3 == _T_16[1:0] ? _T_18_cf_exceptionVec_12 : REG__3_cf_exceptionVec_12; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [38:0] _GEN_240 = 2'h0 == _T_16[1:0] ? _T_18_cf_pnpc : REG__0_cf_pnpc; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [38:0] _GEN_241 = 2'h1 == _T_16[1:0] ? _T_18_cf_pnpc : REG__1_cf_pnpc; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [38:0] _GEN_242 = 2'h2 == _T_16[1:0] ? _T_18_cf_pnpc : REG__2_cf_pnpc; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [38:0] _GEN_243 = 2'h3 == _T_16[1:0] ? _T_18_cf_pnpc : REG__3_cf_pnpc; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [38:0] _GEN_244 = 2'h0 == _T_16[1:0] ? _T_18_cf_pc : REG__0_cf_pc; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [38:0] _GEN_245 = 2'h1 == _T_16[1:0] ? _T_18_cf_pc : REG__1_cf_pc; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [38:0] _GEN_246 = 2'h2 == _T_16[1:0] ? _T_18_cf_pc : REG__2_cf_pc; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [38:0] _GEN_247 = 2'h3 == _T_16[1:0] ? _T_18_cf_pc : REG__3_cf_pc; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [63:0] _GEN_248 = 2'h0 == _T_16[1:0] ? _T_18_cf_instr : REG__0_cf_instr; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [63:0] _GEN_249 = 2'h1 == _T_16[1:0] ? _T_18_cf_instr : REG__1_cf_instr; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [63:0] _GEN_250 = 2'h2 == _T_16[1:0] ? _T_18_cf_instr : REG__2_cf_instr; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [63:0] _GEN_251 = 2'h3 == _T_16[1:0] ? _T_18_cf_instr : REG__3_cf_instr; // @[PipelineVector.scala 45:63 PipelineVector.scala 45:63 PipelineVector.scala 29:29]
  wire [63:0] _GEN_256 = _T_11 ? _GEN_4 : REG__0_data_imm; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [63:0] _GEN_257 = _T_11 ? _GEN_5 : REG__1_data_imm; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [63:0] _GEN_258 = _T_11 ? _GEN_6 : REG__2_data_imm; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [63:0] _GEN_259 = _T_11 ? _GEN_7 : REG__3_data_imm; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [4:0] _GEN_300 = _T_11 ? _GEN_48 : REG__0_ctrl_rfDest; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [4:0] _GEN_301 = _T_11 ? _GEN_49 : REG__1_ctrl_rfDest; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [4:0] _GEN_302 = _T_11 ? _GEN_50 : REG__2_ctrl_rfDest; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [4:0] _GEN_303 = _T_11 ? _GEN_51 : REG__3_ctrl_rfDest; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_304 = _T_11 ? _GEN_52 : REG__0_ctrl_rfWen; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_305 = _T_11 ? _GEN_53 : REG__1_ctrl_rfWen; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_306 = _T_11 ? _GEN_54 : REG__2_ctrl_rfWen; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_307 = _T_11 ? _GEN_55 : REG__3_ctrl_rfWen; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [4:0] _GEN_308 = _T_11 ? _GEN_56 : REG__0_ctrl_rfSrc2; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [4:0] _GEN_309 = _T_11 ? _GEN_57 : REG__1_ctrl_rfSrc2; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [4:0] _GEN_310 = _T_11 ? _GEN_58 : REG__2_ctrl_rfSrc2; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [4:0] _GEN_311 = _T_11 ? _GEN_59 : REG__3_ctrl_rfSrc2; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [4:0] _GEN_312 = _T_11 ? _GEN_60 : REG__0_ctrl_rfSrc1; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [4:0] _GEN_313 = _T_11 ? _GEN_61 : REG__1_ctrl_rfSrc1; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [4:0] _GEN_314 = _T_11 ? _GEN_62 : REG__2_ctrl_rfSrc1; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [4:0] _GEN_315 = _T_11 ? _GEN_63 : REG__3_ctrl_rfSrc1; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [6:0] _GEN_316 = _T_11 ? _GEN_64 : REG__0_ctrl_fuOpType; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [6:0] _GEN_317 = _T_11 ? _GEN_65 : REG__1_ctrl_fuOpType; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [6:0] _GEN_318 = _T_11 ? _GEN_66 : REG__2_ctrl_fuOpType; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [6:0] _GEN_319 = _T_11 ? _GEN_67 : REG__3_ctrl_fuOpType; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [2:0] _GEN_320 = _T_11 ? _GEN_68 : REG__0_ctrl_fuType; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [2:0] _GEN_321 = _T_11 ? _GEN_69 : REG__1_ctrl_fuType; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [2:0] _GEN_322 = _T_11 ? _GEN_70 : REG__2_ctrl_fuType; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [2:0] _GEN_323 = _T_11 ? _GEN_71 : REG__3_ctrl_fuType; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_324 = _T_11 ? _GEN_72 : REG__0_ctrl_src2Type; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_325 = _T_11 ? _GEN_73 : REG__1_ctrl_src2Type; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_326 = _T_11 ? _GEN_74 : REG__2_ctrl_src2Type; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_327 = _T_11 ? _GEN_75 : REG__3_ctrl_src2Type; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_328 = _T_11 ? _GEN_76 : REG__0_ctrl_src1Type; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_329 = _T_11 ? _GEN_77 : REG__1_ctrl_src1Type; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_330 = _T_11 ? _GEN_78 : REG__2_ctrl_src1Type; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_331 = _T_11 ? _GEN_79 : REG__3_ctrl_src1Type; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_332 = _T_11 ? _GEN_80 : REG__0_cf_crossPageIPFFix; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_333 = _T_11 ? _GEN_81 : REG__1_cf_crossPageIPFFix; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_334 = _T_11 ? _GEN_82 : REG__2_cf_crossPageIPFFix; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_335 = _T_11 ? _GEN_83 : REG__3_cf_crossPageIPFFix; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [3:0] _GEN_340 = _T_11 ? _GEN_88 : REG__0_cf_brIdx; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [3:0] _GEN_341 = _T_11 ? _GEN_89 : REG__1_cf_brIdx; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [3:0] _GEN_342 = _T_11 ? _GEN_90 : REG__2_cf_brIdx; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [3:0] _GEN_343 = _T_11 ? _GEN_91 : REG__3_cf_brIdx; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_344 = _T_11 ? _GEN_92 : REG__0_cf_intrVec_0; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_345 = _T_11 ? _GEN_93 : REG__1_cf_intrVec_0; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_346 = _T_11 ? _GEN_94 : REG__2_cf_intrVec_0; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_347 = _T_11 ? _GEN_95 : REG__3_cf_intrVec_0; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_348 = _T_11 ? _GEN_96 : REG__0_cf_intrVec_1; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_349 = _T_11 ? _GEN_97 : REG__1_cf_intrVec_1; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_350 = _T_11 ? _GEN_98 : REG__2_cf_intrVec_1; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_351 = _T_11 ? _GEN_99 : REG__3_cf_intrVec_1; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_352 = _T_11 ? _GEN_100 : REG__0_cf_intrVec_2; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_353 = _T_11 ? _GEN_101 : REG__1_cf_intrVec_2; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_354 = _T_11 ? _GEN_102 : REG__2_cf_intrVec_2; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_355 = _T_11 ? _GEN_103 : REG__3_cf_intrVec_2; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_356 = _T_11 ? _GEN_104 : REG__0_cf_intrVec_3; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_357 = _T_11 ? _GEN_105 : REG__1_cf_intrVec_3; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_358 = _T_11 ? _GEN_106 : REG__2_cf_intrVec_3; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_359 = _T_11 ? _GEN_107 : REG__3_cf_intrVec_3; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_360 = _T_11 ? _GEN_108 : REG__0_cf_intrVec_4; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_361 = _T_11 ? _GEN_109 : REG__1_cf_intrVec_4; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_362 = _T_11 ? _GEN_110 : REG__2_cf_intrVec_4; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_363 = _T_11 ? _GEN_111 : REG__3_cf_intrVec_4; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_364 = _T_11 ? _GEN_112 : REG__0_cf_intrVec_5; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_365 = _T_11 ? _GEN_113 : REG__1_cf_intrVec_5; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_366 = _T_11 ? _GEN_114 : REG__2_cf_intrVec_5; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_367 = _T_11 ? _GEN_115 : REG__3_cf_intrVec_5; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_368 = _T_11 ? _GEN_116 : REG__0_cf_intrVec_6; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_369 = _T_11 ? _GEN_117 : REG__1_cf_intrVec_6; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_370 = _T_11 ? _GEN_118 : REG__2_cf_intrVec_6; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_371 = _T_11 ? _GEN_119 : REG__3_cf_intrVec_6; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_372 = _T_11 ? _GEN_120 : REG__0_cf_intrVec_7; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_373 = _T_11 ? _GEN_121 : REG__1_cf_intrVec_7; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_374 = _T_11 ? _GEN_122 : REG__2_cf_intrVec_7; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_375 = _T_11 ? _GEN_123 : REG__3_cf_intrVec_7; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_376 = _T_11 ? _GEN_124 : REG__0_cf_intrVec_8; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_377 = _T_11 ? _GEN_125 : REG__1_cf_intrVec_8; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_378 = _T_11 ? _GEN_126 : REG__2_cf_intrVec_8; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_379 = _T_11 ? _GEN_127 : REG__3_cf_intrVec_8; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_380 = _T_11 ? _GEN_128 : REG__0_cf_intrVec_9; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_381 = _T_11 ? _GEN_129 : REG__1_cf_intrVec_9; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_382 = _T_11 ? _GEN_130 : REG__2_cf_intrVec_9; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_383 = _T_11 ? _GEN_131 : REG__3_cf_intrVec_9; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_384 = _T_11 ? _GEN_132 : REG__0_cf_intrVec_10; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_385 = _T_11 ? _GEN_133 : REG__1_cf_intrVec_10; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_386 = _T_11 ? _GEN_134 : REG__2_cf_intrVec_10; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_387 = _T_11 ? _GEN_135 : REG__3_cf_intrVec_10; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_388 = _T_11 ? _GEN_136 : REG__0_cf_intrVec_11; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_389 = _T_11 ? _GEN_137 : REG__1_cf_intrVec_11; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_390 = _T_11 ? _GEN_138 : REG__2_cf_intrVec_11; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_391 = _T_11 ? _GEN_139 : REG__3_cf_intrVec_11; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_396 = _T_11 ? _GEN_144 : REG__0_cf_exceptionVec_1; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_397 = _T_11 ? _GEN_145 : REG__1_cf_exceptionVec_1; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_398 = _T_11 ? _GEN_146 : REG__2_cf_exceptionVec_1; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_399 = _T_11 ? _GEN_147 : REG__3_cf_exceptionVec_1; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_400 = _T_11 ? _GEN_148 : REG__0_cf_exceptionVec_2; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_401 = _T_11 ? _GEN_149 : REG__1_cf_exceptionVec_2; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_402 = _T_11 ? _GEN_150 : REG__2_cf_exceptionVec_2; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_403 = _T_11 ? _GEN_151 : REG__3_cf_exceptionVec_2; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_440 = _T_11 ? _GEN_188 : REG__0_cf_exceptionVec_12; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_441 = _T_11 ? _GEN_189 : REG__1_cf_exceptionVec_12; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_442 = _T_11 ? _GEN_190 : REG__2_cf_exceptionVec_12; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire  _GEN_443 = _T_11 ? _GEN_191 : REG__3_cf_exceptionVec_12; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [38:0] _GEN_492 = _T_11 ? _GEN_240 : REG__0_cf_pnpc; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [38:0] _GEN_493 = _T_11 ? _GEN_241 : REG__1_cf_pnpc; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [38:0] _GEN_494 = _T_11 ? _GEN_242 : REG__2_cf_pnpc; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [38:0] _GEN_495 = _T_11 ? _GEN_243 : REG__3_cf_pnpc; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [38:0] _GEN_496 = _T_11 ? _GEN_244 : REG__0_cf_pc; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [38:0] _GEN_497 = _T_11 ? _GEN_245 : REG__1_cf_pc; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [38:0] _GEN_498 = _T_11 ? _GEN_246 : REG__2_cf_pc; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [38:0] _GEN_499 = _T_11 ? _GEN_247 : REG__3_cf_pc; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [63:0] _GEN_500 = _T_11 ? _GEN_248 : REG__0_cf_instr; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [63:0] _GEN_501 = _T_11 ? _GEN_249 : REG__1_cf_instr; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [63:0] _GEN_502 = _T_11 ? _GEN_250 : REG__2_cf_instr; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [63:0] _GEN_503 = _T_11 ? _GEN_251 : REG__3_cf_instr; // @[PipelineVector.scala 45:29 PipelineVector.scala 29:29]
  wire [1:0] _T_20 = 2'h1 + REG_1; // @[PipelineVector.scala 46:45]
  wire [63:0] _REG_T_20_data_imm = frontend_io_out_1_bits_data_imm; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire [4:0] _REG_T_20_ctrl_rfDest = frontend_io_out_1_bits_ctrl_rfDest; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire [4:0] _REG_T_20_ctrl_rfSrc2 = frontend_io_out_1_bits_ctrl_rfSrc2; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire [4:0] _REG_T_20_ctrl_rfSrc1 = frontend_io_out_1_bits_ctrl_rfSrc1; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire [6:0] _REG_T_20_ctrl_fuOpType = frontend_io_out_1_bits_ctrl_fuOpType; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire [2:0] _REG_T_20_ctrl_fuType = frontend_io_out_1_bits_ctrl_fuType; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire [3:0] _REG_T_20_cf_brIdx = frontend_io_out_1_bits_cf_brIdx; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire [38:0] _REG_T_20_cf_pnpc = frontend_io_out_1_bits_cf_pnpc; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire [38:0] _REG_T_20_cf_pc = frontend_io_out_1_bits_cf_pc; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire [63:0] _REG_T_20_cf_instr = frontend_io_out_1_bits_cf_instr; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire [1:0] _T_22 = REG_1 + _T_10; // @[PipelineVector.scala 47:42]
  wire [63:0] _GEN_1266 = 2'h1 == REG_2 ? REG__1_data_imm : REG__0_data_imm; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [63:0] _GEN_1267 = 2'h2 == REG_2 ? REG__2_data_imm : _GEN_1266; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [4:0] _GEN_1310 = 2'h1 == REG_2 ? REG__1_ctrl_rfDest : REG__0_ctrl_rfDest; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [4:0] _GEN_1311 = 2'h2 == REG_2 ? REG__2_ctrl_rfDest : _GEN_1310; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1314 = 2'h1 == REG_2 ? REG__1_ctrl_rfWen : REG__0_ctrl_rfWen; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1315 = 2'h2 == REG_2 ? REG__2_ctrl_rfWen : _GEN_1314; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [4:0] _GEN_1318 = 2'h1 == REG_2 ? REG__1_ctrl_rfSrc2 : REG__0_ctrl_rfSrc2; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [4:0] _GEN_1319 = 2'h2 == REG_2 ? REG__2_ctrl_rfSrc2 : _GEN_1318; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [4:0] _GEN_1322 = 2'h1 == REG_2 ? REG__1_ctrl_rfSrc1 : REG__0_ctrl_rfSrc1; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [4:0] _GEN_1323 = 2'h2 == REG_2 ? REG__2_ctrl_rfSrc1 : _GEN_1322; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [6:0] _GEN_1326 = 2'h1 == REG_2 ? REG__1_ctrl_fuOpType : REG__0_ctrl_fuOpType; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [6:0] _GEN_1327 = 2'h2 == REG_2 ? REG__2_ctrl_fuOpType : _GEN_1326; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [2:0] _GEN_1330 = 2'h1 == REG_2 ? REG__1_ctrl_fuType : REG__0_ctrl_fuType; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [2:0] _GEN_1331 = 2'h2 == REG_2 ? REG__2_ctrl_fuType : _GEN_1330; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1334 = 2'h1 == REG_2 ? REG__1_ctrl_src2Type : REG__0_ctrl_src2Type; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1335 = 2'h2 == REG_2 ? REG__2_ctrl_src2Type : _GEN_1334; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1338 = 2'h1 == REG_2 ? REG__1_ctrl_src1Type : REG__0_ctrl_src1Type; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1339 = 2'h2 == REG_2 ? REG__2_ctrl_src1Type : _GEN_1338; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1342 = 2'h1 == REG_2 ? REG__1_cf_crossPageIPFFix : REG__0_cf_crossPageIPFFix; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1343 = 2'h2 == REG_2 ? REG__2_cf_crossPageIPFFix : _GEN_1342; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [3:0] _GEN_1350 = 2'h1 == REG_2 ? REG__1_cf_brIdx : REG__0_cf_brIdx; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [3:0] _GEN_1351 = 2'h2 == REG_2 ? REG__2_cf_brIdx : _GEN_1350; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1354 = 2'h1 == REG_2 ? REG__1_cf_intrVec_0 : REG__0_cf_intrVec_0; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1355 = 2'h2 == REG_2 ? REG__2_cf_intrVec_0 : _GEN_1354; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1358 = 2'h1 == REG_2 ? REG__1_cf_intrVec_1 : REG__0_cf_intrVec_1; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1359 = 2'h2 == REG_2 ? REG__2_cf_intrVec_1 : _GEN_1358; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1362 = 2'h1 == REG_2 ? REG__1_cf_intrVec_2 : REG__0_cf_intrVec_2; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1363 = 2'h2 == REG_2 ? REG__2_cf_intrVec_2 : _GEN_1362; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1366 = 2'h1 == REG_2 ? REG__1_cf_intrVec_3 : REG__0_cf_intrVec_3; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1367 = 2'h2 == REG_2 ? REG__2_cf_intrVec_3 : _GEN_1366; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1370 = 2'h1 == REG_2 ? REG__1_cf_intrVec_4 : REG__0_cf_intrVec_4; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1371 = 2'h2 == REG_2 ? REG__2_cf_intrVec_4 : _GEN_1370; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1374 = 2'h1 == REG_2 ? REG__1_cf_intrVec_5 : REG__0_cf_intrVec_5; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1375 = 2'h2 == REG_2 ? REG__2_cf_intrVec_5 : _GEN_1374; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1378 = 2'h1 == REG_2 ? REG__1_cf_intrVec_6 : REG__0_cf_intrVec_6; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1379 = 2'h2 == REG_2 ? REG__2_cf_intrVec_6 : _GEN_1378; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1382 = 2'h1 == REG_2 ? REG__1_cf_intrVec_7 : REG__0_cf_intrVec_7; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1383 = 2'h2 == REG_2 ? REG__2_cf_intrVec_7 : _GEN_1382; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1386 = 2'h1 == REG_2 ? REG__1_cf_intrVec_8 : REG__0_cf_intrVec_8; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1387 = 2'h2 == REG_2 ? REG__2_cf_intrVec_8 : _GEN_1386; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1390 = 2'h1 == REG_2 ? REG__1_cf_intrVec_9 : REG__0_cf_intrVec_9; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1391 = 2'h2 == REG_2 ? REG__2_cf_intrVec_9 : _GEN_1390; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1394 = 2'h1 == REG_2 ? REG__1_cf_intrVec_10 : REG__0_cf_intrVec_10; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1395 = 2'h2 == REG_2 ? REG__2_cf_intrVec_10 : _GEN_1394; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1398 = 2'h1 == REG_2 ? REG__1_cf_intrVec_11 : REG__0_cf_intrVec_11; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1399 = 2'h2 == REG_2 ? REG__2_cf_intrVec_11 : _GEN_1398; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1406 = 2'h1 == REG_2 ? REG__1_cf_exceptionVec_1 : REG__0_cf_exceptionVec_1; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1407 = 2'h2 == REG_2 ? REG__2_cf_exceptionVec_1 : _GEN_1406; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1410 = 2'h1 == REG_2 ? REG__1_cf_exceptionVec_2 : REG__0_cf_exceptionVec_2; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1411 = 2'h2 == REG_2 ? REG__2_cf_exceptionVec_2 : _GEN_1410; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1450 = 2'h1 == REG_2 ? REG__1_cf_exceptionVec_12 : REG__0_cf_exceptionVec_12; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _GEN_1451 = 2'h2 == REG_2 ? REG__2_cf_exceptionVec_12 : _GEN_1450; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [38:0] _GEN_1502 = 2'h1 == REG_2 ? REG__1_cf_pnpc : REG__0_cf_pnpc; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [38:0] _GEN_1503 = 2'h2 == REG_2 ? REG__2_cf_pnpc : _GEN_1502; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [38:0] _GEN_1506 = 2'h1 == REG_2 ? REG__1_cf_pc : REG__0_cf_pc; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [38:0] _GEN_1507 = 2'h2 == REG_2 ? REG__2_cf_pc : _GEN_1506; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [63:0] _GEN_1510 = 2'h1 == REG_2 ? REG__1_cf_instr : REG__0_cf_instr; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire [63:0] _GEN_1511 = 2'h2 == REG_2 ? REG__2_cf_instr : _GEN_1510; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  wire  _T_32 = Backend_inorder_io_in_0_ready & Backend_inorder_io_in_0_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_34 = {{1'd0}, _T_32}; // @[PipelineVector.scala 64:44]
  wire  _T_35 = _T_34 > 2'h0; // @[PipelineVector.scala 65:35]
  wire [1:0] _T_37 = REG_2 + _T_34; // @[PipelineVector.scala 67:42]
  ysyx_210000_Frontend_inorder frontend ( // @[NutCore.scala 215:34]
    .clock(frontend_clock),
    .reset(frontend_reset),
    .io_out_0_ready(frontend_io_out_0_ready),
    .io_out_0_valid(frontend_io_out_0_valid),
    .io_out_0_bits_cf_instr(frontend_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(frontend_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(frontend_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(frontend_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(frontend_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(frontend_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_0(frontend_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(frontend_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(frontend_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(frontend_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(frontend_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(frontend_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(frontend_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(frontend_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(frontend_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(frontend_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(frontend_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(frontend_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(frontend_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossPageIPFFix(frontend_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_ctrl_src1Type(frontend_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(frontend_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(frontend_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(frontend_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(frontend_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(frontend_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(frontend_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(frontend_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_data_imm(frontend_io_out_0_bits_data_imm),
    .io_out_1_ready(frontend_io_out_1_ready),
    .io_out_1_valid(frontend_io_out_1_valid),
    .io_out_1_bits_cf_instr(frontend_io_out_1_bits_cf_instr),
    .io_out_1_bits_cf_pc(frontend_io_out_1_bits_cf_pc),
    .io_out_1_bits_cf_pnpc(frontend_io_out_1_bits_cf_pnpc),
    .io_out_1_bits_cf_exceptionVec_1(frontend_io_out_1_bits_cf_exceptionVec_1),
    .io_out_1_bits_cf_exceptionVec_2(frontend_io_out_1_bits_cf_exceptionVec_2),
    .io_out_1_bits_cf_exceptionVec_12(frontend_io_out_1_bits_cf_exceptionVec_12),
    .io_out_1_bits_cf_intrVec_0(frontend_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(frontend_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(frontend_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(frontend_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(frontend_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(frontend_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(frontend_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(frontend_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(frontend_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(frontend_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(frontend_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(frontend_io_out_1_bits_cf_intrVec_11),
    .io_out_1_bits_cf_brIdx(frontend_io_out_1_bits_cf_brIdx),
    .io_out_1_bits_cf_crossPageIPFFix(frontend_io_out_1_bits_cf_crossPageIPFFix),
    .io_out_1_bits_ctrl_src1Type(frontend_io_out_1_bits_ctrl_src1Type),
    .io_out_1_bits_ctrl_src2Type(frontend_io_out_1_bits_ctrl_src2Type),
    .io_out_1_bits_ctrl_fuType(frontend_io_out_1_bits_ctrl_fuType),
    .io_out_1_bits_ctrl_fuOpType(frontend_io_out_1_bits_ctrl_fuOpType),
    .io_out_1_bits_ctrl_rfSrc1(frontend_io_out_1_bits_ctrl_rfSrc1),
    .io_out_1_bits_ctrl_rfSrc2(frontend_io_out_1_bits_ctrl_rfSrc2),
    .io_out_1_bits_ctrl_rfWen(frontend_io_out_1_bits_ctrl_rfWen),
    .io_out_1_bits_ctrl_rfDest(frontend_io_out_1_bits_ctrl_rfDest),
    .io_out_1_bits_data_imm(frontend_io_out_1_bits_data_imm),
    .io_imem_req_ready(frontend_io_imem_req_ready),
    .io_imem_req_valid(frontend_io_imem_req_valid),
    .io_imem_req_bits_addr(frontend_io_imem_req_bits_addr),
    .io_imem_req_bits_user(frontend_io_imem_req_bits_user),
    .io_imem_resp_ready(frontend_io_imem_resp_ready),
    .io_imem_resp_valid(frontend_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(frontend_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(frontend_io_imem_resp_bits_user),
    .io_flushVec(frontend_io_flushVec),
    .io_ipf(frontend_io_ipf),
    .io_redirect_target(frontend_io_redirect_target),
    .io_redirect_valid(frontend_io_redirect_valid),
    .flushICache(frontend_flushICache),
    .REG_6_valid(frontend_REG_6_valid),
    .REG_6_pc(frontend_REG_6_pc),
    .REG_6_isMissPredict(frontend_REG_6_isMissPredict),
    .REG_6_actualTarget(frontend_REG_6_actualTarget),
    .REG_6_actualTaken(frontend_REG_6_actualTaken),
    .REG_6_fuOpType(frontend_REG_6_fuOpType),
    .REG_6_btbType(frontend_REG_6_btbType),
    .REG_6_isRVC(frontend_REG_6_isRVC),
    .vmEnable(frontend_vmEnable),
    .intrVec(frontend_intrVec),
    .flushTLB(frontend_flushTLB)
  );
  ysyx_210000_Backend_inorder Backend_inorder ( // @[NutCore.scala 257:25]
    .clock(Backend_inorder_clock),
    .reset(Backend_inorder_reset),
    .io_in_0_ready(Backend_inorder_io_in_0_ready),
    .io_in_0_valid(Backend_inorder_io_in_0_valid),
    .io_in_0_bits_cf_instr(Backend_inorder_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(Backend_inorder_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(Backend_inorder_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(Backend_inorder_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(Backend_inorder_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(Backend_inorder_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_0(Backend_inorder_io_in_0_bits_cf_intrVec_0),
    .io_in_0_bits_cf_intrVec_1(Backend_inorder_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_2(Backend_inorder_io_in_0_bits_cf_intrVec_2),
    .io_in_0_bits_cf_intrVec_3(Backend_inorder_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_4(Backend_inorder_io_in_0_bits_cf_intrVec_4),
    .io_in_0_bits_cf_intrVec_5(Backend_inorder_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_6(Backend_inorder_io_in_0_bits_cf_intrVec_6),
    .io_in_0_bits_cf_intrVec_7(Backend_inorder_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_8(Backend_inorder_io_in_0_bits_cf_intrVec_8),
    .io_in_0_bits_cf_intrVec_9(Backend_inorder_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_10(Backend_inorder_io_in_0_bits_cf_intrVec_10),
    .io_in_0_bits_cf_intrVec_11(Backend_inorder_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(Backend_inorder_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossPageIPFFix(Backend_inorder_io_in_0_bits_cf_crossPageIPFFix),
    .io_in_0_bits_ctrl_src1Type(Backend_inorder_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(Backend_inorder_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(Backend_inorder_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(Backend_inorder_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(Backend_inorder_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(Backend_inorder_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(Backend_inorder_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(Backend_inorder_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_data_imm(Backend_inorder_io_in_0_bits_data_imm),
    .io_flush(Backend_inorder_io_flush),
    .io_dmem_req_ready(Backend_inorder_io_dmem_req_ready),
    .io_dmem_req_valid(Backend_inorder_io_dmem_req_valid),
    .io_dmem_req_bits_addr(Backend_inorder_io_dmem_req_bits_addr),
    .io_dmem_req_bits_size(Backend_inorder_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(Backend_inorder_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_wmask(Backend_inorder_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wdata(Backend_inorder_io_dmem_req_bits_wdata),
    .io_dmem_resp_valid(Backend_inorder_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(Backend_inorder_io_dmem_resp_bits_rdata),
    .io_memMMU_imem_priviledgeMode(Backend_inorder_io_memMMU_imem_priviledgeMode),
    .io_memMMU_dmem_priviledgeMode(Backend_inorder_io_memMMU_dmem_priviledgeMode),
    .io_memMMU_dmem_status_sum(Backend_inorder_io_memMMU_dmem_status_sum),
    .io_memMMU_dmem_status_mxr(Backend_inorder_io_memMMU_dmem_status_mxr),
    .io_memMMU_dmem_loadPF(Backend_inorder_io_memMMU_dmem_loadPF),
    .io_memMMU_dmem_storePF(Backend_inorder_io_memMMU_dmem_storePF),
    .io_memMMU_dmem_addr(Backend_inorder_io_memMMU_dmem_addr),
    .io_redirect_target(Backend_inorder_io_redirect_target),
    .io_redirect_valid(Backend_inorder_io_redirect_valid),
    ._T_28(Backend_inorder__T_28),
    .flushICache(Backend_inorder_flushICache),
    .satp(Backend_inorder_satp),
    .REG_6_valid(Backend_inorder_REG_6_valid),
    .REG_6_pc(Backend_inorder_REG_6_pc),
    .REG_6_isMissPredict(Backend_inorder_REG_6_isMissPredict),
    .REG_6_actualTarget(Backend_inorder_REG_6_actualTarget),
    .REG_6_actualTaken(Backend_inorder_REG_6_actualTaken),
    .REG_6_fuOpType(Backend_inorder_REG_6_fuOpType),
    .REG_6_btbType(Backend_inorder_REG_6_btbType),
    .REG_6_isRVC(Backend_inorder_REG_6_isRVC),
    .io_extra_mtip(Backend_inorder_io_extra_mtip),
    .amoReq(Backend_inorder_amoReq),
    .io_extra_meip_0(Backend_inorder_io_extra_meip_0),
    .vmEnable(Backend_inorder_vmEnable),
    .intrVec(Backend_inorder_intrVec),
    ._T_27(Backend_inorder__T_27),
    .io_extra_msip(Backend_inorder_io_extra_msip),
    .flushTLB(Backend_inorder_flushTLB)
  );
  ysyx_210000_SimpleBusCrossbarNto1 SimpleBusCrossbarNto1 ( // @[NutCore.scala 261:26]
    .clock(SimpleBusCrossbarNto1_clock),
    .reset(SimpleBusCrossbarNto1_reset),
    .io_in_0_req_ready(SimpleBusCrossbarNto1_io_in_0_req_ready),
    .io_in_0_req_valid(SimpleBusCrossbarNto1_io_in_0_req_valid),
    .io_in_0_req_bits_addr(SimpleBusCrossbarNto1_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(SimpleBusCrossbarNto1_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(SimpleBusCrossbarNto1_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(SimpleBusCrossbarNto1_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(SimpleBusCrossbarNto1_io_in_0_req_bits_wdata),
    .io_in_0_resp_ready(SimpleBusCrossbarNto1_io_in_0_resp_ready),
    .io_in_0_resp_valid(SimpleBusCrossbarNto1_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(SimpleBusCrossbarNto1_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(SimpleBusCrossbarNto1_io_in_1_req_ready),
    .io_in_1_req_valid(SimpleBusCrossbarNto1_io_in_1_req_valid),
    .io_in_1_req_bits_addr(SimpleBusCrossbarNto1_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(SimpleBusCrossbarNto1_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(SimpleBusCrossbarNto1_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(SimpleBusCrossbarNto1_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(SimpleBusCrossbarNto1_io_in_1_req_bits_wdata),
    .io_in_1_resp_ready(SimpleBusCrossbarNto1_io_in_1_resp_ready),
    .io_in_1_resp_valid(SimpleBusCrossbarNto1_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(SimpleBusCrossbarNto1_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata),
    .io_out_req_ready(SimpleBusCrossbarNto1_io_out_req_ready),
    .io_out_req_valid(SimpleBusCrossbarNto1_io_out_req_valid),
    .io_out_req_bits_addr(SimpleBusCrossbarNto1_io_out_req_bits_addr),
    .io_out_req_bits_size(SimpleBusCrossbarNto1_io_out_req_bits_size),
    .io_out_req_bits_cmd(SimpleBusCrossbarNto1_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(SimpleBusCrossbarNto1_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(SimpleBusCrossbarNto1_io_out_req_bits_wdata),
    .io_out_resp_ready(SimpleBusCrossbarNto1_io_out_resp_ready),
    .io_out_resp_valid(SimpleBusCrossbarNto1_io_out_resp_valid),
    .io_out_resp_bits_cmd(SimpleBusCrossbarNto1_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(SimpleBusCrossbarNto1_io_out_resp_bits_rdata)
  );
  ysyx_210000_SimpleBusCrossbarNto1_1 SimpleBusCrossbarNto1_1 ( // @[NutCore.scala 262:26]
    .clock(SimpleBusCrossbarNto1_1_clock),
    .reset(SimpleBusCrossbarNto1_1_reset),
    .io_in_0_req_ready(SimpleBusCrossbarNto1_1_io_in_0_req_ready),
    .io_in_0_req_valid(SimpleBusCrossbarNto1_1_io_in_0_req_valid),
    .io_in_0_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(SimpleBusCrossbarNto1_1_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(SimpleBusCrossbarNto1_1_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(SimpleBusCrossbarNto1_1_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(SimpleBusCrossbarNto1_1_io_in_1_req_ready),
    .io_in_1_req_valid(SimpleBusCrossbarNto1_1_io_in_1_req_valid),
    .io_in_1_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_1_req_bits_addr),
    .io_in_1_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(SimpleBusCrossbarNto1_1_io_in_1_resp_valid),
    .io_in_1_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_1_resp_bits_rdata),
    .io_in_2_req_ready(SimpleBusCrossbarNto1_1_io_in_2_req_ready),
    .io_in_2_req_valid(SimpleBusCrossbarNto1_1_io_in_2_req_valid),
    .io_in_2_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_2_req_bits_addr),
    .io_in_2_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_2_req_bits_cmd),
    .io_in_2_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_2_req_bits_wdata),
    .io_in_2_resp_valid(SimpleBusCrossbarNto1_1_io_in_2_resp_valid),
    .io_in_2_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_2_resp_bits_rdata),
    .io_in_3_req_ready(SimpleBusCrossbarNto1_1_io_in_3_req_ready),
    .io_in_3_req_valid(SimpleBusCrossbarNto1_1_io_in_3_req_valid),
    .io_in_3_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_3_req_bits_addr),
    .io_in_3_req_bits_size(SimpleBusCrossbarNto1_1_io_in_3_req_bits_size),
    .io_in_3_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_3_req_bits_cmd),
    .io_in_3_req_bits_wmask(SimpleBusCrossbarNto1_1_io_in_3_req_bits_wmask),
    .io_in_3_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_3_req_bits_wdata),
    .io_in_3_resp_ready(SimpleBusCrossbarNto1_1_io_in_3_resp_ready),
    .io_in_3_resp_valid(SimpleBusCrossbarNto1_1_io_in_3_resp_valid),
    .io_in_3_resp_bits_cmd(SimpleBusCrossbarNto1_1_io_in_3_resp_bits_cmd),
    .io_in_3_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_3_resp_bits_rdata),
    .io_out_req_ready(SimpleBusCrossbarNto1_1_io_out_req_ready),
    .io_out_req_valid(SimpleBusCrossbarNto1_1_io_out_req_valid),
    .io_out_req_bits_addr(SimpleBusCrossbarNto1_1_io_out_req_bits_addr),
    .io_out_req_bits_size(SimpleBusCrossbarNto1_1_io_out_req_bits_size),
    .io_out_req_bits_cmd(SimpleBusCrossbarNto1_1_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(SimpleBusCrossbarNto1_1_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(SimpleBusCrossbarNto1_1_io_out_req_bits_wdata),
    .io_out_resp_ready(SimpleBusCrossbarNto1_1_io_out_resp_ready),
    .io_out_resp_valid(SimpleBusCrossbarNto1_1_io_out_resp_valid),
    .io_out_resp_bits_cmd(SimpleBusCrossbarNto1_1_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_out_resp_bits_rdata)
  );
  ysyx_210000_MMIOBridge MMIOBridge ( // @[NutCore.scala 264:28]
    .clock(MMIOBridge_clock),
    .reset(MMIOBridge_reset),
    .io_in_req_ready(MMIOBridge_io_in_req_ready),
    .io_in_req_valid(MMIOBridge_io_in_req_valid),
    .io_in_req_bits_addr(MMIOBridge_io_in_req_bits_addr),
    .io_in_req_bits_size(MMIOBridge_io_in_req_bits_size),
    .io_in_resp_valid(MMIOBridge_io_in_resp_valid),
    .io_in_resp_bits_rdata(MMIOBridge_io_in_resp_bits_rdata),
    .io_out_req_ready(MMIOBridge_io_out_req_ready),
    .io_out_req_valid(MMIOBridge_io_out_req_valid),
    .io_out_req_bits_addr(MMIOBridge_io_out_req_bits_addr),
    .io_out_req_bits_size(MMIOBridge_io_out_req_bits_size),
    .io_out_resp_ready(MMIOBridge_io_out_resp_ready),
    .io_out_resp_valid(MMIOBridge_io_out_resp_valid),
    .io_out_resp_bits_rdata(MMIOBridge_io_out_resp_bits_rdata)
  );
  ysyx_210000_EmbeddedTLB EmbeddedTLB ( // @[EmbeddedTLB.scala 427:23]
    .clock(EmbeddedTLB_clock),
    .reset(EmbeddedTLB_reset),
    .io_in_req_ready(EmbeddedTLB_io_in_req_ready),
    .io_in_req_valid(EmbeddedTLB_io_in_req_valid),
    .io_in_req_bits_addr(EmbeddedTLB_io_in_req_bits_addr),
    .io_in_req_bits_user(EmbeddedTLB_io_in_req_bits_user),
    .io_in_resp_ready(EmbeddedTLB_io_in_resp_ready),
    .io_in_resp_valid(EmbeddedTLB_io_in_resp_valid),
    .io_in_resp_bits_rdata(EmbeddedTLB_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(EmbeddedTLB_io_in_resp_bits_user),
    .io_out_req_ready(EmbeddedTLB_io_out_req_ready),
    .io_out_req_valid(EmbeddedTLB_io_out_req_valid),
    .io_out_req_bits_addr(EmbeddedTLB_io_out_req_bits_addr),
    .io_out_req_bits_size(EmbeddedTLB_io_out_req_bits_size),
    .io_out_req_bits_user(EmbeddedTLB_io_out_req_bits_user),
    .io_out_resp_ready(EmbeddedTLB_io_out_resp_ready),
    .io_out_resp_valid(EmbeddedTLB_io_out_resp_valid),
    .io_out_resp_bits_rdata(EmbeddedTLB_io_out_resp_bits_rdata),
    .io_out_resp_bits_user(EmbeddedTLB_io_out_resp_bits_user),
    .io_mem_req_ready(EmbeddedTLB_io_mem_req_ready),
    .io_mem_req_valid(EmbeddedTLB_io_mem_req_valid),
    .io_mem_req_bits_addr(EmbeddedTLB_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(EmbeddedTLB_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(EmbeddedTLB_io_mem_req_bits_wdata),
    .io_mem_resp_valid(EmbeddedTLB_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(EmbeddedTLB_io_mem_resp_bits_rdata),
    .io_flush(EmbeddedTLB_io_flush),
    .io_csrMMU_priviledgeMode(EmbeddedTLB_io_csrMMU_priviledgeMode),
    .io_cacheEmpty(EmbeddedTLB_io_cacheEmpty),
    .io_ipf(EmbeddedTLB_io_ipf),
    .CSRSATP(EmbeddedTLB_CSRSATP),
    .MOUFlushTLB(EmbeddedTLB_MOUFlushTLB)
  );
  ysyx_210000_Cache Cache ( // @[Cache.scala 679:35]
    .clock(Cache_clock),
    .reset(Cache_reset),
    .io_in_req_ready(Cache_io_in_req_ready),
    .io_in_req_valid(Cache_io_in_req_valid),
    .io_in_req_bits_addr(Cache_io_in_req_bits_addr),
    .io_in_req_bits_size(Cache_io_in_req_bits_size),
    .io_in_req_bits_user(Cache_io_in_req_bits_user),
    .io_in_resp_ready(Cache_io_in_resp_ready),
    .io_in_resp_valid(Cache_io_in_resp_valid),
    .io_in_resp_bits_rdata(Cache_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(Cache_io_in_resp_bits_user),
    .io_flush(Cache_io_flush),
    .io_out_mem_req_ready(Cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(Cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(Cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(Cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(Cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(Cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(Cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(Cache_io_out_mem_resp_bits_rdata),
    .io_mmio_req_ready(Cache_io_mmio_req_ready),
    .io_mmio_req_valid(Cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(Cache_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(Cache_io_mmio_req_bits_size),
    .io_mmio_resp_valid(Cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(Cache_io_mmio_resp_bits_rdata),
    .io_empty(Cache_io_empty),
    .MOUFlushICache(Cache_MOUFlushICache)
  );
  ysyx_210000_EmbeddedTLB_1 EmbeddedTLB_1 ( // @[EmbeddedTLB.scala 427:23]
    .clock(EmbeddedTLB_1_clock),
    .reset(EmbeddedTLB_1_reset),
    .io_in_req_ready(EmbeddedTLB_1_io_in_req_ready),
    .io_in_req_valid(EmbeddedTLB_1_io_in_req_valid),
    .io_in_req_bits_addr(EmbeddedTLB_1_io_in_req_bits_addr),
    .io_in_req_bits_size(EmbeddedTLB_1_io_in_req_bits_size),
    .io_in_req_bits_cmd(EmbeddedTLB_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(EmbeddedTLB_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(EmbeddedTLB_1_io_in_req_bits_wdata),
    .io_in_resp_valid(EmbeddedTLB_1_io_in_resp_valid),
    .io_in_resp_bits_rdata(EmbeddedTLB_1_io_in_resp_bits_rdata),
    .io_out_req_ready(EmbeddedTLB_1_io_out_req_ready),
    .io_out_req_valid(EmbeddedTLB_1_io_out_req_valid),
    .io_out_req_bits_addr(EmbeddedTLB_1_io_out_req_bits_addr),
    .io_out_req_bits_size(EmbeddedTLB_1_io_out_req_bits_size),
    .io_out_req_bits_cmd(EmbeddedTLB_1_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(EmbeddedTLB_1_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(EmbeddedTLB_1_io_out_req_bits_wdata),
    .io_out_resp_valid(EmbeddedTLB_1_io_out_resp_valid),
    .io_out_resp_bits_rdata(EmbeddedTLB_1_io_out_resp_bits_rdata),
    .io_mem_req_ready(EmbeddedTLB_1_io_mem_req_ready),
    .io_mem_req_valid(EmbeddedTLB_1_io_mem_req_valid),
    .io_mem_req_bits_addr(EmbeddedTLB_1_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(EmbeddedTLB_1_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(EmbeddedTLB_1_io_mem_req_bits_wdata),
    .io_mem_resp_valid(EmbeddedTLB_1_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(EmbeddedTLB_1_io_mem_resp_bits_rdata),
    .io_csrMMU_priviledgeMode(EmbeddedTLB_1_io_csrMMU_priviledgeMode),
    .io_csrMMU_status_sum(EmbeddedTLB_1_io_csrMMU_status_sum),
    .io_csrMMU_status_mxr(EmbeddedTLB_1_io_csrMMU_status_mxr),
    .io_csrMMU_loadPF(EmbeddedTLB_1_io_csrMMU_loadPF),
    .io_csrMMU_storePF(EmbeddedTLB_1_io_csrMMU_storePF),
    .io_csrMMU_addr(EmbeddedTLB_1_io_csrMMU_addr),
    ._T_28_0(EmbeddedTLB_1__T_28_0),
    .CSRSATP(EmbeddedTLB_1_CSRSATP),
    .amoReq(EmbeddedTLB_1_amoReq),
    .vmEnable_0(EmbeddedTLB_1_vmEnable_0),
    ._T_27_0(EmbeddedTLB_1__T_27_0),
    .MOUFlushTLB(EmbeddedTLB_1_MOUFlushTLB)
  );
  ysyx_210000_Cache_1 Cache_1 ( // @[Cache.scala 679:35]
    .clock(Cache_1_clock),
    .reset(Cache_1_reset),
    .io_in_req_ready(Cache_1_io_in_req_ready),
    .io_in_req_valid(Cache_1_io_in_req_valid),
    .io_in_req_bits_addr(Cache_1_io_in_req_bits_addr),
    .io_in_req_bits_size(Cache_1_io_in_req_bits_size),
    .io_in_req_bits_cmd(Cache_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(Cache_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(Cache_1_io_in_req_bits_wdata),
    .io_in_resp_ready(Cache_1_io_in_resp_ready),
    .io_in_resp_valid(Cache_1_io_in_resp_valid),
    .io_in_resp_bits_cmd(Cache_1_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(Cache_1_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(Cache_1_io_out_mem_req_ready),
    .io_out_mem_req_valid(Cache_1_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(Cache_1_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(Cache_1_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(Cache_1_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(Cache_1_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(Cache_1_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(Cache_1_io_out_mem_resp_bits_rdata),
    .io_out_coh_req_ready(Cache_1_io_out_coh_req_ready),
    .io_out_coh_req_valid(Cache_1_io_out_coh_req_valid),
    .io_out_coh_req_bits_addr(Cache_1_io_out_coh_req_bits_addr),
    .io_out_coh_req_bits_wdata(Cache_1_io_out_coh_req_bits_wdata),
    .io_out_coh_resp_valid(Cache_1_io_out_coh_resp_valid),
    .io_out_coh_resp_bits_cmd(Cache_1_io_out_coh_resp_bits_cmd),
    .io_out_coh_resp_bits_rdata(Cache_1_io_out_coh_resp_bits_rdata),
    .io_mmio_req_ready(Cache_1_io_mmio_req_ready),
    .io_mmio_req_valid(Cache_1_io_mmio_req_valid),
    .io_mmio_req_bits_addr(Cache_1_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(Cache_1_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(Cache_1_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(Cache_1_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(Cache_1_io_mmio_req_bits_wdata),
    .io_mmio_resp_valid(Cache_1_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(Cache_1_io_mmio_resp_bits_rdata)
  );
  assign io_imem_mem_req_valid = Cache_io_out_mem_req_valid; // @[NutCore.scala 269:13]
  assign io_imem_mem_req_bits_addr = Cache_io_out_mem_req_bits_addr; // @[NutCore.scala 269:13]
  assign io_imem_mem_req_bits_cmd = Cache_io_out_mem_req_bits_cmd; // @[NutCore.scala 269:13]
  assign io_imem_mem_req_bits_wdata = Cache_io_out_mem_req_bits_wdata; // @[NutCore.scala 269:13]
  assign io_dmem_mem_req_valid = Cache_1_io_out_mem_req_valid; // @[NutCore.scala 277:13]
  assign io_dmem_mem_req_bits_addr = Cache_1_io_out_mem_req_bits_addr; // @[NutCore.scala 277:13]
  assign io_dmem_mem_req_bits_cmd = Cache_1_io_out_mem_req_bits_cmd; // @[NutCore.scala 277:13]
  assign io_dmem_mem_req_bits_wdata = Cache_1_io_out_mem_req_bits_wdata; // @[NutCore.scala 277:13]
  assign io_dmem_coh_req_ready = Cache_1_io_out_coh_req_ready; // @[NutCore.scala 277:13]
  assign io_dmem_coh_resp_valid = Cache_1_io_out_coh_resp_valid; // @[NutCore.scala 277:13]
  assign io_dmem_coh_resp_bits_cmd = Cache_1_io_out_coh_resp_bits_cmd; // @[NutCore.scala 277:13]
  assign io_dmem_coh_resp_bits_rdata = Cache_1_io_out_coh_resp_bits_rdata; // @[NutCore.scala 277:13]
  assign io_mmio_req_valid = SimpleBusCrossbarNto1_io_out_req_valid; // @[NutCore.scala 286:13]
  assign io_mmio_req_bits_addr = SimpleBusCrossbarNto1_io_out_req_bits_addr; // @[NutCore.scala 286:13]
  assign io_mmio_req_bits_size = SimpleBusCrossbarNto1_io_out_req_bits_size; // @[NutCore.scala 286:13]
  assign io_mmio_req_bits_cmd = SimpleBusCrossbarNto1_io_out_req_bits_cmd; // @[NutCore.scala 286:13]
  assign io_mmio_req_bits_wmask = SimpleBusCrossbarNto1_io_out_req_bits_wmask; // @[NutCore.scala 286:13]
  assign io_mmio_req_bits_wdata = SimpleBusCrossbarNto1_io_out_req_bits_wdata; // @[NutCore.scala 286:13]
  assign io_mmio_resp_ready = SimpleBusCrossbarNto1_io_out_resp_ready; // @[NutCore.scala 286:13]
  assign io_frontend_req_ready = SimpleBusCrossbarNto1_1_io_in_3_req_ready; // @[NutCore.scala 284:23]
  assign io_frontend_resp_valid = SimpleBusCrossbarNto1_1_io_in_3_resp_valid; // @[NutCore.scala 284:23]
  assign io_frontend_resp_bits_cmd = SimpleBusCrossbarNto1_1_io_in_3_resp_bits_cmd; // @[NutCore.scala 284:23]
  assign io_frontend_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_3_resp_bits_rdata; // @[NutCore.scala 284:23]
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_io_out_0_ready = _T_9 | ~frontend_io_out_0_valid; // @[PipelineVector.scala 50:36]
  assign frontend_io_out_1_ready = _T_9 | ~frontend_io_out_1_valid; // @[PipelineVector.scala 51:36]
  assign frontend_io_imem_req_ready = EmbeddedTLB_io_in_req_ready; // @[EmbeddedTLB.scala 428:17]
  assign frontend_io_imem_resp_valid = EmbeddedTLB_io_in_resp_valid; // @[EmbeddedTLB.scala 428:17]
  assign frontend_io_imem_resp_bits_rdata = EmbeddedTLB_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 428:17]
  assign frontend_io_imem_resp_bits_user = EmbeddedTLB_io_in_resp_bits_user; // @[EmbeddedTLB.scala 428:17]
  assign frontend_io_ipf = EmbeddedTLB_io_ipf; // @[NutCore.scala 268:21]
  assign frontend_io_redirect_target = Backend_inorder_io_redirect_target; // @[NutCore.scala 280:26]
  assign frontend_io_redirect_valid = Backend_inorder_io_redirect_valid; // @[NutCore.scala 280:26]
  assign frontend_flushICache = Backend_inorder_flushICache;
  assign frontend_REG_6_valid = Backend_inorder_REG_6_valid;
  assign frontend_REG_6_pc = Backend_inorder_REG_6_pc;
  assign frontend_REG_6_isMissPredict = Backend_inorder_REG_6_isMissPredict;
  assign frontend_REG_6_actualTarget = Backend_inorder_REG_6_actualTarget;
  assign frontend_REG_6_actualTaken = Backend_inorder_REG_6_actualTaken;
  assign frontend_REG_6_fuOpType = Backend_inorder_REG_6_fuOpType;
  assign frontend_REG_6_btbType = Backend_inorder_REG_6_btbType;
  assign frontend_REG_6_isRVC = Backend_inorder_REG_6_isRVC;
  assign frontend_vmEnable = EmbeddedTLB_1_vmEnable_0;
  assign frontend_intrVec = Backend_inorder_intrVec;
  assign frontend_flushTLB = Backend_inorder_flushTLB;
  assign Backend_inorder_clock = clock;
  assign Backend_inorder_reset = reset;
  assign Backend_inorder_io_in_0_valid = REG_1 != REG_2; // @[PipelineVector.scala 56:34]
  assign Backend_inorder_io_in_0_bits_cf_instr = 2'h3 == REG_2 ? REG__3_cf_instr : _GEN_1511; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_pc = 2'h3 == REG_2 ? REG__3_cf_pc : _GEN_1507; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_pnpc = 2'h3 == REG_2 ? REG__3_cf_pnpc : _GEN_1503; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_exceptionVec_1 = 2'h3 == REG_2 ? REG__3_cf_exceptionVec_1 : _GEN_1407; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_exceptionVec_2 = 2'h3 == REG_2 ? REG__3_cf_exceptionVec_2 : _GEN_1411; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_exceptionVec_12 = 2'h3 == REG_2 ? REG__3_cf_exceptionVec_12 : _GEN_1451; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_0 = 2'h3 == REG_2 ? REG__3_cf_intrVec_0 : _GEN_1355; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_1 = 2'h3 == REG_2 ? REG__3_cf_intrVec_1 : _GEN_1359; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_2 = 2'h3 == REG_2 ? REG__3_cf_intrVec_2 : _GEN_1363; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_3 = 2'h3 == REG_2 ? REG__3_cf_intrVec_3 : _GEN_1367; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_4 = 2'h3 == REG_2 ? REG__3_cf_intrVec_4 : _GEN_1371; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_5 = 2'h3 == REG_2 ? REG__3_cf_intrVec_5 : _GEN_1375; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_6 = 2'h3 == REG_2 ? REG__3_cf_intrVec_6 : _GEN_1379; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_7 = 2'h3 == REG_2 ? REG__3_cf_intrVec_7 : _GEN_1383; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_8 = 2'h3 == REG_2 ? REG__3_cf_intrVec_8 : _GEN_1387; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_9 = 2'h3 == REG_2 ? REG__3_cf_intrVec_9 : _GEN_1391; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_10 = 2'h3 == REG_2 ? REG__3_cf_intrVec_10 : _GEN_1395; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_11 = 2'h3 == REG_2 ? REG__3_cf_intrVec_11 : _GEN_1399; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_brIdx = 2'h3 == REG_2 ? REG__3_cf_brIdx : _GEN_1351; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_crossPageIPFFix = 2'h3 == REG_2 ? REG__3_cf_crossPageIPFFix : _GEN_1343; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_src1Type = 2'h3 == REG_2 ? REG__3_ctrl_src1Type : _GEN_1339; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_src2Type = 2'h3 == REG_2 ? REG__3_ctrl_src2Type : _GEN_1335; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_fuType = 2'h3 == REG_2 ? REG__3_ctrl_fuType : _GEN_1331; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_fuOpType = 2'h3 == REG_2 ? REG__3_ctrl_fuOpType : _GEN_1327; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_rfSrc1 = 2'h3 == REG_2 ? REG__3_ctrl_rfSrc1 : _GEN_1323; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_rfSrc2 = 2'h3 == REG_2 ? REG__3_ctrl_rfSrc2 : _GEN_1319; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_rfWen = 2'h3 == REG_2 ? REG__3_ctrl_rfWen : _GEN_1315; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_rfDest = 2'h3 == REG_2 ? REG__3_ctrl_rfDest : _GEN_1311; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_data_imm = 2'h3 == REG_2 ? REG__3_data_imm : _GEN_1267; // @[PipelineVector.scala 55:15 PipelineVector.scala 55:15]
  assign Backend_inorder_io_flush = frontend_io_flushVec[3:2]; // @[NutCore.scala 281:45]
  assign Backend_inorder_io_dmem_req_ready = EmbeddedTLB_1_io_in_req_ready; // @[EmbeddedTLB.scala 428:17]
  assign Backend_inorder_io_dmem_resp_valid = EmbeddedTLB_1_io_in_resp_valid; // @[EmbeddedTLB.scala 428:17]
  assign Backend_inorder_io_dmem_resp_bits_rdata = EmbeddedTLB_1_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 428:17]
  assign Backend_inorder_io_memMMU_dmem_loadPF = EmbeddedTLB_1_io_csrMMU_loadPF; // @[EmbeddedTLB.scala 431:21]
  assign Backend_inorder_io_memMMU_dmem_storePF = EmbeddedTLB_1_io_csrMMU_storePF; // @[EmbeddedTLB.scala 431:21]
  assign Backend_inorder_io_memMMU_dmem_addr = EmbeddedTLB_1_io_csrMMU_addr; // @[EmbeddedTLB.scala 431:21]
  assign Backend_inorder__T_28 = EmbeddedTLB_1__T_28_0;
  assign Backend_inorder_io_extra_mtip = io_extra_mtip;
  assign Backend_inorder_io_extra_meip_0 = io_extra_meip_0;
  assign Backend_inorder_vmEnable = EmbeddedTLB_1_vmEnable_0;
  assign Backend_inorder__T_27 = EmbeddedTLB_1__T_27_0;
  assign Backend_inorder_io_extra_msip = io_extra_msip;
  assign SimpleBusCrossbarNto1_clock = clock;
  assign SimpleBusCrossbarNto1_reset = reset;
  assign SimpleBusCrossbarNto1_io_in_0_req_valid = MMIOBridge_io_out_req_valid; // @[NutCore.scala 272:23]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_addr = MMIOBridge_io_out_req_bits_addr; // @[NutCore.scala 272:23]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_size = MMIOBridge_io_out_req_bits_size; // @[NutCore.scala 272:23]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_cmd = 4'h0; // @[NutCore.scala 272:23]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_wmask = 8'h0; // @[NutCore.scala 272:23]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_wdata = 64'h0; // @[NutCore.scala 272:23]
  assign SimpleBusCrossbarNto1_io_in_0_resp_ready = 1'h1; // @[NutCore.scala 272:23]
  assign SimpleBusCrossbarNto1_io_in_1_req_valid = Cache_1_io_mmio_req_valid; // @[Cache.scala 686:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_addr = Cache_1_io_mmio_req_bits_addr; // @[Cache.scala 686:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_size = Cache_1_io_mmio_req_bits_size; // @[Cache.scala 686:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_cmd = Cache_1_io_mmio_req_bits_cmd; // @[Cache.scala 686:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_wmask = Cache_1_io_mmio_req_bits_wmask; // @[Cache.scala 686:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_wdata = Cache_1_io_mmio_req_bits_wdata; // @[Cache.scala 686:13]
  assign SimpleBusCrossbarNto1_io_in_1_resp_ready = 1'h1; // @[Cache.scala 686:13]
  assign SimpleBusCrossbarNto1_io_out_req_ready = io_mmio_req_ready; // @[NutCore.scala 286:13]
  assign SimpleBusCrossbarNto1_io_out_resp_valid = io_mmio_resp_valid; // @[NutCore.scala 286:13]
  assign SimpleBusCrossbarNto1_io_out_resp_bits_cmd = io_mmio_resp_bits_cmd; // @[NutCore.scala 286:13]
  assign SimpleBusCrossbarNto1_io_out_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[NutCore.scala 286:13]
  assign SimpleBusCrossbarNto1_1_clock = clock;
  assign SimpleBusCrossbarNto1_1_reset = reset;
  assign SimpleBusCrossbarNto1_1_io_in_0_req_valid = EmbeddedTLB_1_io_out_req_valid; // @[NutCore.scala 276:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_addr = EmbeddedTLB_1_io_out_req_bits_addr; // @[NutCore.scala 276:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_size = EmbeddedTLB_1_io_out_req_bits_size; // @[NutCore.scala 276:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_cmd = EmbeddedTLB_1_io_out_req_bits_cmd; // @[NutCore.scala 276:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_wmask = EmbeddedTLB_1_io_out_req_bits_wmask; // @[NutCore.scala 276:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_wdata = EmbeddedTLB_1_io_out_req_bits_wdata; // @[NutCore.scala 276:23]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_valid = EmbeddedTLB_io_mem_req_valid; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_bits_addr = EmbeddedTLB_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_bits_cmd = EmbeddedTLB_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_bits_wdata = EmbeddedTLB_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_valid = EmbeddedTLB_1_io_mem_req_valid; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_bits_addr = EmbeddedTLB_1_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_bits_cmd = EmbeddedTLB_1_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_bits_wdata = EmbeddedTLB_1_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_valid = io_frontend_req_valid; // @[NutCore.scala 284:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_addr = io_frontend_req_bits_addr; // @[NutCore.scala 284:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_size = io_frontend_req_bits_size; // @[NutCore.scala 284:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_cmd = io_frontend_req_bits_cmd; // @[NutCore.scala 284:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_wmask = io_frontend_req_bits_wmask; // @[NutCore.scala 284:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_wdata = io_frontend_req_bits_wdata; // @[NutCore.scala 284:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_resp_ready = io_frontend_resp_ready; // @[NutCore.scala 284:23]
  assign SimpleBusCrossbarNto1_1_io_out_req_ready = Cache_1_io_in_req_ready; // @[Cache.scala 685:17]
  assign SimpleBusCrossbarNto1_1_io_out_resp_valid = Cache_1_io_in_resp_valid; // @[Cache.scala 685:17]
  assign SimpleBusCrossbarNto1_1_io_out_resp_bits_cmd = Cache_1_io_in_resp_bits_cmd; // @[Cache.scala 685:17]
  assign SimpleBusCrossbarNto1_1_io_out_resp_bits_rdata = Cache_1_io_in_resp_bits_rdata; // @[Cache.scala 685:17]
  assign MMIOBridge_clock = clock;
  assign MMIOBridge_reset = reset;
  assign MMIOBridge_io_in_req_valid = Cache_io_mmio_req_valid; // @[NutCore.scala 271:14]
  assign MMIOBridge_io_in_req_bits_addr = Cache_io_mmio_req_bits_addr; // @[NutCore.scala 271:14]
  assign MMIOBridge_io_in_req_bits_size = Cache_io_mmio_req_bits_size; // @[NutCore.scala 271:14]
  assign MMIOBridge_io_out_req_ready = SimpleBusCrossbarNto1_io_in_0_req_ready; // @[NutCore.scala 272:23]
  assign MMIOBridge_io_out_resp_valid = SimpleBusCrossbarNto1_io_in_0_resp_valid; // @[NutCore.scala 272:23]
  assign MMIOBridge_io_out_resp_bits_rdata = SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata; // @[NutCore.scala 272:23]
  assign EmbeddedTLB_clock = clock;
  assign EmbeddedTLB_reset = reset;
  assign EmbeddedTLB_io_in_req_valid = frontend_io_imem_req_valid; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_io_in_req_bits_addr = frontend_io_imem_req_bits_addr; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_io_in_req_bits_user = frontend_io_imem_req_bits_user; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_io_in_resp_ready = frontend_io_imem_resp_ready; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_io_out_req_ready = Cache_io_in_req_ready; // @[Cache.scala 685:17]
  assign EmbeddedTLB_io_out_resp_valid = Cache_io_in_resp_valid; // @[Cache.scala 685:17]
  assign EmbeddedTLB_io_out_resp_bits_rdata = Cache_io_in_resp_bits_rdata; // @[Cache.scala 685:17]
  assign EmbeddedTLB_io_out_resp_bits_user = Cache_io_in_resp_bits_user; // @[Cache.scala 685:17]
  assign EmbeddedTLB_io_mem_req_ready = SimpleBusCrossbarNto1_1_io_in_1_req_ready; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_io_mem_resp_valid = SimpleBusCrossbarNto1_1_io_in_1_resp_valid; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_io_mem_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_1_resp_bits_rdata; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_io_flush = frontend_io_flushVec[0]; // @[NutCore.scala 267:104]
  assign EmbeddedTLB_io_csrMMU_priviledgeMode = Backend_inorder_io_memMMU_imem_priviledgeMode; // @[EmbeddedTLB.scala 431:21]
  assign EmbeddedTLB_io_cacheEmpty = Cache_io_empty; // @[Cache.scala 687:11]
  assign EmbeddedTLB_CSRSATP = Backend_inorder_satp;
  assign EmbeddedTLB_MOUFlushTLB = Backend_inorder_flushTLB;
  assign Cache_clock = clock;
  assign Cache_reset = reset;
  assign Cache_io_in_req_valid = EmbeddedTLB_io_out_req_valid; // @[Cache.scala 685:17]
  assign Cache_io_in_req_bits_addr = EmbeddedTLB_io_out_req_bits_addr; // @[Cache.scala 685:17]
  assign Cache_io_in_req_bits_size = EmbeddedTLB_io_out_req_bits_size; // @[Cache.scala 685:17]
  assign Cache_io_in_req_bits_user = EmbeddedTLB_io_out_req_bits_user; // @[Cache.scala 685:17]
  assign Cache_io_in_resp_ready = EmbeddedTLB_io_out_resp_ready; // @[Cache.scala 685:17]
  assign Cache_io_flush = frontend_io_flushVec[0] ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  assign Cache_io_out_mem_req_ready = io_imem_mem_req_ready; // @[NutCore.scala 269:13]
  assign Cache_io_out_mem_resp_valid = io_imem_mem_resp_valid; // @[NutCore.scala 269:13]
  assign Cache_io_out_mem_resp_bits_cmd = io_imem_mem_resp_bits_cmd; // @[NutCore.scala 269:13]
  assign Cache_io_out_mem_resp_bits_rdata = io_imem_mem_resp_bits_rdata; // @[NutCore.scala 269:13]
  assign Cache_io_mmio_req_ready = MMIOBridge_io_in_req_ready; // @[Cache.scala 686:13]
  assign Cache_io_mmio_resp_valid = MMIOBridge_io_in_resp_valid; // @[Cache.scala 686:13]
  assign Cache_io_mmio_resp_bits_rdata = MMIOBridge_io_in_resp_bits_rdata; // @[Cache.scala 686:13]
  assign Cache_MOUFlushICache = Backend_inorder_flushICache;
  assign EmbeddedTLB_1_clock = clock;
  assign EmbeddedTLB_1_reset = reset;
  assign EmbeddedTLB_1_io_in_req_valid = Backend_inorder_io_dmem_req_valid; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_addr = Backend_inorder_io_dmem_req_bits_addr; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_size = Backend_inorder_io_dmem_req_bits_size; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_cmd = Backend_inorder_io_dmem_req_bits_cmd; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_wmask = Backend_inorder_io_dmem_req_bits_wmask; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_wdata = Backend_inorder_io_dmem_req_bits_wdata; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_out_req_ready = SimpleBusCrossbarNto1_1_io_in_0_req_ready; // @[NutCore.scala 276:23]
  assign EmbeddedTLB_1_io_out_resp_valid = SimpleBusCrossbarNto1_1_io_in_0_resp_valid; // @[NutCore.scala 276:23]
  assign EmbeddedTLB_1_io_out_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_0_resp_bits_rdata; // @[NutCore.scala 276:23]
  assign EmbeddedTLB_1_io_mem_req_ready = SimpleBusCrossbarNto1_1_io_in_2_req_ready; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_1_io_mem_resp_valid = SimpleBusCrossbarNto1_1_io_in_2_resp_valid; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_1_io_mem_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_2_resp_bits_rdata; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_1_io_csrMMU_priviledgeMode = Backend_inorder_io_memMMU_dmem_priviledgeMode; // @[EmbeddedTLB.scala 431:21]
  assign EmbeddedTLB_1_io_csrMMU_status_sum = Backend_inorder_io_memMMU_dmem_status_sum; // @[EmbeddedTLB.scala 431:21]
  assign EmbeddedTLB_1_io_csrMMU_status_mxr = Backend_inorder_io_memMMU_dmem_status_mxr; // @[EmbeddedTLB.scala 431:21]
  assign EmbeddedTLB_1_CSRSATP = Backend_inorder_satp;
  assign EmbeddedTLB_1_amoReq = Backend_inorder_amoReq;
  assign EmbeddedTLB_1_MOUFlushTLB = Backend_inorder_flushTLB;
  assign Cache_1_clock = clock;
  assign Cache_1_reset = reset;
  assign Cache_1_io_in_req_valid = SimpleBusCrossbarNto1_1_io_out_req_valid; // @[Cache.scala 685:17]
  assign Cache_1_io_in_req_bits_addr = SimpleBusCrossbarNto1_1_io_out_req_bits_addr; // @[Cache.scala 685:17]
  assign Cache_1_io_in_req_bits_size = SimpleBusCrossbarNto1_1_io_out_req_bits_size; // @[Cache.scala 685:17]
  assign Cache_1_io_in_req_bits_cmd = SimpleBusCrossbarNto1_1_io_out_req_bits_cmd; // @[Cache.scala 685:17]
  assign Cache_1_io_in_req_bits_wmask = SimpleBusCrossbarNto1_1_io_out_req_bits_wmask; // @[Cache.scala 685:17]
  assign Cache_1_io_in_req_bits_wdata = SimpleBusCrossbarNto1_1_io_out_req_bits_wdata; // @[Cache.scala 685:17]
  assign Cache_1_io_in_resp_ready = SimpleBusCrossbarNto1_1_io_out_resp_ready; // @[Cache.scala 685:17]
  assign Cache_1_io_out_mem_req_ready = io_dmem_mem_req_ready; // @[NutCore.scala 277:13]
  assign Cache_1_io_out_mem_resp_valid = io_dmem_mem_resp_valid; // @[NutCore.scala 277:13]
  assign Cache_1_io_out_mem_resp_bits_cmd = io_dmem_mem_resp_bits_cmd; // @[NutCore.scala 277:13]
  assign Cache_1_io_out_mem_resp_bits_rdata = io_dmem_mem_resp_bits_rdata; // @[NutCore.scala 277:13]
  assign Cache_1_io_out_coh_req_valid = io_dmem_coh_req_valid; // @[NutCore.scala 277:13]
  assign Cache_1_io_out_coh_req_bits_addr = io_dmem_coh_req_bits_addr; // @[NutCore.scala 277:13]
  assign Cache_1_io_out_coh_req_bits_wdata = io_dmem_coh_req_bits_wdata; // @[NutCore.scala 277:13]
  assign Cache_1_io_mmio_req_ready = SimpleBusCrossbarNto1_io_in_1_req_ready; // @[Cache.scala 686:13]
  assign Cache_1_io_mmio_resp_valid = SimpleBusCrossbarNto1_io_in_1_resp_valid; // @[Cache.scala 686:13]
  assign Cache_1_io_mmio_resp_bits_rdata = SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata; // @[Cache.scala 686:13]
  always @(posedge clock) begin
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_instr <= _REG_T_20_cf_instr; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_instr <= _GEN_500;
        end
      end else begin
        REG__0_cf_instr <= _GEN_500;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_pc <= _REG_T_20_cf_pc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_pc <= _GEN_496;
        end
      end else begin
        REG__0_cf_pc <= _GEN_496;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_pnpc <= _REG_T_20_cf_pnpc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_pnpc <= _GEN_492;
        end
      end else begin
        REG__0_cf_pnpc <= _GEN_492;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_exceptionVec_1 <= frontend_io_out_1_bits_cf_exceptionVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_exceptionVec_1 <= _GEN_396;
        end
      end else begin
        REG__0_cf_exceptionVec_1 <= _GEN_396;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_exceptionVec_2 <= frontend_io_out_1_bits_cf_exceptionVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_exceptionVec_2 <= _GEN_400;
        end
      end else begin
        REG__0_cf_exceptionVec_2 <= _GEN_400;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_exceptionVec_12 <= frontend_io_out_1_bits_cf_exceptionVec_12; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_exceptionVec_12 <= _GEN_440;
        end
      end else begin
        REG__0_cf_exceptionVec_12 <= _GEN_440;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_0 <= _GEN_344;
        end
      end else begin
        REG__0_cf_intrVec_0 <= _GEN_344;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_1 <= _GEN_348;
        end
      end else begin
        REG__0_cf_intrVec_1 <= _GEN_348;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_2 <= _GEN_352;
        end
      end else begin
        REG__0_cf_intrVec_2 <= _GEN_352;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_3 <= _GEN_356;
        end
      end else begin
        REG__0_cf_intrVec_3 <= _GEN_356;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_4 <= _GEN_360;
        end
      end else begin
        REG__0_cf_intrVec_4 <= _GEN_360;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_5 <= _GEN_364;
        end
      end else begin
        REG__0_cf_intrVec_5 <= _GEN_364;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_6 <= _GEN_368;
        end
      end else begin
        REG__0_cf_intrVec_6 <= _GEN_368;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_7 <= _GEN_372;
        end
      end else begin
        REG__0_cf_intrVec_7 <= _GEN_372;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_8 <= _GEN_376;
        end
      end else begin
        REG__0_cf_intrVec_8 <= _GEN_376;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_9 <= _GEN_380;
        end
      end else begin
        REG__0_cf_intrVec_9 <= _GEN_380;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_10 <= _GEN_384;
        end
      end else begin
        REG__0_cf_intrVec_10 <= _GEN_384;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_intrVec_11 <= _GEN_388;
        end
      end else begin
        REG__0_cf_intrVec_11 <= _GEN_388;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_brIdx <= _REG_T_20_cf_brIdx; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_brIdx <= _GEN_340;
        end
      end else begin
        REG__0_cf_brIdx <= _GEN_340;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_cf_crossPageIPFFix <= frontend_io_out_1_bits_cf_crossPageIPFFix; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_cf_crossPageIPFFix <= _GEN_332;
        end
      end else begin
        REG__0_cf_crossPageIPFFix <= _GEN_332;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_src1Type <= frontend_io_out_1_bits_ctrl_src1Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_src1Type <= _GEN_328;
        end
      end else begin
        REG__0_ctrl_src1Type <= _GEN_328;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_src2Type <= frontend_io_out_1_bits_ctrl_src2Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_src2Type <= _GEN_324;
        end
      end else begin
        REG__0_ctrl_src2Type <= _GEN_324;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_fuType <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_fuType <= _REG_T_20_ctrl_fuType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_fuType <= _GEN_320;
        end
      end else begin
        REG__0_ctrl_fuType <= _GEN_320;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_fuOpType <= _REG_T_20_ctrl_fuOpType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_fuOpType <= _GEN_316;
        end
      end else begin
        REG__0_ctrl_fuOpType <= _GEN_316;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_rfSrc1 <= _REG_T_20_ctrl_rfSrc1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_rfSrc1 <= _GEN_312;
        end
      end else begin
        REG__0_ctrl_rfSrc1 <= _GEN_312;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_rfSrc2 <= _REG_T_20_ctrl_rfSrc2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_rfSrc2 <= _GEN_308;
        end
      end else begin
        REG__0_ctrl_rfSrc2 <= _GEN_308;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_rfWen <= frontend_io_out_1_bits_ctrl_rfWen; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_rfWen <= _GEN_304;
        end
      end else begin
        REG__0_ctrl_rfWen <= _GEN_304;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_ctrl_rfDest <= _REG_T_20_ctrl_rfDest; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_ctrl_rfDest <= _GEN_300;
        end
      end else begin
        REG__0_ctrl_rfDest <= _GEN_300;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__0_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h0 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__0_data_imm <= _REG_T_20_data_imm; // @[PipelineVector.scala 46:63]
        end else begin
          REG__0_data_imm <= _GEN_256;
        end
      end else begin
        REG__0_data_imm <= _GEN_256;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_instr <= _REG_T_20_cf_instr; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_instr <= _GEN_501;
        end
      end else begin
        REG__1_cf_instr <= _GEN_501;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_pc <= _REG_T_20_cf_pc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_pc <= _GEN_497;
        end
      end else begin
        REG__1_cf_pc <= _GEN_497;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_pnpc <= _REG_T_20_cf_pnpc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_pnpc <= _GEN_493;
        end
      end else begin
        REG__1_cf_pnpc <= _GEN_493;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_exceptionVec_1 <= frontend_io_out_1_bits_cf_exceptionVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_exceptionVec_1 <= _GEN_397;
        end
      end else begin
        REG__1_cf_exceptionVec_1 <= _GEN_397;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_exceptionVec_2 <= frontend_io_out_1_bits_cf_exceptionVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_exceptionVec_2 <= _GEN_401;
        end
      end else begin
        REG__1_cf_exceptionVec_2 <= _GEN_401;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_exceptionVec_12 <= frontend_io_out_1_bits_cf_exceptionVec_12; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_exceptionVec_12 <= _GEN_441;
        end
      end else begin
        REG__1_cf_exceptionVec_12 <= _GEN_441;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_0 <= _GEN_345;
        end
      end else begin
        REG__1_cf_intrVec_0 <= _GEN_345;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_1 <= _GEN_349;
        end
      end else begin
        REG__1_cf_intrVec_1 <= _GEN_349;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_2 <= _GEN_353;
        end
      end else begin
        REG__1_cf_intrVec_2 <= _GEN_353;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_3 <= _GEN_357;
        end
      end else begin
        REG__1_cf_intrVec_3 <= _GEN_357;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_4 <= _GEN_361;
        end
      end else begin
        REG__1_cf_intrVec_4 <= _GEN_361;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_5 <= _GEN_365;
        end
      end else begin
        REG__1_cf_intrVec_5 <= _GEN_365;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_6 <= _GEN_369;
        end
      end else begin
        REG__1_cf_intrVec_6 <= _GEN_369;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_7 <= _GEN_373;
        end
      end else begin
        REG__1_cf_intrVec_7 <= _GEN_373;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_8 <= _GEN_377;
        end
      end else begin
        REG__1_cf_intrVec_8 <= _GEN_377;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_9 <= _GEN_381;
        end
      end else begin
        REG__1_cf_intrVec_9 <= _GEN_381;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_10 <= _GEN_385;
        end
      end else begin
        REG__1_cf_intrVec_10 <= _GEN_385;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_intrVec_11 <= _GEN_389;
        end
      end else begin
        REG__1_cf_intrVec_11 <= _GEN_389;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_brIdx <= _REG_T_20_cf_brIdx; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_brIdx <= _GEN_341;
        end
      end else begin
        REG__1_cf_brIdx <= _GEN_341;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_cf_crossPageIPFFix <= frontend_io_out_1_bits_cf_crossPageIPFFix; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_cf_crossPageIPFFix <= _GEN_333;
        end
      end else begin
        REG__1_cf_crossPageIPFFix <= _GEN_333;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_src1Type <= frontend_io_out_1_bits_ctrl_src1Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_src1Type <= _GEN_329;
        end
      end else begin
        REG__1_ctrl_src1Type <= _GEN_329;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_src2Type <= frontend_io_out_1_bits_ctrl_src2Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_src2Type <= _GEN_325;
        end
      end else begin
        REG__1_ctrl_src2Type <= _GEN_325;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_fuType <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_fuType <= _REG_T_20_ctrl_fuType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_fuType <= _GEN_321;
        end
      end else begin
        REG__1_ctrl_fuType <= _GEN_321;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_fuOpType <= _REG_T_20_ctrl_fuOpType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_fuOpType <= _GEN_317;
        end
      end else begin
        REG__1_ctrl_fuOpType <= _GEN_317;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_rfSrc1 <= _REG_T_20_ctrl_rfSrc1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_rfSrc1 <= _GEN_313;
        end
      end else begin
        REG__1_ctrl_rfSrc1 <= _GEN_313;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_rfSrc2 <= _REG_T_20_ctrl_rfSrc2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_rfSrc2 <= _GEN_309;
        end
      end else begin
        REG__1_ctrl_rfSrc2 <= _GEN_309;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_rfWen <= frontend_io_out_1_bits_ctrl_rfWen; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_rfWen <= _GEN_305;
        end
      end else begin
        REG__1_ctrl_rfWen <= _GEN_305;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_ctrl_rfDest <= _REG_T_20_ctrl_rfDest; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_ctrl_rfDest <= _GEN_301;
        end
      end else begin
        REG__1_ctrl_rfDest <= _GEN_301;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__1_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h1 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__1_data_imm <= _REG_T_20_data_imm; // @[PipelineVector.scala 46:63]
        end else begin
          REG__1_data_imm <= _GEN_257;
        end
      end else begin
        REG__1_data_imm <= _GEN_257;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_instr <= _REG_T_20_cf_instr; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_instr <= _GEN_502;
        end
      end else begin
        REG__2_cf_instr <= _GEN_502;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_pc <= _REG_T_20_cf_pc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_pc <= _GEN_498;
        end
      end else begin
        REG__2_cf_pc <= _GEN_498;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_pnpc <= _REG_T_20_cf_pnpc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_pnpc <= _GEN_494;
        end
      end else begin
        REG__2_cf_pnpc <= _GEN_494;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_exceptionVec_1 <= frontend_io_out_1_bits_cf_exceptionVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_exceptionVec_1 <= _GEN_398;
        end
      end else begin
        REG__2_cf_exceptionVec_1 <= _GEN_398;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_exceptionVec_2 <= frontend_io_out_1_bits_cf_exceptionVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_exceptionVec_2 <= _GEN_402;
        end
      end else begin
        REG__2_cf_exceptionVec_2 <= _GEN_402;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_exceptionVec_12 <= frontend_io_out_1_bits_cf_exceptionVec_12; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_exceptionVec_12 <= _GEN_442;
        end
      end else begin
        REG__2_cf_exceptionVec_12 <= _GEN_442;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_0 <= _GEN_346;
        end
      end else begin
        REG__2_cf_intrVec_0 <= _GEN_346;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_1 <= _GEN_350;
        end
      end else begin
        REG__2_cf_intrVec_1 <= _GEN_350;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_2 <= _GEN_354;
        end
      end else begin
        REG__2_cf_intrVec_2 <= _GEN_354;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_3 <= _GEN_358;
        end
      end else begin
        REG__2_cf_intrVec_3 <= _GEN_358;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_4 <= _GEN_362;
        end
      end else begin
        REG__2_cf_intrVec_4 <= _GEN_362;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_5 <= _GEN_366;
        end
      end else begin
        REG__2_cf_intrVec_5 <= _GEN_366;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_6 <= _GEN_370;
        end
      end else begin
        REG__2_cf_intrVec_6 <= _GEN_370;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_7 <= _GEN_374;
        end
      end else begin
        REG__2_cf_intrVec_7 <= _GEN_374;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_8 <= _GEN_378;
        end
      end else begin
        REG__2_cf_intrVec_8 <= _GEN_378;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_9 <= _GEN_382;
        end
      end else begin
        REG__2_cf_intrVec_9 <= _GEN_382;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_10 <= _GEN_386;
        end
      end else begin
        REG__2_cf_intrVec_10 <= _GEN_386;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_intrVec_11 <= _GEN_390;
        end
      end else begin
        REG__2_cf_intrVec_11 <= _GEN_390;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_brIdx <= _REG_T_20_cf_brIdx; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_brIdx <= _GEN_342;
        end
      end else begin
        REG__2_cf_brIdx <= _GEN_342;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_cf_crossPageIPFFix <= frontend_io_out_1_bits_cf_crossPageIPFFix; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_cf_crossPageIPFFix <= _GEN_334;
        end
      end else begin
        REG__2_cf_crossPageIPFFix <= _GEN_334;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_src1Type <= frontend_io_out_1_bits_ctrl_src1Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_src1Type <= _GEN_330;
        end
      end else begin
        REG__2_ctrl_src1Type <= _GEN_330;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_src2Type <= frontend_io_out_1_bits_ctrl_src2Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_src2Type <= _GEN_326;
        end
      end else begin
        REG__2_ctrl_src2Type <= _GEN_326;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_fuType <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_fuType <= _REG_T_20_ctrl_fuType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_fuType <= _GEN_322;
        end
      end else begin
        REG__2_ctrl_fuType <= _GEN_322;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_fuOpType <= _REG_T_20_ctrl_fuOpType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_fuOpType <= _GEN_318;
        end
      end else begin
        REG__2_ctrl_fuOpType <= _GEN_318;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_rfSrc1 <= _REG_T_20_ctrl_rfSrc1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_rfSrc1 <= _GEN_314;
        end
      end else begin
        REG__2_ctrl_rfSrc1 <= _GEN_314;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_rfSrc2 <= _REG_T_20_ctrl_rfSrc2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_rfSrc2 <= _GEN_310;
        end
      end else begin
        REG__2_ctrl_rfSrc2 <= _GEN_310;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_rfWen <= frontend_io_out_1_bits_ctrl_rfWen; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_rfWen <= _GEN_306;
        end
      end else begin
        REG__2_ctrl_rfWen <= _GEN_306;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_ctrl_rfDest <= _REG_T_20_ctrl_rfDest; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_ctrl_rfDest <= _GEN_302;
        end
      end else begin
        REG__2_ctrl_rfDest <= _GEN_302;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__2_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h2 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__2_data_imm <= _REG_T_20_data_imm; // @[PipelineVector.scala 46:63]
        end else begin
          REG__2_data_imm <= _GEN_258;
        end
      end else begin
        REG__2_data_imm <= _GEN_258;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_instr <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_instr <= _REG_T_20_cf_instr; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_instr <= _GEN_503;
        end
      end else begin
        REG__3_cf_instr <= _GEN_503;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_pc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_pc <= _REG_T_20_cf_pc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_pc <= _GEN_499;
        end
      end else begin
        REG__3_cf_pc <= _GEN_499;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_pnpc <= 39'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_pnpc <= _REG_T_20_cf_pnpc; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_pnpc <= _GEN_495;
        end
      end else begin
        REG__3_cf_pnpc <= _GEN_495;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_exceptionVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_exceptionVec_1 <= frontend_io_out_1_bits_cf_exceptionVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_exceptionVec_1 <= _GEN_399;
        end
      end else begin
        REG__3_cf_exceptionVec_1 <= _GEN_399;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_exceptionVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_exceptionVec_2 <= frontend_io_out_1_bits_cf_exceptionVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_exceptionVec_2 <= _GEN_403;
        end
      end else begin
        REG__3_cf_exceptionVec_2 <= _GEN_403;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_exceptionVec_12 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_exceptionVec_12 <= frontend_io_out_1_bits_cf_exceptionVec_12; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_exceptionVec_12 <= _GEN_443;
        end
      end else begin
        REG__3_cf_exceptionVec_12 <= _GEN_443;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_0 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_0 <= _GEN_347;
        end
      end else begin
        REG__3_cf_intrVec_0 <= _GEN_347;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_1 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_1 <= _GEN_351;
        end
      end else begin
        REG__3_cf_intrVec_1 <= _GEN_351;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_2 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_2 <= _GEN_355;
        end
      end else begin
        REG__3_cf_intrVec_2 <= _GEN_355;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_3 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_3 <= _GEN_359;
        end
      end else begin
        REG__3_cf_intrVec_3 <= _GEN_359;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_4 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_4 <= _GEN_363;
        end
      end else begin
        REG__3_cf_intrVec_4 <= _GEN_363;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_5 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_5 <= _GEN_367;
        end
      end else begin
        REG__3_cf_intrVec_5 <= _GEN_367;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_6 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_6 <= _GEN_371;
        end
      end else begin
        REG__3_cf_intrVec_6 <= _GEN_371;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_7 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_7 <= _GEN_375;
        end
      end else begin
        REG__3_cf_intrVec_7 <= _GEN_375;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_8 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_8 <= _GEN_379;
        end
      end else begin
        REG__3_cf_intrVec_8 <= _GEN_379;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_9 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_9 <= _GEN_383;
        end
      end else begin
        REG__3_cf_intrVec_9 <= _GEN_383;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_10 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_10 <= _GEN_387;
        end
      end else begin
        REG__3_cf_intrVec_10 <= _GEN_387;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_intrVec_11 <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_intrVec_11 <= _GEN_391;
        end
      end else begin
        REG__3_cf_intrVec_11 <= _GEN_391;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_brIdx <= 4'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_brIdx <= _REG_T_20_cf_brIdx; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_brIdx <= _GEN_343;
        end
      end else begin
        REG__3_cf_brIdx <= _GEN_343;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_cf_crossPageIPFFix <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_cf_crossPageIPFFix <= frontend_io_out_1_bits_cf_crossPageIPFFix; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_cf_crossPageIPFFix <= _GEN_335;
        end
      end else begin
        REG__3_cf_crossPageIPFFix <= _GEN_335;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_src1Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_src1Type <= frontend_io_out_1_bits_ctrl_src1Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_src1Type <= _GEN_331;
        end
      end else begin
        REG__3_ctrl_src1Type <= _GEN_331;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_src2Type <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_src2Type <= frontend_io_out_1_bits_ctrl_src2Type; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_src2Type <= _GEN_327;
        end
      end else begin
        REG__3_ctrl_src2Type <= _GEN_327;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_fuType <= 3'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_fuType <= _REG_T_20_ctrl_fuType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_fuType <= _GEN_323;
        end
      end else begin
        REG__3_ctrl_fuType <= _GEN_323;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_fuOpType <= 7'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_fuOpType <= _REG_T_20_ctrl_fuOpType; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_fuOpType <= _GEN_319;
        end
      end else begin
        REG__3_ctrl_fuOpType <= _GEN_319;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_rfSrc1 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_rfSrc1 <= _REG_T_20_ctrl_rfSrc1; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_rfSrc1 <= _GEN_315;
        end
      end else begin
        REG__3_ctrl_rfSrc1 <= _GEN_315;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_rfSrc2 <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_rfSrc2 <= _REG_T_20_ctrl_rfSrc2; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_rfSrc2 <= _GEN_311;
        end
      end else begin
        REG__3_ctrl_rfSrc2 <= _GEN_311;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_rfWen <= 1'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_rfWen <= frontend_io_out_1_bits_ctrl_rfWen; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_rfWen <= _GEN_307;
        end
      end else begin
        REG__3_ctrl_rfWen <= _GEN_307;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_ctrl_rfDest <= 5'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_ctrl_rfDest <= _REG_T_20_ctrl_rfDest; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_ctrl_rfDest <= _GEN_303;
        end
      end else begin
        REG__3_ctrl_rfDest <= _GEN_303;
      end
    end
    if (reset) begin // @[PipelineVector.scala 29:29]
      REG__3_data_imm <= 64'h0; // @[PipelineVector.scala 29:29]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      if (_T_12) begin // @[PipelineVector.scala 46:29]
        if (2'h3 == _T_20) begin // @[PipelineVector.scala 46:63]
          REG__3_data_imm <= _REG_T_20_data_imm; // @[PipelineVector.scala 46:63]
        end else begin
          REG__3_data_imm <= _GEN_259;
        end
      end else begin
        REG__3_data_imm <= _GEN_259;
      end
    end
    if (reset) begin // @[PipelineVector.scala 30:33]
      REG_1 <= 2'h0; // @[PipelineVector.scala 30:33]
    end else if (frontend_io_flushVec[1]) begin // @[PipelineVector.scala 71:16]
      REG_1 <= 2'h0; // @[PipelineVector.scala 72:24]
    end else if (_T_15) begin // @[PipelineVector.scala 44:14]
      REG_1 <= _T_22; // @[PipelineVector.scala 47:24]
    end
    if (reset) begin // @[PipelineVector.scala 31:33]
      REG_2 <= 2'h0; // @[PipelineVector.scala 31:33]
    end else if (frontend_io_flushVec[1]) begin // @[PipelineVector.scala 71:16]
      REG_2 <= 2'h0; // @[PipelineVector.scala 73:24]
    end else if (_T_35) begin // @[PipelineVector.scala 66:22]
      REG_2 <= _T_37; // @[PipelineVector.scala 67:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  REG__0_cf_instr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  REG__0_cf_pc = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  REG__0_cf_pnpc = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  REG__0_cf_exceptionVec_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG__0_cf_exceptionVec_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG__0_cf_exceptionVec_12 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  REG__0_cf_intrVec_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  REG__0_cf_intrVec_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  REG__0_cf_intrVec_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  REG__0_cf_intrVec_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  REG__0_cf_intrVec_4 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG__0_cf_intrVec_5 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  REG__0_cf_intrVec_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  REG__0_cf_intrVec_7 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  REG__0_cf_intrVec_8 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  REG__0_cf_intrVec_9 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  REG__0_cf_intrVec_10 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  REG__0_cf_intrVec_11 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  REG__0_cf_brIdx = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  REG__0_cf_crossPageIPFFix = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  REG__0_ctrl_src1Type = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  REG__0_ctrl_src2Type = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  REG__0_ctrl_fuType = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  REG__0_ctrl_fuOpType = _RAND_23[6:0];
  _RAND_24 = {1{`RANDOM}};
  REG__0_ctrl_rfSrc1 = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  REG__0_ctrl_rfSrc2 = _RAND_25[4:0];
  _RAND_26 = {1{`RANDOM}};
  REG__0_ctrl_rfWen = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  REG__0_ctrl_rfDest = _RAND_27[4:0];
  _RAND_28 = {2{`RANDOM}};
  REG__0_data_imm = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  REG__1_cf_instr = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  REG__1_cf_pc = _RAND_30[38:0];
  _RAND_31 = {2{`RANDOM}};
  REG__1_cf_pnpc = _RAND_31[38:0];
  _RAND_32 = {1{`RANDOM}};
  REG__1_cf_exceptionVec_1 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  REG__1_cf_exceptionVec_2 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  REG__1_cf_exceptionVec_12 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  REG__1_cf_intrVec_0 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  REG__1_cf_intrVec_1 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  REG__1_cf_intrVec_2 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  REG__1_cf_intrVec_3 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  REG__1_cf_intrVec_4 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  REG__1_cf_intrVec_5 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  REG__1_cf_intrVec_6 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  REG__1_cf_intrVec_7 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  REG__1_cf_intrVec_8 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  REG__1_cf_intrVec_9 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  REG__1_cf_intrVec_10 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  REG__1_cf_intrVec_11 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  REG__1_cf_brIdx = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  REG__1_cf_crossPageIPFFix = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  REG__1_ctrl_src1Type = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  REG__1_ctrl_src2Type = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  REG__1_ctrl_fuType = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  REG__1_ctrl_fuOpType = _RAND_52[6:0];
  _RAND_53 = {1{`RANDOM}};
  REG__1_ctrl_rfSrc1 = _RAND_53[4:0];
  _RAND_54 = {1{`RANDOM}};
  REG__1_ctrl_rfSrc2 = _RAND_54[4:0];
  _RAND_55 = {1{`RANDOM}};
  REG__1_ctrl_rfWen = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  REG__1_ctrl_rfDest = _RAND_56[4:0];
  _RAND_57 = {2{`RANDOM}};
  REG__1_data_imm = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  REG__2_cf_instr = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  REG__2_cf_pc = _RAND_59[38:0];
  _RAND_60 = {2{`RANDOM}};
  REG__2_cf_pnpc = _RAND_60[38:0];
  _RAND_61 = {1{`RANDOM}};
  REG__2_cf_exceptionVec_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  REG__2_cf_exceptionVec_2 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  REG__2_cf_exceptionVec_12 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  REG__2_cf_intrVec_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  REG__2_cf_intrVec_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  REG__2_cf_intrVec_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  REG__2_cf_intrVec_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  REG__2_cf_intrVec_4 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  REG__2_cf_intrVec_5 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  REG__2_cf_intrVec_6 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  REG__2_cf_intrVec_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  REG__2_cf_intrVec_8 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  REG__2_cf_intrVec_9 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  REG__2_cf_intrVec_10 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  REG__2_cf_intrVec_11 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  REG__2_cf_brIdx = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  REG__2_cf_crossPageIPFFix = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  REG__2_ctrl_src1Type = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  REG__2_ctrl_src2Type = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  REG__2_ctrl_fuType = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  REG__2_ctrl_fuOpType = _RAND_81[6:0];
  _RAND_82 = {1{`RANDOM}};
  REG__2_ctrl_rfSrc1 = _RAND_82[4:0];
  _RAND_83 = {1{`RANDOM}};
  REG__2_ctrl_rfSrc2 = _RAND_83[4:0];
  _RAND_84 = {1{`RANDOM}};
  REG__2_ctrl_rfWen = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  REG__2_ctrl_rfDest = _RAND_85[4:0];
  _RAND_86 = {2{`RANDOM}};
  REG__2_data_imm = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  REG__3_cf_instr = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  REG__3_cf_pc = _RAND_88[38:0];
  _RAND_89 = {2{`RANDOM}};
  REG__3_cf_pnpc = _RAND_89[38:0];
  _RAND_90 = {1{`RANDOM}};
  REG__3_cf_exceptionVec_1 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  REG__3_cf_exceptionVec_2 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  REG__3_cf_exceptionVec_12 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  REG__3_cf_intrVec_0 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  REG__3_cf_intrVec_1 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  REG__3_cf_intrVec_2 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  REG__3_cf_intrVec_3 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  REG__3_cf_intrVec_4 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  REG__3_cf_intrVec_5 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  REG__3_cf_intrVec_6 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  REG__3_cf_intrVec_7 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  REG__3_cf_intrVec_8 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  REG__3_cf_intrVec_9 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  REG__3_cf_intrVec_10 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  REG__3_cf_intrVec_11 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  REG__3_cf_brIdx = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  REG__3_cf_crossPageIPFFix = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  REG__3_ctrl_src1Type = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  REG__3_ctrl_src2Type = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  REG__3_ctrl_fuType = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  REG__3_ctrl_fuOpType = _RAND_110[6:0];
  _RAND_111 = {1{`RANDOM}};
  REG__3_ctrl_rfSrc1 = _RAND_111[4:0];
  _RAND_112 = {1{`RANDOM}};
  REG__3_ctrl_rfSrc2 = _RAND_112[4:0];
  _RAND_113 = {1{`RANDOM}};
  REG__3_ctrl_rfWen = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  REG__3_ctrl_rfDest = _RAND_114[4:0];
  _RAND_115 = {2{`RANDOM}};
  REG__3_data_imm = _RAND_115[63:0];
  _RAND_116 = {1{`RANDOM}};
  REG_1 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  REG_2 = _RAND_117[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_CoherenceManager(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [2:0]  io_out_mem_req_bits_size,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [7:0]  io_out_mem_req_bits_wmask,
  output [63:0] io_out_mem_req_bits_wdata,
  output        io_out_mem_resp_ready,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  input         io_out_coh_req_ready,
  output        io_out_coh_req_valid,
  output [31:0] io_out_coh_req_bits_addr,
  output [63:0] io_out_coh_req_bits_wdata,
  output        io_out_coh_resp_ready,
  input         io_out_coh_resp_valid,
  input  [3:0]  io_out_coh_resp_bits_cmd,
  input  [63:0] io_out_coh_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Coherence.scala 45:22]
  wire  inflight = state != 3'h0; // @[Coherence.scala 46:24]
  wire  _T_1 = ~io_in_req_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_4 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_14 = ~inflight; // @[Coherence.scala 52:70]
  wire  _T_20 = ~inflight & _T_4; // @[Coherence.scala 52:80]
  reg [31:0] reqLatch_addr; // @[Reg.scala 27:20]
  reg [2:0] reqLatch_size; // @[Reg.scala 27:20]
  reg [3:0] reqLatch_cmd; // @[Reg.scala 27:20]
  reg [7:0] reqLatch_wmask; // @[Reg.scala 27:20]
  reg [63:0] reqLatch_wdata; // @[Reg.scala 27:20]
  wire  _T_23 = io_in_req_valid & _T_14; // @[Coherence.scala 65:43]
  wire  _GEN_5 = _T_4 & _T_23; // @[Coherence.scala 67:39 Coherence.scala 68:26 Coherence.scala 63:24]
  wire  _GEN_6 = _T_4 & (io_out_coh_req_ready & _T_14); // @[Coherence.scala 67:39 Coherence.scala 69:19 Coherence.scala 62:17]
  wire  _GEN_7 = io_in_req_bits_cmd[0] & (io_in_req_valid & _T_14); // @[Coherence.scala 64:61 Coherence.scala 65:26 Coherence.scala 61:24]
  wire  _T_35 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_36 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_43 = io_in_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire [2:0] _GEN_10 = _T_43 ? 3'h5 : state; // @[Coherence.scala 78:48 Coherence.scala 78:56 Coherence.scala 45:22]
  wire  _T_44 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_45 = io_out_coh_resp_ready & io_out_coh_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_46 = io_out_coh_resp_bits_cmd == 4'hc; // @[SimpleBus.scala 92:26]
  wire [2:0] _T_47 = _T_46 ? 3'h2 : 3'h3; // @[Coherence.scala 83:21]
  wire  _T_48 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_50 = io_in_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [2:0] _GEN_14 = io_in_resp_valid & _T_50 ? 3'h0 : state; // @[Coherence.scala 89:60 Coherence.scala 89:68 Coherence.scala 45:22]
  wire  _T_52 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_53 = io_out_mem_req_ready & io_out_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_15 = _T_53 ? 3'h4 : state; // @[Coherence.scala 94:36 Coherence.scala 94:44 Coherence.scala 45:22]
  wire  _T_54 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_55 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_56 = io_out_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire [2:0] _GEN_16 = _T_55 & _T_56 ? 3'h0 : state; // @[Coherence.scala 96:93 Coherence.scala 96:101 Coherence.scala 45:22]
  wire  _T_58 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_17 = _T_55 ? 3'h0 : state; // @[Coherence.scala 97:57 Coherence.scala 97:65 Coherence.scala 45:22]
  wire [2:0] _GEN_18 = _T_58 ? _GEN_17 : state; // @[Conditional.scala 39:67 Coherence.scala 45:22]
  wire [2:0] _GEN_19 = _T_54 ? _GEN_16 : _GEN_18; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_20 = _T_52 ? reqLatch_wdata : io_in_req_bits_wdata; // @[Conditional.scala 39:67 Coherence.scala 92:27 Coherence.scala 59:23]
  wire [7:0] _GEN_21 = _T_52 ? reqLatch_wmask : 8'hff; // @[Conditional.scala 39:67 Coherence.scala 92:27 Coherence.scala 59:23]
  wire [3:0] _GEN_22 = _T_52 ? reqLatch_cmd : io_in_req_bits_cmd; // @[Conditional.scala 39:67 Coherence.scala 92:27 Coherence.scala 59:23]
  wire [2:0] _GEN_23 = _T_52 ? reqLatch_size : 3'h3; // @[Conditional.scala 39:67 Coherence.scala 92:27 Coherence.scala 59:23]
  wire [31:0] _GEN_24 = _T_52 ? reqLatch_addr : io_in_req_bits_addr; // @[Conditional.scala 39:67 Coherence.scala 92:27 Coherence.scala 59:23]
  wire  _GEN_25 = _T_52 | _GEN_7; // @[Conditional.scala 39:67 Coherence.scala 93:28]
  wire [2:0] _GEN_26 = _T_52 ? _GEN_15 : _GEN_19; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_27 = _T_48 ? io_out_coh_resp_bits_rdata : io_out_mem_resp_bits_rdata; // @[Conditional.scala 39:67 Coherence.scala 88:16 Coherence.scala 72:14]
  wire [3:0] _GEN_28 = _T_48 ? io_out_coh_resp_bits_cmd : io_out_mem_resp_bits_cmd; // @[Conditional.scala 39:67 Coherence.scala 88:16 Coherence.scala 72:14]
  wire  _GEN_29 = _T_48 ? io_out_coh_resp_valid : io_out_mem_resp_valid; // @[Conditional.scala 39:67 Coherence.scala 88:16 Coherence.scala 72:14]
  wire [63:0] _GEN_32 = _T_48 ? io_in_req_bits_wdata : _GEN_20; // @[Conditional.scala 39:67 Coherence.scala 59:23]
  wire [7:0] _GEN_33 = _T_48 ? 8'hff : _GEN_21; // @[Conditional.scala 39:67 Coherence.scala 59:23]
  wire [3:0] _GEN_34 = _T_48 ? io_in_req_bits_cmd : _GEN_22; // @[Conditional.scala 39:67 Coherence.scala 59:23]
  wire [2:0] _GEN_35 = _T_48 ? 3'h3 : _GEN_23; // @[Conditional.scala 39:67 Coherence.scala 59:23]
  wire [31:0] _GEN_36 = _T_48 ? io_in_req_bits_addr : _GEN_24; // @[Conditional.scala 39:67 Coherence.scala 59:23]
  wire  _GEN_37 = _T_48 ? _GEN_7 : _GEN_25; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_39 = _T_44 ? io_out_mem_resp_bits_rdata : _GEN_27; // @[Conditional.scala 39:67 Coherence.scala 72:14]
  wire [3:0] _GEN_40 = _T_44 ? io_out_mem_resp_bits_cmd : _GEN_28; // @[Conditional.scala 39:67 Coherence.scala 72:14]
  wire  _GEN_41 = _T_44 ? io_out_mem_resp_valid : _GEN_29; // @[Conditional.scala 39:67 Coherence.scala 72:14]
  wire [63:0] _GEN_43 = _T_44 ? io_in_req_bits_wdata : _GEN_32; // @[Conditional.scala 39:67 Coherence.scala 59:23]
  wire [7:0] _GEN_44 = _T_44 ? 8'hff : _GEN_33; // @[Conditional.scala 39:67 Coherence.scala 59:23]
  wire [3:0] _GEN_45 = _T_44 ? io_in_req_bits_cmd : _GEN_34; // @[Conditional.scala 39:67 Coherence.scala 59:23]
  wire [2:0] _GEN_46 = _T_44 ? 3'h3 : _GEN_35; // @[Conditional.scala 39:67 Coherence.scala 59:23]
  wire [31:0] _GEN_47 = _T_44 ? io_in_req_bits_addr : _GEN_36; // @[Conditional.scala 39:67 Coherence.scala 59:23]
  wire  _GEN_48 = _T_44 ? _GEN_7 : _GEN_37; // @[Conditional.scala 39:67]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? io_out_mem_req_ready & _T_14 : _GEN_6; // @[Coherence.scala 64:61 Coherence.scala 66:19]
  assign io_in_resp_valid = _T_35 ? io_out_mem_resp_valid : _GEN_41; // @[Conditional.scala 40:58 Coherence.scala 72:14]
  assign io_in_resp_bits_cmd = _T_35 ? io_out_mem_resp_bits_cmd : _GEN_40; // @[Conditional.scala 40:58 Coherence.scala 72:14]
  assign io_in_resp_bits_rdata = _T_35 ? io_out_mem_resp_bits_rdata : _GEN_39; // @[Conditional.scala 40:58 Coherence.scala 72:14]
  assign io_out_mem_req_valid = _T_35 ? _GEN_7 : _GEN_48; // @[Conditional.scala 40:58]
  assign io_out_mem_req_bits_addr = _T_35 ? io_in_req_bits_addr : _GEN_47; // @[Conditional.scala 40:58 Coherence.scala 59:23]
  assign io_out_mem_req_bits_size = _T_35 ? 3'h3 : _GEN_46; // @[Conditional.scala 40:58 Coherence.scala 59:23]
  assign io_out_mem_req_bits_cmd = _T_35 ? io_in_req_bits_cmd : _GEN_45; // @[Conditional.scala 40:58 Coherence.scala 59:23]
  assign io_out_mem_req_bits_wmask = _T_35 ? 8'hff : _GEN_44; // @[Conditional.scala 40:58 Coherence.scala 59:23]
  assign io_out_mem_req_bits_wdata = _T_35 ? io_in_req_bits_wdata : _GEN_43; // @[Conditional.scala 40:58 Coherence.scala 59:23]
  assign io_out_mem_resp_ready = 1'h1; // @[Coherence.scala 72:14]
  assign io_out_coh_req_valid = io_in_req_bits_cmd[0] ? 1'h0 : _GEN_5; // @[Coherence.scala 64:61 Coherence.scala 63:24]
  assign io_out_coh_req_bits_addr = io_in_req_bits_addr; // @[Coherence.scala 54:16]
  assign io_out_coh_req_bits_wdata = io_in_req_bits_wdata; // @[Coherence.scala 54:16]
  assign io_out_coh_resp_ready = 1'h1; // @[Conditional.scala 40:58 Coherence.scala 56:18]
  always @(posedge clock) begin
    if (reset) begin // @[Coherence.scala 45:22]
      state <= 3'h0; // @[Coherence.scala 45:22]
    end else if (_T_35) begin // @[Conditional.scala 40:58]
      if (_T_36) begin // @[Coherence.scala 76:29]
        if (_T_4) begin // @[Coherence.scala 77:38]
          state <= 3'h1; // @[Coherence.scala 77:46]
        end else begin
          state <= _GEN_10;
        end
      end
    end else if (_T_44) begin // @[Conditional.scala 39:67]
      if (_T_45) begin // @[Coherence.scala 82:37]
        state <= _T_47; // @[Coherence.scala 83:15]
      end
    end else if (_T_48) begin // @[Conditional.scala 39:67]
      state <= _GEN_14;
    end else begin
      state <= _GEN_26;
    end
    if (reset) begin // @[Reg.scala 27:20]
      reqLatch_addr <= 32'h0; // @[Reg.scala 27:20]
    end else if (_T_20) begin // @[Reg.scala 28:19]
      reqLatch_addr <= io_in_req_bits_addr; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reqLatch_size <= 3'h0; // @[Reg.scala 27:20]
    end else if (_T_20) begin // @[Reg.scala 28:19]
      reqLatch_size <= 3'h3; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reqLatch_cmd <= 4'h0; // @[Reg.scala 27:20]
    end else if (_T_20) begin // @[Reg.scala 28:19]
      reqLatch_cmd <= io_in_req_bits_cmd; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reqLatch_wmask <= 8'h0; // @[Reg.scala 27:20]
    end else if (_T_20) begin // @[Reg.scala 28:19]
      reqLatch_wmask <= 8'hff; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      reqLatch_wdata <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_20) begin // @[Reg.scala 28:19]
      reqLatch_wdata <= io_in_req_bits_wdata; // @[Reg.scala 28:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~(io_in_req_valid & ~_T_4 & _T_1) | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Coherence.scala:49 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"
            ); // @[Coherence.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~(io_in_req_valid & ~_T_4 & _T_1) | reset)) begin
          $fatal; // @[Coherence.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  reqLatch_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reqLatch_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  reqLatch_cmd = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  reqLatch_wmask = _RAND_4[7:0];
  _RAND_5 = {2{`RANDOM}};
  reqLatch_wdata = _RAND_5[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_AXI42SimpleBusConverter(
  input         clock,
  input         reset,
  output        io_in_awready,
  input         io_in_awvalid,
  input  [31:0] io_in_awaddr,
  input  [17:0] io_in_awid,
  input  [7:0]  io_in_awlen,
  input  [2:0]  io_in_awsize,
  output        io_in_wready,
  input         io_in_wvalid,
  input  [63:0] io_in_wdata,
  input  [7:0]  io_in_wstrb,
  input         io_in_wlast,
  input         io_in_bready,
  output        io_in_bvalid,
  output        io_in_arready,
  input         io_in_arvalid,
  input  [31:0] io_in_araddr,
  input  [17:0] io_in_arid,
  input  [7:0]  io_in_arlen,
  input  [2:0]  io_in_arsize,
  input         io_in_rready,
  output        io_in_rvalid,
  output [63:0] io_in_rdata,
  output        io_in_rlast,
  output [17:0] io_in_rid,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [17:0] inflight_id_reg; // @[ToAXI4.scala 38:32]
  reg [1:0] inflight_type; // @[ToAXI4.scala 40:30]
  wire  _T = inflight_type == 2'h0; // @[ToAXI4.scala 50:19]
  wire  _T_1 = ~_T; // @[ToAXI4.scala 53:5]
  wire  _T_2 = ~_T_1; // @[ToAXI4.scala 64:9]
  wire  _T_3 = ~_T_1 & io_in_arvalid; // @[ToAXI4.scala 64:23]
  wire [1:0] _T_5 = io_in_arlen == 8'h0 ? 2'h0 : 2'h2; // @[ToAXI4.scala 67:19]
  wire  _T_6 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire [17:0] _GEN_0 = _T_6 ? io_in_arid : inflight_id_reg; // @[ToAXI4.scala 74:25 ToAXI4.scala 42:21 ToAXI4.scala 38:32]
  wire [1:0] _GEN_1 = _T_6 ? 2'h1 : inflight_type; // @[ToAXI4.scala 74:25 ToAXI4.scala 43:19 ToAXI4.scala 40:30]
  wire [31:0] _GEN_2 = ~_T_1 & io_in_arvalid ? io_in_araddr : 32'h0; // @[ToAXI4.scala 64:40 ToAXI4.scala 66:14 ToAXI4.scala 59:7]
  wire [3:0] _GEN_3 = ~_T_1 & io_in_arvalid ? {{2'd0}, _T_5} : 4'h0; // @[ToAXI4.scala 64:40 ToAXI4.scala 67:13 ToAXI4.scala 59:7]
  wire [2:0] _GEN_4 = ~_T_1 & io_in_arvalid ? io_in_arsize : 3'h0; // @[ToAXI4.scala 64:40 ToAXI4.scala 69:14 ToAXI4.scala 59:7]
  wire [17:0] _GEN_7 = ~_T_1 & io_in_arvalid ? _GEN_0 : inflight_id_reg; // @[ToAXI4.scala 64:40 ToAXI4.scala 38:32]
  wire [1:0] _GEN_8 = ~_T_1 & io_in_arvalid ? _GEN_1 : inflight_type; // @[ToAXI4.scala 64:40 ToAXI4.scala 40:30]
  wire  _T_7 = inflight_type == 2'h1; // @[ToAXI4.scala 50:19]
  wire  _T_9 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_10 = io_in_rready & io_in_rvalid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_9 = _T_10 & _T_9 ? 2'h0 : _GEN_8; // @[ToAXI4.scala 88:42 ToAXI4.scala 46:19]
  wire [17:0] _GEN_10 = _T_10 & _T_9 ? 18'h0 : _GEN_7; // @[ToAXI4.scala 88:42 ToAXI4.scala 47:21]
  wire [1:0] _GEN_15 = _T_7 & io_out_resp_valid ? _GEN_9 : _GEN_8; // @[ToAXI4.scala 79:46]
  wire [17:0] _GEN_16 = _T_7 & io_out_resp_valid ? _GEN_10 : _GEN_7; // @[ToAXI4.scala 79:46]
  reg [31:0] aw_reg_addr; // @[ToAXI4.scala 94:23]
  reg [7:0] aw_reg_len; // @[ToAXI4.scala 94:23]
  reg [2:0] aw_reg_size; // @[ToAXI4.scala 94:23]
  reg  bresp_en; // @[ToAXI4.scala 95:25]
  wire  _T_17 = ~io_in_arvalid; // @[ToAXI4.scala 97:42]
  wire  _T_19 = io_in_awready & io_in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_20 = inflight_type == 2'h2; // @[ToAXI4.scala 50:19]
  wire  _T_21 = io_in_wready & io_in_wvalid; // @[Decoupled.scala 40:37]
  wire [2:0] _T_24 = io_in_wlast ? 3'h7 : 3'h3; // @[ToAXI4.scala 108:10]
  wire [2:0] _T_25 = aw_reg_len == 8'h0 ? 3'h1 : _T_24; // @[ToAXI4.scala 107:19]
  wire  _GEN_27 = io_in_wlast | bresp_en; // @[ToAXI4.scala 115:19 ToAXI4.scala 116:16 ToAXI4.scala 95:25]
  wire  _T_26 = io_in_bready & io_in_bvalid; // @[Decoupled.scala 40:37]
  wire  _T_57 = io_in_arready & io_in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_81 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  assign io_in_awready = _T_2 & _T_17; // @[ToAXI4.scala 132:33]
  assign io_in_wready = _T_20 & io_out_req_ready; // @[ToAXI4.scala 133:38]
  assign io_in_bvalid = bresp_en & io_out_resp_valid; // @[ToAXI4.scala 134:27]
  assign io_in_arready = _T_2 & io_out_req_ready; // @[ToAXI4.scala 129:33]
  assign io_in_rvalid = _T_7 & io_out_resp_valid; // @[ToAXI4.scala 130:36]
  assign io_in_rdata = _T_7 & io_out_resp_valid ? io_out_resp_bits_rdata : 64'h0; // @[ToAXI4.scala 79:46 ToAXI4.scala 81:12 ToAXI4.scala 60:5]
  assign io_in_rlast = _T_7 & io_out_resp_valid & _T_9; // @[ToAXI4.scala 79:46 ToAXI4.scala 85:12 ToAXI4.scala 60:5]
  assign io_in_rid = _T_7 & io_out_resp_valid ? inflight_id_reg : 18'h0; // @[ToAXI4.scala 79:46 ToAXI4.scala 82:10 ToAXI4.scala 60:5]
  assign io_out_req_valid = _T_3 | _T_20 & io_in_wvalid; // @[ToAXI4.scala 127:52]
  assign io_out_req_bits_addr = _T_20 & _T_21 ? aw_reg_addr : _GEN_2; // @[ToAXI4.scala 105:45 ToAXI4.scala 109:14]
  assign io_out_req_bits_size = _T_20 & _T_21 ? aw_reg_size : _GEN_4; // @[ToAXI4.scala 105:45 ToAXI4.scala 110:14]
  assign io_out_req_bits_cmd = _T_20 & _T_21 ? {{1'd0}, _T_25} : _GEN_3; // @[ToAXI4.scala 105:45 ToAXI4.scala 107:13]
  assign io_out_req_bits_wmask = _T_20 & _T_21 ? io_in_wstrb : 8'h0; // @[ToAXI4.scala 105:45 ToAXI4.scala 111:15]
  assign io_out_req_bits_wdata = _T_20 & _T_21 ? io_in_wdata : 64'h0; // @[ToAXI4.scala 105:45 ToAXI4.scala 112:15]
  assign io_out_resp_ready = _T_2 | _T_7 & io_in_rready | _T_20 & io_in_bready; // @[ToAXI4.scala 128:73]
  always @(posedge clock) begin
    if (reset) begin // @[ToAXI4.scala 38:32]
      inflight_id_reg <= 18'h0; // @[ToAXI4.scala 38:32]
    end else if (_T_26) begin // @[ToAXI4.scala 120:21]
      inflight_id_reg <= 18'h0; // @[ToAXI4.scala 47:21]
    end else if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      if (_T_19) begin // @[ToAXI4.scala 100:24]
        inflight_id_reg <= io_in_awid; // @[ToAXI4.scala 42:21]
      end else begin
        inflight_id_reg <= _GEN_16;
      end
    end else begin
      inflight_id_reg <= _GEN_16;
    end
    if (reset) begin // @[ToAXI4.scala 40:30]
      inflight_type <= 2'h0; // @[ToAXI4.scala 40:30]
    end else if (_T_26) begin // @[ToAXI4.scala 120:21]
      inflight_type <= 2'h0; // @[ToAXI4.scala 46:19]
    end else if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      if (_T_19) begin // @[ToAXI4.scala 100:24]
        inflight_type <= 2'h2; // @[ToAXI4.scala 43:19]
      end else begin
        inflight_type <= _GEN_15;
      end
    end else begin
      inflight_type <= _GEN_15;
    end
    if (reset) begin // @[ToAXI4.scala 94:23]
      aw_reg_addr <= 32'h0; // @[ToAXI4.scala 94:23]
    end else if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      aw_reg_addr <= io_in_awaddr; // @[ToAXI4.scala 98:12]
    end
    if (reset) begin // @[ToAXI4.scala 94:23]
      aw_reg_len <= 8'h0; // @[ToAXI4.scala 94:23]
    end else if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      aw_reg_len <= io_in_awlen; // @[ToAXI4.scala 98:12]
    end
    if (reset) begin // @[ToAXI4.scala 94:23]
      aw_reg_size <= 3'h0; // @[ToAXI4.scala 94:23]
    end else if (_T_2 & io_in_awvalid & ~io_in_arvalid) begin // @[ToAXI4.scala 97:57]
      aw_reg_size <= io_in_awsize; // @[ToAXI4.scala 98:12]
    end
    if (reset) begin // @[ToAXI4.scala 95:25]
      bresp_en <= 1'h0; // @[ToAXI4.scala 95:25]
    end else if (_T_26) begin // @[ToAXI4.scala 120:21]
      bresp_en <= 1'h0; // @[ToAXI4.scala 121:14]
    end else if (_T_20 & _T_21) begin // @[ToAXI4.scala 105:45]
      bresp_en <= _GEN_27;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_57 & ~(_T_6 & _T_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:137 when (axi.ar.fire()) { assert(mem.req.fire() && !isInflight()); }\n"
            ); // @[ToAXI4.scala 137:32]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_57 & ~(_T_6 & _T_2 | reset)) begin
          $fatal; // @[ToAXI4.scala 137:32]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_19 & ~(_T_2 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:138 when (axi.aw.fire()) { assert(!isInflight()); }\n"); // @[ToAXI4.scala 138:32]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_19 & ~(_T_2 | reset)) begin
          $fatal; // @[ToAXI4.scala 138:32]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & ~(_T_6 & _T_20 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:139 when (axi.w.fire()) { assert(mem.req .fire() && isState(axi_write)); }\n"
            ); // @[ToAXI4.scala 139:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_21 & ~(_T_6 & _T_20 | reset)) begin
          $fatal; // @[ToAXI4.scala 139:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_26 & ~(_T_81 & _T_20 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:140 when (axi.b.fire()) { assert(mem.resp.fire() && isState(axi_write)); }\n"
            ); // @[ToAXI4.scala 140:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_26 & ~(_T_81 & _T_20 | reset)) begin
          $fatal; // @[ToAXI4.scala 140:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(_T_81 & _T_7 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at ToAXI4.scala:141 when (axi.r.fire()) { assert(mem.resp.fire() && isState(axi_read)); }\n"
            ); // @[ToAXI4.scala 141:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10 & ~(_T_81 & _T_7 | reset)) begin
          $fatal; // @[ToAXI4.scala 141:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inflight_id_reg = _RAND_0[17:0];
  _RAND_1 = {1{`RANDOM}};
  inflight_type = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  aw_reg_addr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  aw_reg_len = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  aw_reg_size = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  bresp_en = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_SimpleBusAddressMapper(
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
  assign io_in_req_ready = io_out_req_ready; // @[AddressMapper.scala 31:10]
  assign io_in_resp_valid = io_out_resp_valid; // @[AddressMapper.scala 31:10]
  assign io_in_resp_bits_cmd = io_out_resp_bits_cmd; // @[AddressMapper.scala 31:10]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[AddressMapper.scala 31:10]
  assign io_out_req_valid = io_in_req_valid; // @[AddressMapper.scala 31:10]
  assign io_out_req_bits_addr = io_in_req_bits_addr; // @[AddressMapper.scala 31:10]
  assign io_out_req_bits_size = io_in_req_bits_size; // @[AddressMapper.scala 31:10]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[AddressMapper.scala 31:10]
  assign io_out_req_bits_wmask = io_in_req_bits_wmask; // @[AddressMapper.scala 31:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[AddressMapper.scala 31:10]
  assign io_out_resp_ready = io_in_resp_ready; // @[AddressMapper.scala 31:10]
endmodule
module ysyx_210000_SimpleBusCrossbar1toN(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_0_req_ready,
  output        io_out_0_req_valid,
  output [31:0] io_out_0_req_bits_addr,
  output [2:0]  io_out_0_req_bits_size,
  output [3:0]  io_out_0_req_bits_cmd,
  output [7:0]  io_out_0_req_bits_wmask,
  output [63:0] io_out_0_req_bits_wdata,
  output        io_out_0_resp_ready,
  input         io_out_0_resp_valid,
  input  [3:0]  io_out_0_resp_bits_cmd,
  input  [63:0] io_out_0_resp_bits_rdata,
  input         io_out_1_req_ready,
  output        io_out_1_req_valid,
  output [31:0] io_out_1_req_bits_addr,
  output [3:0]  io_out_1_req_bits_cmd,
  output [7:0]  io_out_1_req_bits_wmask,
  output [63:0] io_out_1_req_bits_wdata,
  output        io_out_1_resp_ready,
  input         io_out_1_resp_valid,
  input  [63:0] io_out_1_resp_bits_rdata,
  input         io_out_2_req_ready,
  output        io_out_2_req_valid,
  output [31:0] io_out_2_req_bits_addr,
  output [3:0]  io_out_2_req_bits_cmd,
  output [7:0]  io_out_2_req_bits_wmask,
  output [63:0] io_out_2_req_bits_wdata,
  output        io_out_2_resp_ready,
  input         io_out_2_resp_valid,
  input  [63:0] io_out_2_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[Crossbar.scala 31:22]
  wire  outSelVec_0 = io_in_req_bits_addr >= 32'h10000000 & io_in_req_bits_addr < 32'h80000000; // @[Crossbar.scala 36:34]
  wire  outSelVec_1 = io_in_req_bits_addr >= 32'h2000000 & io_in_req_bits_addr < 32'h2010000; // @[Crossbar.scala 36:34]
  wire  outSelVec_2 = io_in_req_bits_addr >= 32'hc000000 & io_in_req_bits_addr < 32'h10000000; // @[Crossbar.scala 36:34]
  wire [1:0] _T_9 = outSelVec_1 ? 2'h1 : 2'h2; // @[Mux.scala 47:69]
  wire [1:0] outSelIdx = outSelVec_0 ? 2'h0 : _T_9; // @[Mux.scala 47:69]
  wire  _GEN_1 = 2'h1 == outSelIdx ? io_out_1_req_ready : io_out_0_req_ready; // @[Decoupled.scala 40:37 Decoupled.scala 40:37]
  wire  _GEN_2 = 2'h2 == outSelIdx ? io_out_2_req_ready : _GEN_1; // @[Decoupled.scala 40:37 Decoupled.scala 40:37]
  wire  _GEN_4 = 2'h1 == outSelIdx ? io_out_1_req_valid : io_out_0_req_valid; // @[Decoupled.scala 40:37 Decoupled.scala 40:37]
  wire  _GEN_5 = 2'h2 == outSelIdx ? io_out_2_req_valid : _GEN_4; // @[Decoupled.scala 40:37 Decoupled.scala 40:37]
  wire  _T_10 = _GEN_2 & _GEN_5; // @[Decoupled.scala 40:37]
  wire  _T_11 = state == 2'h0; // @[Crossbar.scala 39:97]
  wire  _T_12 = _T_10 & state == 2'h0; // @[Crossbar.scala 39:87]
  reg [1:0] outSelIdxResp; // @[Reg.scala 27:20]
  wire [2:0] _T_15 = {outSelVec_2,outSelVec_1,outSelVec_0}; // @[Crossbar.scala 41:54]
  wire  reqInvalidAddr = io_in_req_valid & ~(|_T_15); // @[Crossbar.scala 41:40]
  wire  _T_24 = io_in_req_valid & &_T_15; // @[Crossbar.scala 43:71]
  wire  _T_42 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_44 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _GEN_10 = 2'h1 == outSelIdxResp ? io_out_1_resp_ready : io_out_0_resp_ready; // @[Decoupled.scala 40:37 Decoupled.scala 40:37]
  wire  _GEN_11 = 2'h2 == outSelIdxResp ? io_out_2_resp_ready : _GEN_10; // @[Decoupled.scala 40:37 Decoupled.scala 40:37]
  wire  _GEN_13 = 2'h1 == outSelIdxResp ? io_out_1_resp_valid : io_out_0_resp_valid; // @[Decoupled.scala 40:37 Decoupled.scala 40:37]
  wire  _GEN_14 = 2'h2 == outSelIdxResp ? io_out_2_resp_valid : _GEN_13; // @[Decoupled.scala 40:37 Decoupled.scala 40:37]
  wire  _T_45 = _GEN_11 & _GEN_14; // @[Decoupled.scala 40:37]
  wire  _T_46 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_47 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_16 = _T_47 ? 2'h0 : state; // @[Crossbar.scala 64:43 Crossbar.scala 64:51 Crossbar.scala 31:22]
  wire [63:0] _GEN_21 = 2'h1 == outSelIdxResp ? io_out_1_resp_bits_rdata : io_out_0_resp_bits_rdata; // @[Crossbar.scala 68:19 Crossbar.scala 68:19]
  wire [3:0] _GEN_24 = 2'h1 == outSelIdxResp ? 4'h6 : io_out_0_resp_bits_cmd; // @[Crossbar.scala 68:19 Crossbar.scala 68:19]
  assign io_in_req_ready = _GEN_2 | reqInvalidAddr; // @[Crossbar.scala 71:39]
  assign io_in_resp_valid = _T_45 | state == 2'h2; // @[Crossbar.scala 67:46]
  assign io_in_resp_bits_cmd = 2'h2 == outSelIdxResp ? 4'h6 : _GEN_24; // @[Crossbar.scala 68:19 Crossbar.scala 68:19]
  assign io_in_resp_bits_rdata = 2'h2 == outSelIdxResp ? io_out_2_resp_bits_rdata : _GEN_21; // @[Crossbar.scala 68:19 Crossbar.scala 68:19]
  assign io_out_0_req_valid = outSelVec_0 & (io_in_req_valid & _T_11); // @[Crossbar.scala 54:22]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_0_resp_ready = 2'h0 == outSelIdxResp ? io_in_resp_ready : outSelVec_0; // @[Crossbar.scala 70:25 Crossbar.scala 70:25 Crossbar.scala 55:18]
  assign io_out_1_req_valid = outSelVec_1 & (io_in_req_valid & _T_11); // @[Crossbar.scala 54:22]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_1_resp_ready = 2'h1 == outSelIdxResp ? io_in_resp_ready : outSelVec_1; // @[Crossbar.scala 70:25 Crossbar.scala 70:25 Crossbar.scala 55:18]
  assign io_out_2_req_valid = outSelVec_2 & (io_in_req_valid & _T_11); // @[Crossbar.scala 54:22]
  assign io_out_2_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_2_resp_ready = 2'h2 == outSelIdxResp ? io_in_resp_ready : outSelVec_2; // @[Crossbar.scala 70:25 Crossbar.scala 70:25 Crossbar.scala 55:18]
  always @(posedge clock) begin
    if (reset) begin // @[Crossbar.scala 31:22]
      state <= 2'h0; // @[Crossbar.scala 31:22]
    end else if (_T_42) begin // @[Conditional.scala 40:58]
      if (reqInvalidAddr) begin // @[Crossbar.scala 61:29]
        state <= 2'h2; // @[Crossbar.scala 61:37]
      end else if (_T_10) begin // @[Crossbar.scala 60:32]
        state <= 2'h1; // @[Crossbar.scala 60:40]
      end
    end else if (_T_44) begin // @[Conditional.scala 39:67]
      if (_T_45) begin // @[Crossbar.scala 63:49]
        state <= 2'h0; // @[Crossbar.scala 63:57]
      end
    end else if (_T_46) begin // @[Conditional.scala 39:67]
      state <= _GEN_16;
    end
    if (reset) begin // @[Reg.scala 27:20]
      outSelIdxResp <= 2'h0; // @[Reg.scala 27:20]
    end else if (_T_12) begin // @[Reg.scala 28:19]
      if (outSelVec_0) begin // @[Mux.scala 47:69]
        outSelIdxResp <= 2'h0;
      end else if (outSelVec_1) begin // @[Mux.scala 47:69]
        outSelIdxResp <= 2'h1;
      end else begin
        outSelIdxResp <= 2'h2;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(~_T_24 | reset)) begin
          $fwrite(32'h80000002,
            "Assertion failed: address decode error, bad addr = 0x%x\n\n    at Crossbar.scala:49 assert(!(io.in.req.valid && outSelVec.asUInt.andR), \"address decode error, bad addr = 0x%%x\\n\", addr)\n"
            ,io_in_req_bits_addr); // @[Crossbar.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(~_T_24 | reset)) begin
          $fatal; // @[Crossbar.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelIdxResp = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_ReqBlocker(
  input         clock,
  input         reset,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [31:0] io_in_0_req_bits_addr,
  input  [2:0]  io_in_0_req_bits_size,
  input  [3:0]  io_in_0_req_bits_cmd,
  input  [7:0]  io_in_0_req_bits_wmask,
  input  [63:0] io_in_0_req_bits_wdata,
  input         io_in_0_resp_ready,
  output        io_in_0_resp_valid,
  output [3:0]  io_in_0_resp_bits_cmd,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [31:0] io_in_1_req_bits_addr,
  input  [2:0]  io_in_1_req_bits_size,
  input  [3:0]  io_in_1_req_bits_cmd,
  input  [7:0]  io_in_1_req_bits_wmask,
  input  [63:0] io_in_1_req_bits_wdata,
  input         io_in_1_resp_ready,
  output        io_in_1_resp_valid,
  output [3:0]  io_in_1_resp_bits_cmd,
  output [63:0] io_in_1_resp_bits_rdata,
  input         io_out_0_req_ready,
  output        io_out_0_req_valid,
  output [31:0] io_out_0_req_bits_addr,
  output [2:0]  io_out_0_req_bits_size,
  output [3:0]  io_out_0_req_bits_cmd,
  output [7:0]  io_out_0_req_bits_wmask,
  output [63:0] io_out_0_req_bits_wdata,
  output        io_out_0_resp_ready,
  input         io_out_0_resp_valid,
  input  [3:0]  io_out_0_resp_bits_cmd,
  input  [63:0] io_out_0_resp_bits_rdata,
  input         io_out_1_req_ready,
  output        io_out_1_req_valid,
  output [31:0] io_out_1_req_bits_addr,
  output [2:0]  io_out_1_req_bits_size,
  output [3:0]  io_out_1_req_bits_cmd,
  output [7:0]  io_out_1_req_bits_wmask,
  output [63:0] io_out_1_req_bits_wdata,
  output        io_out_1_resp_ready,
  input         io_out_1_resp_valid,
  input  [3:0]  io_out_1_resp_bits_cmd,
  input  [63:0] io_out_1_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Crossbar.scala 203:22]
  wire  chooseLo = io_in_0_req_valid & ~io_in_1_req_valid; // @[Crossbar.scala 206:37]
  wire  _T_1 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_2 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_3 = io_in_1_req_ready & io_in_1_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = io_in_0_req_ready & io_in_0_req_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_3 = _T_5 ? 3'h4 : state; // @[Crossbar.scala 217:34 Crossbar.scala 217:42 Crossbar.scala 203:22]
  wire  _T_6 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_7 = io_in_1_resp_ready & io_in_1_resp_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_4 = _T_7 ? 3'h0 : state; // @[Crossbar.scala 220:35 Crossbar.scala 220:43 Crossbar.scala 203:22]
  wire  _T_8 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_9 = io_in_0_resp_ready & io_in_0_resp_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_5 = _T_9 ? 3'h0 : state; // @[Crossbar.scala 223:35 Crossbar.scala 223:43 Crossbar.scala 203:22]
  wire [2:0] _GEN_6 = _T_8 ? _GEN_5 : state; // @[Conditional.scala 39:67 Crossbar.scala 203:22]
  wire [2:0] _GEN_7 = _T_6 ? _GEN_4 : _GEN_6; // @[Conditional.scala 39:67]
  wire  do_hi = state == 3'h1 | state == 3'h3; // @[Crossbar.scala 227:31]
  wire  do_lo = state == 3'h2 | state == 3'h4; // @[Crossbar.scala 228:31]
  assign io_in_0_req_ready = io_out_0_req_ready & do_lo; // @[Crossbar.scala 237:45]
  assign io_in_0_resp_valid = io_out_0_resp_valid; // @[Crossbar.scala 230:13]
  assign io_in_0_resp_bits_cmd = io_out_0_resp_bits_cmd; // @[Crossbar.scala 230:13]
  assign io_in_0_resp_bits_rdata = io_out_0_resp_bits_rdata; // @[Crossbar.scala 230:13]
  assign io_in_1_req_ready = io_out_1_req_ready & do_hi; // @[Crossbar.scala 234:45]
  assign io_in_1_resp_valid = io_out_1_resp_valid; // @[Crossbar.scala 231:13]
  assign io_in_1_resp_bits_cmd = io_out_1_resp_bits_cmd; // @[Crossbar.scala 231:13]
  assign io_in_1_resp_bits_rdata = io_out_1_resp_bits_rdata; // @[Crossbar.scala 231:13]
  assign io_out_0_req_valid = io_in_0_req_valid & do_lo; // @[Crossbar.scala 236:45]
  assign io_out_0_req_bits_addr = io_in_0_req_bits_addr; // @[Crossbar.scala 230:13]
  assign io_out_0_req_bits_size = io_in_0_req_bits_size; // @[Crossbar.scala 230:13]
  assign io_out_0_req_bits_cmd = io_in_0_req_bits_cmd; // @[Crossbar.scala 230:13]
  assign io_out_0_req_bits_wmask = io_in_0_req_bits_wmask; // @[Crossbar.scala 230:13]
  assign io_out_0_req_bits_wdata = io_in_0_req_bits_wdata; // @[Crossbar.scala 230:13]
  assign io_out_0_resp_ready = io_in_0_resp_ready; // @[Crossbar.scala 230:13]
  assign io_out_1_req_valid = io_in_1_req_valid & do_hi; // @[Crossbar.scala 233:45]
  assign io_out_1_req_bits_addr = io_in_1_req_bits_addr; // @[Crossbar.scala 231:13]
  assign io_out_1_req_bits_size = io_in_1_req_bits_size; // @[Crossbar.scala 231:13]
  assign io_out_1_req_bits_cmd = io_in_1_req_bits_cmd; // @[Crossbar.scala 231:13]
  assign io_out_1_req_bits_wmask = io_in_1_req_bits_wmask; // @[Crossbar.scala 231:13]
  assign io_out_1_req_bits_wdata = io_in_1_req_bits_wdata; // @[Crossbar.scala 231:13]
  assign io_out_1_resp_ready = io_in_1_resp_ready; // @[Crossbar.scala 231:13]
  always @(posedge clock) begin
    if (reset) begin // @[Crossbar.scala 203:22]
      state <= 3'h0; // @[Crossbar.scala 203:22]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      if (chooseLo) begin // @[Crossbar.scala 211:22]
        state <= 3'h2; // @[Crossbar.scala 211:30]
      end else if (io_in_1_req_valid) begin // @[Crossbar.scala 210:22]
        state <= 3'h1; // @[Crossbar.scala 210:30]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[Crossbar.scala 214:34]
        state <= 3'h3; // @[Crossbar.scala 214:42]
      end
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      state <= _GEN_3;
    end else begin
      state <= _GEN_7;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_SimpleBus2AXI4Converter(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_awready,
  output        io_out_awvalid,
  output [31:0] io_out_awaddr,
  output [3:0]  io_out_awid,
  output [7:0]  io_out_awlen,
  output [2:0]  io_out_awsize,
  output [1:0]  io_out_awburst,
  input         io_out_wready,
  output        io_out_wvalid,
  output [63:0] io_out_wdata,
  output [7:0]  io_out_wstrb,
  output        io_out_wlast,
  output        io_out_bready,
  input         io_out_bvalid,
  input         io_out_arready,
  output        io_out_arvalid,
  output [31:0] io_out_araddr,
  output [3:0]  io_out_arid,
  output [7:0]  io_out_arlen,
  output [2:0]  io_out_arsize,
  output [1:0]  io_out_arburst,
  output        io_out_rready,
  input         io_out_rvalid,
  input  [63:0] io_out_rdata,
  input         io_out_rlast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] _T_8 = io_in_req_bits_cmd[1] ? 3'h7 : 3'h0; // @[ToAXI4.scala 169:30]
  wire  _T_9 = io_in_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_10 = io_in_req_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire [2:0] _T_12 = io_out_rlast ? 3'h6 : 3'h0; // @[ToAXI4.scala 184:28]
  wire  _T_13 = io_out_awready & io_out_awvalid; // @[Decoupled.scala 40:37]
  reg  awAck; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_13 | awAck; // @[StopWatch.scala 30:20 StopWatch.scala 30:24 StopWatch.scala 24:20]
  wire  _T_17 = io_out_wready & io_out_wvalid; // @[Decoupled.scala 40:37]
  reg  wAck; // @[StopWatch.scala 24:20]
  wire  wSend = _T_13 & _T_17 & io_out_wlast | awAck & wAck; // @[ToAXI4.scala 189:53]
  wire  _T_15 = _T_17 & io_out_wlast; // @[ToAXI4.scala 188:41]
  wire  _GEN_2 = _T_15 | wAck; // @[StopWatch.scala 30:20 StopWatch.scala 30:24 StopWatch.scala 24:20]
  wire  _T_23 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg  wen; // @[Reg.scala 27:20]
  wire  _T_28 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_31 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  wire  _T_36 = ~wAck; // @[ToAXI4.scala 194:36]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_36 & io_out_wready : io_out_arready; // @[ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_bvalid : io_out_rvalid; // @[ToAXI4.scala 199:25]
  assign io_in_resp_bits_cmd = {{1'd0}, _T_12}; // @[ToAXI4.scala 184:28]
  assign io_in_resp_bits_rdata = io_out_rdata; // @[ToAXI4.scala 183:23]
  assign io_out_awvalid = _T_31 & ~awAck; // @[ToAXI4.scala 193:33]
  assign io_out_awaddr = io_out_araddr; // @[ToAXI4.scala 182:6]
  assign io_out_awid = io_out_arid; // @[ToAXI4.scala 182:6]
  assign io_out_awlen = io_out_arlen; // @[ToAXI4.scala 182:6]
  assign io_out_awsize = io_out_arsize; // @[ToAXI4.scala 182:6]
  assign io_out_awburst = io_out_arburst; // @[ToAXI4.scala 182:6]
  assign io_out_wvalid = _T_31 & ~wAck; // @[ToAXI4.scala 194:33]
  assign io_out_wdata = io_in_req_bits_wdata; // @[ToAXI4.scala 160:10]
  assign io_out_wstrb = io_in_req_bits_wmask; // @[ToAXI4.scala 161:10]
  assign io_out_wlast = _T_9 | _T_10; // @[ToAXI4.scala 177:54]
  assign io_out_bready = io_in_resp_ready; // @[ToAXI4.scala 198:16]
  assign io_out_arvalid = io_in_req_valid & _T_28; // @[SimpleBus.scala 104:29]
  assign io_out_araddr = io_in_req_bits_addr; // @[ToAXI4.scala 158:12]
  assign io_out_arid = 4'h0; // @[ToAXI4.scala 168:24]
  assign io_out_arlen = {{5'd0}, _T_8}; // @[ToAXI4.scala 169:30]
  assign io_out_arsize = io_in_req_bits_size; // @[ToAXI4.scala 170:24]
  assign io_out_arburst = 2'h2; // @[ToAXI4.scala 171:24]
  assign io_out_rready = io_in_resp_ready; // @[ToAXI4.scala 197:16]
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      awAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      awAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      wAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      wAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (reset) begin // @[Reg.scala 27:20]
      wen <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_23) begin // @[Reg.scala 28:19]
      wen <= io_in_req_bits_cmd[0]; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_AXI4CLINT(
  input         clock,
  input         reset,
  output        io__in_awready,
  input         io__in_awvalid,
  input  [31:0] io__in_awaddr,
  output        io__in_wready,
  input         io__in_wvalid,
  input  [63:0] io__in_wdata,
  input  [7:0]  io__in_wstrb,
  input         io__in_bready,
  output        io__in_bvalid,
  output        io__in_arready,
  input         io__in_arvalid,
  input  [31:0] io__in_araddr,
  input         io__in_rready,
  output        io__in_rvalid,
  output [63:0] io__in_rdata,
  output        io__extra_mtip,
  output        io__extra_msip,
  output        io_extra_mtip,
  output        io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] lo_lo_lo = io__in_wstrb[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lo_lo_hi = io__in_wstrb[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lo_hi_lo = io__in_wstrb[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lo_hi_hi = io__in_wstrb[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_lo_lo = io__in_wstrb[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_lo_hi = io__in_wstrb[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_hi_lo = io__in_wstrb[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_hi_hi = io__in_wstrb[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] fullMask = {hi_hi_hi,hi_hi_lo,hi_lo_hi,hi_lo_lo,lo_hi_hi,lo_hi_lo,lo_lo_hi,lo_lo_lo}; // @[Cat.scala 30:58]
  wire  _T_16 = io__in_arready & io__in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_17 = io__in_rready & io__in_rvalid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_17 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19 StopWatch.scala 26:23 StopWatch.scala 24:20]
  wire  _GEN_1 = _T_16 | _GEN_0; // @[StopWatch.scala 27:20 StopWatch.scala 27:24]
  reg  REG; // @[AXI4Slave.scala 73:17]
  wire  _T_28 = REG & (_T_16 | r_busy); // @[AXI4Slave.scala 74:35]
  reg  REG_1; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_17 ? 1'h0 : REG_1; // @[StopWatch.scala 26:19 StopWatch.scala 26:23 StopWatch.scala 24:20]
  wire  _GEN_3 = _T_28 | _GEN_2; // @[StopWatch.scala 27:20 StopWatch.scala 27:24]
  wire  _T_30 = io__in_awready & io__in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_31 = io__in_bready & io__in_bvalid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_31 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19 StopWatch.scala 26:23 StopWatch.scala 24:20]
  wire  _GEN_5 = _T_30 | _GEN_4; // @[StopWatch.scala 27:20 StopWatch.scala 27:24]
  wire  _T_34 = io__in_wready & io__in_wvalid; // @[Decoupled.scala 40:37]
  reg  REG_2; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_31 ? 1'h0 : REG_2; // @[StopWatch.scala 26:19 StopWatch.scala 26:23 StopWatch.scala 24:20]
  wire  _GEN_7 = _T_34 | _GEN_6; // @[StopWatch.scala 27:20 StopWatch.scala 27:24]
  reg [63:0] mtime; // @[AXI4CLINT.scala 32:22]
  reg [63:0] mtimecmp; // @[AXI4CLINT.scala 33:25]
  reg [63:0] msip; // @[AXI4CLINT.scala 34:21]
  reg [15:0] freq; // @[AXI4CLINT.scala 37:21]
  reg [15:0] inc; // @[AXI4CLINT.scala 38:20]
  reg [15:0] cnt; // @[AXI4CLINT.scala 40:20]
  wire [15:0] nextCnt = cnt + 16'h1; // @[AXI4CLINT.scala 41:21]
  wire  tick = nextCnt == freq; // @[AXI4CLINT.scala 43:23]
  wire [63:0] _GEN_14 = {{48'd0}, inc}; // @[AXI4CLINT.scala 44:32]
  wire [63:0] _T_41 = mtime + _GEN_14; // @[AXI4CLINT.scala 44:32]
  wire  _T_62 = 16'h0 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_63 = 16'h8000 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_64 = 16'hbff8 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_65 = 16'h8008 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_66 = 16'h4000 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_67 = _T_62 ? msip : 64'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_68 = _T_63 ? freq : 16'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_69 = _T_64 ? mtime : 64'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_70 = _T_65 ? inc : 16'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_71 = _T_66 ? mtimecmp : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_15 = {{48'd0}, _T_68}; // @[Mux.scala 27:72]
  wire [63:0] _T_72 = _T_67 | _GEN_15; // @[Mux.scala 27:72]
  wire [63:0] _T_73 = _T_72 | _T_69; // @[Mux.scala 27:72]
  wire [63:0] _GEN_16 = {{48'd0}, _T_70}; // @[Mux.scala 27:72]
  wire [63:0] _T_74 = _T_73 | _GEN_16; // @[Mux.scala 27:72]
  wire [63:0] _T_78 = io__in_wdata & fullMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_79 = ~fullMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_80 = msip & _T_79; // @[BitUtils.scala 32:36]
  wire [63:0] _T_81 = _T_78 | _T_80; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_17 = {{48'd0}, freq}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_86 = _GEN_17 & _T_79; // @[BitUtils.scala 32:36]
  wire [63:0] _T_87 = _T_78 | _T_86; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_10 = _T_34 & io__in_awaddr[15:0] == 16'h8000 ? _T_87 : {{48'd0}, freq}; // @[RegMap.scala 32:48 RegMap.scala 32:52 AXI4CLINT.scala 37:21]
  wire [63:0] _T_92 = mtime & _T_79; // @[BitUtils.scala 32:36]
  wire [63:0] _T_93 = _T_78 | _T_92; // @[BitUtils.scala 32:25]
  wire [63:0] _T_98 = _GEN_14 & _T_79; // @[BitUtils.scala 32:36]
  wire [63:0] _T_99 = _T_78 | _T_98; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_12 = _T_34 & io__in_awaddr[15:0] == 16'h8008 ? _T_99 : {{48'd0}, inc}; // @[RegMap.scala 32:48 RegMap.scala 32:52 AXI4CLINT.scala 38:20]
  wire [63:0] _T_104 = mtimecmp & _T_79; // @[BitUtils.scala 32:36]
  wire [63:0] _T_105 = _T_78 | _T_104; // @[BitUtils.scala 32:25]
  reg  REG_3; // @[AXI4CLINT.scala 64:31]
  reg  REG_4; // @[AXI4CLINT.scala 65:31]
  assign io__in_awready = ~w_busy; // @[AXI4Slave.scala 94:18]
  assign io__in_wready = io__in_awvalid | w_busy; // @[AXI4Slave.scala 95:30]
  assign io__in_bvalid = REG_2; // @[AXI4Slave.scala 97:14]
  assign io__in_arready = io__in_rready | ~r_busy; // @[AXI4Slave.scala 71:29]
  assign io__in_rvalid = REG_1; // @[AXI4Slave.scala 74:14]
  assign io__in_rdata = _T_74 | _T_71; // @[Mux.scala 27:72]
  assign io__extra_mtip = REG_3; // @[AXI4CLINT.scala 64:21]
  assign io__extra_msip = REG_4; // @[AXI4CLINT.scala 65:21]
  assign io_extra_mtip = io__extra_mtip;
  assign io_extra_msip = io__extra_msip;
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[AXI4Slave.scala 73:17]
      REG <= 1'h0; // @[AXI4Slave.scala 73:17]
    end else begin
      REG <= _T_16; // @[AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_1 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_1 <= _GEN_3;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_2 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_2 <= _GEN_7;
    end
    if (reset) begin // @[AXI4CLINT.scala 32:22]
      mtime <= 64'h0; // @[AXI4CLINT.scala 32:22]
    end else if (_T_34 & io__in_awaddr[15:0] == 16'hbff8) begin // @[RegMap.scala 32:48]
      mtime <= _T_93; // @[RegMap.scala 32:52]
    end else if (tick) begin // @[AXI4CLINT.scala 44:15]
      mtime <= _T_41; // @[AXI4CLINT.scala 44:23]
    end
    if (reset) begin // @[AXI4CLINT.scala 33:25]
      mtimecmp <= 64'h0; // @[AXI4CLINT.scala 33:25]
    end else if (_T_34 & io__in_awaddr[15:0] == 16'h4000) begin // @[RegMap.scala 32:48]
      mtimecmp <= _T_105; // @[RegMap.scala 32:52]
    end
    if (reset) begin // @[AXI4CLINT.scala 34:21]
      msip <= 64'h0; // @[AXI4CLINT.scala 34:21]
    end else if (_T_34 & io__in_awaddr[15:0] == 16'h0) begin // @[RegMap.scala 32:48]
      msip <= _T_81; // @[RegMap.scala 32:52]
    end
    if (reset) begin // @[AXI4CLINT.scala 37:21]
      freq <= 16'h28; // @[AXI4CLINT.scala 37:21]
    end else begin
      freq <= _GEN_10[15:0];
    end
    if (reset) begin // @[AXI4CLINT.scala 38:20]
      inc <= 16'h1; // @[AXI4CLINT.scala 38:20]
    end else begin
      inc <= _GEN_12[15:0];
    end
    if (reset) begin // @[AXI4CLINT.scala 40:20]
      cnt <= 16'h0; // @[AXI4CLINT.scala 40:20]
    end else if (nextCnt < freq) begin // @[AXI4CLINT.scala 42:13]
      cnt <= nextCnt;
    end else begin
      cnt <= 16'h0;
    end
    if (reset) begin // @[AXI4CLINT.scala 64:31]
      REG_3 <= 1'h0; // @[AXI4CLINT.scala 64:31]
    end else begin
      REG_3 <= mtime >= mtimecmp; // @[AXI4CLINT.scala 64:31]
    end
    if (reset) begin // @[AXI4CLINT.scala 65:31]
      REG_4 <= 1'h0; // @[AXI4CLINT.scala 65:31]
    end else begin
      REG_4 <= msip != 64'h0; // @[AXI4CLINT.scala 65:31]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_2 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  mtime = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mtimecmp = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  msip = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  freq = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  inc = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  cnt = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  REG_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  REG_4 = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_SimpleBus2AXI4Converter_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_awready,
  output        io_out_awvalid,
  output [31:0] io_out_awaddr,
  input         io_out_wready,
  output        io_out_wvalid,
  output [63:0] io_out_wdata,
  output [7:0]  io_out_wstrb,
  output        io_out_bready,
  input         io_out_bvalid,
  input         io_out_arready,
  output        io_out_arvalid,
  output [31:0] io_out_araddr,
  output        io_out_rready,
  input         io_out_rvalid,
  input  [63:0] io_out_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  toAXI4Lite = ~(io_in_req_valid & io_in_req_bits_cmd[1]); // @[ToAXI4.scala 151:20]
  wire  _T_8 = io_out_awready & io_out_awvalid; // @[Decoupled.scala 40:37]
  reg  awAck; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_8 | awAck; // @[StopWatch.scala 30:20 StopWatch.scala 30:24 StopWatch.scala 24:20]
  wire  _T_12 = io_out_wready & io_out_wvalid; // @[Decoupled.scala 40:37]
  reg  wAck; // @[StopWatch.scala 24:20]
  wire  wSend = _T_8 & _T_12 | awAck & wAck; // @[ToAXI4.scala 189:53]
  wire  _GEN_2 = _T_12 | wAck; // @[StopWatch.scala 30:20 StopWatch.scala 30:24 StopWatch.scala 24:20]
  wire  _T_18 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg  wen; // @[Reg.scala 27:20]
  wire  _T_23 = ~io_in_req_bits_cmd[0] & ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:26]
  wire  _T_26 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  wire  _T_31 = ~wAck; // @[ToAXI4.scala 194:36]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_31 & io_out_wready : io_out_arready; // @[ToAXI4.scala 195:24]
  assign io_in_resp_valid = wen ? io_out_bvalid : io_out_rvalid; // @[ToAXI4.scala 199:25]
  assign io_in_resp_bits_rdata = io_out_rdata; // @[ToAXI4.scala 183:23]
  assign io_out_awvalid = _T_26 & ~awAck; // @[ToAXI4.scala 193:33]
  assign io_out_awaddr = io_out_araddr; // @[ToAXI4.scala 182:6]
  assign io_out_wvalid = _T_26 & ~wAck; // @[ToAXI4.scala 194:33]
  assign io_out_wdata = io_in_req_bits_wdata; // @[ToAXI4.scala 160:10]
  assign io_out_wstrb = io_in_req_bits_wmask; // @[ToAXI4.scala 161:10]
  assign io_out_bready = io_in_resp_ready; // @[ToAXI4.scala 198:16]
  assign io_out_arvalid = io_in_req_valid & _T_23; // @[SimpleBus.scala 104:29]
  assign io_out_araddr = io_in_req_bits_addr; // @[ToAXI4.scala 158:12]
  assign io_out_rready = io_in_resp_ready; // @[ToAXI4.scala 197:16]
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      awAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      awAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      wAck <= 1'h0; // @[StopWatch.scala 24:20]
    end else if (wSend) begin // @[StopWatch.scala 31:19]
      wAck <= 1'h0; // @[StopWatch.scala 31:23]
    end else begin
      wAck <= _GEN_2;
    end
    if (reset) begin // @[Reg.scala 27:20]
      wen <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_18) begin // @[Reg.scala 28:19]
      wen <= io_in_req_bits_cmd[0]; // @[Reg.scala 28:23]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~(toAXI4Lite | reset)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (~(toAXI4Lite | reset)) begin
          $fatal; // @[ToAXI4.scala 153:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_AXI4PLIC(
  input         clock,
  input         reset,
  output        io__in_awready,
  input         io__in_awvalid,
  input  [31:0] io__in_awaddr,
  output        io__in_wready,
  input         io__in_wvalid,
  input  [63:0] io__in_wdata,
  input  [7:0]  io__in_wstrb,
  input         io__in_bready,
  output        io__in_bvalid,
  output        io__in_arready,
  input         io__in_arvalid,
  input  [31:0] io__in_araddr,
  input         io__in_rready,
  output        io__in_rvalid,
  output [63:0] io__in_rdata,
  input         io__extra_intrVec,
  output        io__extra_meip_0,
  output        io_extra_meip_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  _T_16 = io__in_arready & io__in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_17 = io__in_rready & io__in_rvalid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_17 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19 StopWatch.scala 26:23 StopWatch.scala 24:20]
  wire  _GEN_1 = _T_16 | _GEN_0; // @[StopWatch.scala 27:20 StopWatch.scala 27:24]
  reg  REG; // @[AXI4Slave.scala 73:17]
  wire  _T_28 = REG & (_T_16 | r_busy); // @[AXI4Slave.scala 74:35]
  reg  REG_1; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_17 ? 1'h0 : REG_1; // @[StopWatch.scala 26:19 StopWatch.scala 26:23 StopWatch.scala 24:20]
  wire  _GEN_3 = _T_28 | _GEN_2; // @[StopWatch.scala 27:20 StopWatch.scala 27:24]
  wire  _T_30 = io__in_awready & io__in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_31 = io__in_bready & io__in_bvalid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_31 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19 StopWatch.scala 26:23 StopWatch.scala 24:20]
  wire  _GEN_5 = _T_30 | _GEN_4; // @[StopWatch.scala 27:20 StopWatch.scala 27:24]
  wire  _T_34 = io__in_wready & io__in_wvalid; // @[Decoupled.scala 40:37]
  reg  REG_2; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_31 ? 1'h0 : REG_2; // @[StopWatch.scala 26:19 StopWatch.scala 26:23 StopWatch.scala 24:20]
  wire  _GEN_7 = _T_34 | _GEN_6; // @[StopWatch.scala 27:20 StopWatch.scala 27:24]
  reg [31:0] priority_0; // @[AXI4PLIC.scala 37:43]
  reg  pending_0_1; // @[AXI4PLIC.scala 43:46]
  wire [31:0] _T_37 = {16'h0,8'h0,4'h0,2'h0,pending_0_1,1'h0}; // @[Cat.scala 30:58]
  reg [31:0] enable_0_0; // @[AXI4PLIC.scala 48:64]
  reg [31:0] threshold_0; // @[AXI4PLIC.scala 53:44]
  reg  inHandle_1; // @[AXI4PLIC.scala 58:25]
  reg [31:0] claimCompletion_0; // @[AXI4PLIC.scala 64:50]
  wire  _GEN_11 = _T_17 & io__in_araddr[25:0] == 26'h200004 ? claimCompletion_0[0] | inHandle_1 : inHandle_1; // @[AXI4PLIC.scala 68:59 AXI4PLIC.scala 58:25]
  wire  _GEN_12 = io__extra_intrVec | pending_0_1; // @[AXI4PLIC.scala 75:17 AXI4PLIC.scala 75:45 AXI4PLIC.scala 43:46]
  wire [31:0] _T_44 = _T_37 & enable_0_0; // @[AXI4PLIC.scala 81:31]
  wire [4:0] _T_78 = _T_44[30] ? 5'h1e : 5'h1f; // @[Mux.scala 47:69]
  wire [4:0] _T_79 = _T_44[29] ? 5'h1d : _T_78; // @[Mux.scala 47:69]
  wire [4:0] _T_80 = _T_44[28] ? 5'h1c : _T_79; // @[Mux.scala 47:69]
  wire [4:0] _T_81 = _T_44[27] ? 5'h1b : _T_80; // @[Mux.scala 47:69]
  wire [4:0] _T_82 = _T_44[26] ? 5'h1a : _T_81; // @[Mux.scala 47:69]
  wire [4:0] _T_83 = _T_44[25] ? 5'h19 : _T_82; // @[Mux.scala 47:69]
  wire [4:0] _T_84 = _T_44[24] ? 5'h18 : _T_83; // @[Mux.scala 47:69]
  wire [4:0] _T_85 = _T_44[23] ? 5'h17 : _T_84; // @[Mux.scala 47:69]
  wire [4:0] _T_86 = _T_44[22] ? 5'h16 : _T_85; // @[Mux.scala 47:69]
  wire [4:0] _T_87 = _T_44[21] ? 5'h15 : _T_86; // @[Mux.scala 47:69]
  wire [4:0] _T_88 = _T_44[20] ? 5'h14 : _T_87; // @[Mux.scala 47:69]
  wire [4:0] _T_89 = _T_44[19] ? 5'h13 : _T_88; // @[Mux.scala 47:69]
  wire [4:0] _T_90 = _T_44[18] ? 5'h12 : _T_89; // @[Mux.scala 47:69]
  wire [4:0] _T_91 = _T_44[17] ? 5'h11 : _T_90; // @[Mux.scala 47:69]
  wire [4:0] _T_92 = _T_44[16] ? 5'h10 : _T_91; // @[Mux.scala 47:69]
  wire [4:0] _T_93 = _T_44[15] ? 5'hf : _T_92; // @[Mux.scala 47:69]
  wire [4:0] _T_94 = _T_44[14] ? 5'he : _T_93; // @[Mux.scala 47:69]
  wire [4:0] _T_95 = _T_44[13] ? 5'hd : _T_94; // @[Mux.scala 47:69]
  wire [4:0] _T_96 = _T_44[12] ? 5'hc : _T_95; // @[Mux.scala 47:69]
  wire [4:0] _T_97 = _T_44[11] ? 5'hb : _T_96; // @[Mux.scala 47:69]
  wire [4:0] _T_98 = _T_44[10] ? 5'ha : _T_97; // @[Mux.scala 47:69]
  wire [4:0] _T_99 = _T_44[9] ? 5'h9 : _T_98; // @[Mux.scala 47:69]
  wire [4:0] _T_100 = _T_44[8] ? 5'h8 : _T_99; // @[Mux.scala 47:69]
  wire [4:0] _T_101 = _T_44[7] ? 5'h7 : _T_100; // @[Mux.scala 47:69]
  wire [4:0] _T_102 = _T_44[6] ? 5'h6 : _T_101; // @[Mux.scala 47:69]
  wire [4:0] _T_103 = _T_44[5] ? 5'h5 : _T_102; // @[Mux.scala 47:69]
  wire [4:0] _T_104 = _T_44[4] ? 5'h4 : _T_103; // @[Mux.scala 47:69]
  wire [4:0] _T_105 = _T_44[3] ? 5'h3 : _T_104; // @[Mux.scala 47:69]
  wire [4:0] _T_106 = _T_44[2] ? 5'h2 : _T_105; // @[Mux.scala 47:69]
  wire [4:0] _T_107 = _T_44[1] ? 5'h1 : _T_106; // @[Mux.scala 47:69]
  wire [4:0] _T_108 = _T_44[0] ? 5'h0 : _T_107; // @[Mux.scala 47:69]
  wire [4:0] _T_109 = _T_44 == 32'h0 ? 5'h0 : _T_108; // @[AXI4PLIC.scala 82:13]
  wire [7:0] _T_114 = io__in_wstrb >> io__in_awaddr[2:0]; // @[AXI4PLIC.scala 89:78]
  wire [7:0] lo_lo_lo_3 = _T_114[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lo_lo_hi_3 = _T_114[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lo_hi_lo_3 = _T_114[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lo_hi_hi_3 = _T_114[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_lo_lo_3 = _T_114[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_lo_hi_3 = _T_114[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_hi_lo_3 = _T_114[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] hi_hi_hi_3 = _T_114[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_131 = {hi_hi_hi_3,hi_hi_lo_3,hi_lo_hi_3,hi_lo_lo_3,lo_hi_hi_3,lo_hi_lo_3,lo_lo_hi_3,lo_lo_lo_3}; // @[Cat.scala 30:58]
  wire  _T_132 = 26'h1000 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_133 = 26'h2000 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_134 = 26'h200004 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_135 = 26'h4 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_136 = 26'h200000 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire [31:0] _T_137 = _T_132 ? _T_37 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_138 = _T_133 ? enable_0_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_139 = _T_134 ? claimCompletion_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_140 = _T_135 ? priority_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_141 = _T_136 ? threshold_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_142 = _T_137 | _T_138; // @[Mux.scala 27:72]
  wire [31:0] _T_143 = _T_142 | _T_139; // @[Mux.scala 27:72]
  wire [31:0] _T_144 = _T_143 | _T_140; // @[Mux.scala 27:72]
  wire [31:0] rdata = _T_144 | _T_141; // @[Mux.scala 27:72]
  wire [63:0] _T_148 = io__in_wdata & _T_131; // @[BitUtils.scala 32:13]
  wire [63:0] _T_149 = ~_T_131; // @[BitUtils.scala 32:38]
  wire [63:0] _GEN_23 = {{32'd0}, enable_0_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_150 = _GEN_23 & _T_149; // @[BitUtils.scala 32:36]
  wire [63:0] _T_151 = _T_148 | _T_150; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_14 = _T_34 & io__in_awaddr[25:0] == 26'h2000 ? _T_151 : {{32'd0}, enable_0_0}; // @[RegMap.scala 32:48 RegMap.scala 32:52 AXI4PLIC.scala 48:64]
  wire [63:0] _GEN_24 = {{32'd0}, claimCompletion_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_156 = _GEN_24 & _T_149; // @[BitUtils.scala 32:36]
  wire [63:0] _T_157 = _T_148 | _T_156; // @[BitUtils.scala 32:25]
  wire [4:0] _GEN_19 = _T_34 & io__in_awaddr[25:0] == 26'h200004 ? 5'h0 : _T_109; // @[RegMap.scala 32:48 RegMap.scala 32:52 AXI4PLIC.scala 82:7]
  wire [63:0] _GEN_25 = {{32'd0}, priority_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_164 = _GEN_25 & _T_149; // @[BitUtils.scala 32:36]
  wire [63:0] _T_165 = _T_148 | _T_164; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_20 = _T_34 & io__in_awaddr[25:0] == 26'h4 ? _T_165 : {{32'd0}, priority_0}; // @[RegMap.scala 32:48 RegMap.scala 32:52 AXI4PLIC.scala 37:43]
  wire [63:0] _GEN_26 = {{32'd0}, threshold_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_170 = _GEN_26 & _T_149; // @[BitUtils.scala 32:36]
  wire [63:0] _T_171 = _T_148 | _T_170; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_21 = _T_34 & io__in_awaddr[25:0] == 26'h200000 ? _T_171 : {{32'd0}, threshold_0}; // @[RegMap.scala 32:48 RegMap.scala 32:52 AXI4PLIC.scala 53:44]
  wire [4:0] _GEN_27 = reset ? 5'h0 : _GEN_19; // @[AXI4PLIC.scala 64:50 AXI4PLIC.scala 64:50]
  assign io__in_awready = ~w_busy; // @[AXI4Slave.scala 94:18]
  assign io__in_wready = io__in_awvalid | w_busy; // @[AXI4Slave.scala 95:30]
  assign io__in_bvalid = REG_2; // @[AXI4Slave.scala 97:14]
  assign io__in_arready = io__in_rready | ~r_busy; // @[AXI4Slave.scala 71:29]
  assign io__in_rvalid = REG_1; // @[AXI4Slave.scala 74:14]
  assign io__in_rdata = {rdata,rdata}; // @[Cat.scala 30:58]
  assign io__extra_meip_0 = claimCompletion_0 != 32'h0; // @[AXI4PLIC.scala 93:87]
  assign io_extra_meip_0 = io__extra_meip_0;
  always @(posedge clock) begin
    if (reset) begin // @[StopWatch.scala 24:20]
      r_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin // @[AXI4Slave.scala 73:17]
      REG <= 1'h0; // @[AXI4Slave.scala 73:17]
    end else begin
      REG <= _T_16; // @[AXI4Slave.scala 73:17]
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_1 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_1 <= _GEN_3;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      w_busy <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin // @[StopWatch.scala 24:20]
      REG_2 <= 1'h0; // @[StopWatch.scala 24:20]
    end else begin
      REG_2 <= _GEN_7;
    end
    if (reset) begin // @[AXI4PLIC.scala 37:43]
      priority_0 <= 32'h0; // @[AXI4PLIC.scala 37:43]
    end else begin
      priority_0 <= _GEN_20[31:0];
    end
    if (reset) begin // @[AXI4PLIC.scala 43:46]
      pending_0_1 <= 1'h0; // @[AXI4PLIC.scala 43:46]
    end else if (inHandle_1) begin // @[AXI4PLIC.scala 76:25]
      pending_0_1 <= 1'h0; // @[AXI4PLIC.scala 76:53]
    end else begin
      pending_0_1 <= _GEN_12;
    end
    if (reset) begin // @[AXI4PLIC.scala 48:64]
      enable_0_0 <= 32'h0; // @[AXI4PLIC.scala 48:64]
    end else begin
      enable_0_0 <= _GEN_14[31:0];
    end
    if (reset) begin // @[AXI4PLIC.scala 53:44]
      threshold_0 <= 32'h0; // @[AXI4PLIC.scala 53:44]
    end else begin
      threshold_0 <= _GEN_21[31:0];
    end
    if (reset) begin // @[AXI4PLIC.scala 58:25]
      inHandle_1 <= 1'h0; // @[AXI4PLIC.scala 58:25]
    end else if (_T_34 & io__in_awaddr[25:0] == 26'h200004) begin // @[RegMap.scala 32:48]
      if (_T_157[0]) begin // @[AXI4PLIC.scala 60:27]
        inHandle_1 <= 1'h0; // @[AXI4PLIC.scala 60:27]
      end else begin
        inHandle_1 <= _GEN_11;
      end
    end else begin
      inHandle_1 <= _GEN_11;
    end
    claimCompletion_0 <= {{27'd0}, _GEN_27}; // @[AXI4PLIC.scala 64:50 AXI4PLIC.scala 64:50]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  priority_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  pending_0_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  enable_0_0 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  threshold_0 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  inHandle_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  claimCompletion_0 = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000(
  input         clock,
  input         reset,
  input         io_master_awready,
  output        io_master_awvalid,
  output [31:0] io_master_awaddr,
  output [3:0]  io_master_awid,
  output [7:0]  io_master_awlen,
  output [2:0]  io_master_awsize,
  output [1:0]  io_master_awburst,
  input         io_master_wready,
  output        io_master_wvalid,
  output [63:0] io_master_wdata,
  output [7:0]  io_master_wstrb,
  output        io_master_wlast,
  output        io_master_bready,
  input         io_master_bvalid,
  input  [1:0]  io_master_bresp,
  input  [3:0]  io_master_bid,
  input         io_master_arready,
  output        io_master_arvalid,
  output [31:0] io_master_araddr,
  output [3:0]  io_master_arid,
  output [7:0]  io_master_arlen,
  output [2:0]  io_master_arsize,
  output [1:0]  io_master_arburst,
  output        io_master_rready,
  input         io_master_rvalid,
  input  [1:0]  io_master_rresp,
  input  [63:0] io_master_rdata,
  input         io_master_rlast,
  input  [3:0]  io_master_rid,
  output        io_slave_awready,
  input         io_slave_awvalid,
  input  [31:0] io_slave_awaddr,
  input  [3:0]  io_slave_awid,
  input  [7:0]  io_slave_awlen,
  input  [2:0]  io_slave_awsize,
  input  [1:0]  io_slave_awburst,
  output        io_slave_wready,
  input         io_slave_wvalid,
  input  [63:0] io_slave_wdata,
  input  [7:0]  io_slave_wstrb,
  input         io_slave_wlast,
  input         io_slave_bready,
  output        io_slave_bvalid,
  output [1:0]  io_slave_bresp,
  output [3:0]  io_slave_bid,
  output        io_slave_arready,
  input         io_slave_arvalid,
  input  [31:0] io_slave_araddr,
  input  [3:0]  io_slave_arid,
  input  [7:0]  io_slave_arlen,
  input  [2:0]  io_slave_arsize,
  input  [1:0]  io_slave_arburst,
  input         io_slave_rready,
  output        io_slave_rvalid,
  output [1:0]  io_slave_rresp,
  output [63:0] io_slave_rdata,
  output        io_slave_rlast,
  output [3:0]  io_slave_rid,
  input         io_interrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  nutcore_clock; // @[NutShell.scala 54:23]
  wire  nutcore_reset; // @[NutShell.scala 54:23]
  wire  nutcore_io_imem_mem_req_ready; // @[NutShell.scala 54:23]
  wire  nutcore_io_imem_mem_req_valid; // @[NutShell.scala 54:23]
  wire [31:0] nutcore_io_imem_mem_req_bits_addr; // @[NutShell.scala 54:23]
  wire [3:0] nutcore_io_imem_mem_req_bits_cmd; // @[NutShell.scala 54:23]
  wire [63:0] nutcore_io_imem_mem_req_bits_wdata; // @[NutShell.scala 54:23]
  wire  nutcore_io_imem_mem_resp_valid; // @[NutShell.scala 54:23]
  wire [3:0] nutcore_io_imem_mem_resp_bits_cmd; // @[NutShell.scala 54:23]
  wire [63:0] nutcore_io_imem_mem_resp_bits_rdata; // @[NutShell.scala 54:23]
  wire  nutcore_io_dmem_mem_req_ready; // @[NutShell.scala 54:23]
  wire  nutcore_io_dmem_mem_req_valid; // @[NutShell.scala 54:23]
  wire [31:0] nutcore_io_dmem_mem_req_bits_addr; // @[NutShell.scala 54:23]
  wire [3:0] nutcore_io_dmem_mem_req_bits_cmd; // @[NutShell.scala 54:23]
  wire [63:0] nutcore_io_dmem_mem_req_bits_wdata; // @[NutShell.scala 54:23]
  wire  nutcore_io_dmem_mem_resp_valid; // @[NutShell.scala 54:23]
  wire [3:0] nutcore_io_dmem_mem_resp_bits_cmd; // @[NutShell.scala 54:23]
  wire [63:0] nutcore_io_dmem_mem_resp_bits_rdata; // @[NutShell.scala 54:23]
  wire  nutcore_io_dmem_coh_req_ready; // @[NutShell.scala 54:23]
  wire  nutcore_io_dmem_coh_req_valid; // @[NutShell.scala 54:23]
  wire [31:0] nutcore_io_dmem_coh_req_bits_addr; // @[NutShell.scala 54:23]
  wire [63:0] nutcore_io_dmem_coh_req_bits_wdata; // @[NutShell.scala 54:23]
  wire  nutcore_io_dmem_coh_resp_valid; // @[NutShell.scala 54:23]
  wire [3:0] nutcore_io_dmem_coh_resp_bits_cmd; // @[NutShell.scala 54:23]
  wire [63:0] nutcore_io_dmem_coh_resp_bits_rdata; // @[NutShell.scala 54:23]
  wire  nutcore_io_mmio_req_ready; // @[NutShell.scala 54:23]
  wire  nutcore_io_mmio_req_valid; // @[NutShell.scala 54:23]
  wire [31:0] nutcore_io_mmio_req_bits_addr; // @[NutShell.scala 54:23]
  wire [2:0] nutcore_io_mmio_req_bits_size; // @[NutShell.scala 54:23]
  wire [3:0] nutcore_io_mmio_req_bits_cmd; // @[NutShell.scala 54:23]
  wire [7:0] nutcore_io_mmio_req_bits_wmask; // @[NutShell.scala 54:23]
  wire [63:0] nutcore_io_mmio_req_bits_wdata; // @[NutShell.scala 54:23]
  wire  nutcore_io_mmio_resp_ready; // @[NutShell.scala 54:23]
  wire  nutcore_io_mmio_resp_valid; // @[NutShell.scala 54:23]
  wire [3:0] nutcore_io_mmio_resp_bits_cmd; // @[NutShell.scala 54:23]
  wire [63:0] nutcore_io_mmio_resp_bits_rdata; // @[NutShell.scala 54:23]
  wire  nutcore_io_frontend_req_ready; // @[NutShell.scala 54:23]
  wire  nutcore_io_frontend_req_valid; // @[NutShell.scala 54:23]
  wire [31:0] nutcore_io_frontend_req_bits_addr; // @[NutShell.scala 54:23]
  wire [2:0] nutcore_io_frontend_req_bits_size; // @[NutShell.scala 54:23]
  wire [3:0] nutcore_io_frontend_req_bits_cmd; // @[NutShell.scala 54:23]
  wire [7:0] nutcore_io_frontend_req_bits_wmask; // @[NutShell.scala 54:23]
  wire [63:0] nutcore_io_frontend_req_bits_wdata; // @[NutShell.scala 54:23]
  wire  nutcore_io_frontend_resp_ready; // @[NutShell.scala 54:23]
  wire  nutcore_io_frontend_resp_valid; // @[NutShell.scala 54:23]
  wire [3:0] nutcore_io_frontend_resp_bits_cmd; // @[NutShell.scala 54:23]
  wire [63:0] nutcore_io_frontend_resp_bits_rdata; // @[NutShell.scala 54:23]
  wire  nutcore_io_extra_mtip; // @[NutShell.scala 54:23]
  wire  nutcore_io_extra_meip_0; // @[NutShell.scala 54:23]
  wire  nutcore_io_extra_msip; // @[NutShell.scala 54:23]
  wire  cohMg_clock; // @[NutShell.scala 55:21]
  wire  cohMg_reset; // @[NutShell.scala 55:21]
  wire  cohMg_io_in_req_ready; // @[NutShell.scala 55:21]
  wire  cohMg_io_in_req_valid; // @[NutShell.scala 55:21]
  wire [31:0] cohMg_io_in_req_bits_addr; // @[NutShell.scala 55:21]
  wire [3:0] cohMg_io_in_req_bits_cmd; // @[NutShell.scala 55:21]
  wire [63:0] cohMg_io_in_req_bits_wdata; // @[NutShell.scala 55:21]
  wire  cohMg_io_in_resp_valid; // @[NutShell.scala 55:21]
  wire [3:0] cohMg_io_in_resp_bits_cmd; // @[NutShell.scala 55:21]
  wire [63:0] cohMg_io_in_resp_bits_rdata; // @[NutShell.scala 55:21]
  wire  cohMg_io_out_mem_req_ready; // @[NutShell.scala 55:21]
  wire  cohMg_io_out_mem_req_valid; // @[NutShell.scala 55:21]
  wire [31:0] cohMg_io_out_mem_req_bits_addr; // @[NutShell.scala 55:21]
  wire [2:0] cohMg_io_out_mem_req_bits_size; // @[NutShell.scala 55:21]
  wire [3:0] cohMg_io_out_mem_req_bits_cmd; // @[NutShell.scala 55:21]
  wire [7:0] cohMg_io_out_mem_req_bits_wmask; // @[NutShell.scala 55:21]
  wire [63:0] cohMg_io_out_mem_req_bits_wdata; // @[NutShell.scala 55:21]
  wire  cohMg_io_out_mem_resp_ready; // @[NutShell.scala 55:21]
  wire  cohMg_io_out_mem_resp_valid; // @[NutShell.scala 55:21]
  wire [3:0] cohMg_io_out_mem_resp_bits_cmd; // @[NutShell.scala 55:21]
  wire [63:0] cohMg_io_out_mem_resp_bits_rdata; // @[NutShell.scala 55:21]
  wire  cohMg_io_out_coh_req_ready; // @[NutShell.scala 55:21]
  wire  cohMg_io_out_coh_req_valid; // @[NutShell.scala 55:21]
  wire [31:0] cohMg_io_out_coh_req_bits_addr; // @[NutShell.scala 55:21]
  wire [63:0] cohMg_io_out_coh_req_bits_wdata; // @[NutShell.scala 55:21]
  wire  cohMg_io_out_coh_resp_ready; // @[NutShell.scala 55:21]
  wire  cohMg_io_out_coh_resp_valid; // @[NutShell.scala 55:21]
  wire [3:0] cohMg_io_out_coh_resp_bits_cmd; // @[NutShell.scala 55:21]
  wire [63:0] cohMg_io_out_coh_resp_bits_rdata; // @[NutShell.scala 55:21]
  wire  xbar_clock; // @[NutShell.scala 56:20]
  wire  xbar_reset; // @[NutShell.scala 56:20]
  wire  xbar_io_in_0_req_ready; // @[NutShell.scala 56:20]
  wire  xbar_io_in_0_req_valid; // @[NutShell.scala 56:20]
  wire [31:0] xbar_io_in_0_req_bits_addr; // @[NutShell.scala 56:20]
  wire [2:0] xbar_io_in_0_req_bits_size; // @[NutShell.scala 56:20]
  wire [3:0] xbar_io_in_0_req_bits_cmd; // @[NutShell.scala 56:20]
  wire [7:0] xbar_io_in_0_req_bits_wmask; // @[NutShell.scala 56:20]
  wire [63:0] xbar_io_in_0_req_bits_wdata; // @[NutShell.scala 56:20]
  wire  xbar_io_in_0_resp_ready; // @[NutShell.scala 56:20]
  wire  xbar_io_in_0_resp_valid; // @[NutShell.scala 56:20]
  wire [3:0] xbar_io_in_0_resp_bits_cmd; // @[NutShell.scala 56:20]
  wire [63:0] xbar_io_in_0_resp_bits_rdata; // @[NutShell.scala 56:20]
  wire  xbar_io_in_1_req_ready; // @[NutShell.scala 56:20]
  wire  xbar_io_in_1_req_valid; // @[NutShell.scala 56:20]
  wire [31:0] xbar_io_in_1_req_bits_addr; // @[NutShell.scala 56:20]
  wire [2:0] xbar_io_in_1_req_bits_size; // @[NutShell.scala 56:20]
  wire [3:0] xbar_io_in_1_req_bits_cmd; // @[NutShell.scala 56:20]
  wire [7:0] xbar_io_in_1_req_bits_wmask; // @[NutShell.scala 56:20]
  wire [63:0] xbar_io_in_1_req_bits_wdata; // @[NutShell.scala 56:20]
  wire  xbar_io_in_1_resp_ready; // @[NutShell.scala 56:20]
  wire  xbar_io_in_1_resp_valid; // @[NutShell.scala 56:20]
  wire [3:0] xbar_io_in_1_resp_bits_cmd; // @[NutShell.scala 56:20]
  wire [63:0] xbar_io_in_1_resp_bits_rdata; // @[NutShell.scala 56:20]
  wire  xbar_io_out_req_ready; // @[NutShell.scala 56:20]
  wire  xbar_io_out_req_valid; // @[NutShell.scala 56:20]
  wire [31:0] xbar_io_out_req_bits_addr; // @[NutShell.scala 56:20]
  wire [2:0] xbar_io_out_req_bits_size; // @[NutShell.scala 56:20]
  wire [3:0] xbar_io_out_req_bits_cmd; // @[NutShell.scala 56:20]
  wire [7:0] xbar_io_out_req_bits_wmask; // @[NutShell.scala 56:20]
  wire [63:0] xbar_io_out_req_bits_wdata; // @[NutShell.scala 56:20]
  wire  xbar_io_out_resp_ready; // @[NutShell.scala 56:20]
  wire  xbar_io_out_resp_valid; // @[NutShell.scala 56:20]
  wire [3:0] xbar_io_out_resp_bits_cmd; // @[NutShell.scala 56:20]
  wire [63:0] xbar_io_out_resp_bits_rdata; // @[NutShell.scala 56:20]
  wire  axi2sb_clock; // @[NutShell.scala 62:22]
  wire  axi2sb_reset; // @[NutShell.scala 62:22]
  wire  axi2sb_io_in_awready; // @[NutShell.scala 62:22]
  wire  axi2sb_io_in_awvalid; // @[NutShell.scala 62:22]
  wire [31:0] axi2sb_io_in_awaddr; // @[NutShell.scala 62:22]
  wire [17:0] axi2sb_io_in_awid; // @[NutShell.scala 62:22]
  wire [7:0] axi2sb_io_in_awlen; // @[NutShell.scala 62:22]
  wire [2:0] axi2sb_io_in_awsize; // @[NutShell.scala 62:22]
  wire  axi2sb_io_in_wready; // @[NutShell.scala 62:22]
  wire  axi2sb_io_in_wvalid; // @[NutShell.scala 62:22]
  wire [63:0] axi2sb_io_in_wdata; // @[NutShell.scala 62:22]
  wire [7:0] axi2sb_io_in_wstrb; // @[NutShell.scala 62:22]
  wire  axi2sb_io_in_wlast; // @[NutShell.scala 62:22]
  wire  axi2sb_io_in_bready; // @[NutShell.scala 62:22]
  wire  axi2sb_io_in_bvalid; // @[NutShell.scala 62:22]
  wire  axi2sb_io_in_arready; // @[NutShell.scala 62:22]
  wire  axi2sb_io_in_arvalid; // @[NutShell.scala 62:22]
  wire [31:0] axi2sb_io_in_araddr; // @[NutShell.scala 62:22]
  wire [17:0] axi2sb_io_in_arid; // @[NutShell.scala 62:22]
  wire [7:0] axi2sb_io_in_arlen; // @[NutShell.scala 62:22]
  wire [2:0] axi2sb_io_in_arsize; // @[NutShell.scala 62:22]
  wire  axi2sb_io_in_rready; // @[NutShell.scala 62:22]
  wire  axi2sb_io_in_rvalid; // @[NutShell.scala 62:22]
  wire [63:0] axi2sb_io_in_rdata; // @[NutShell.scala 62:22]
  wire  axi2sb_io_in_rlast; // @[NutShell.scala 62:22]
  wire [17:0] axi2sb_io_in_rid; // @[NutShell.scala 62:22]
  wire  axi2sb_io_out_req_ready; // @[NutShell.scala 62:22]
  wire  axi2sb_io_out_req_valid; // @[NutShell.scala 62:22]
  wire [31:0] axi2sb_io_out_req_bits_addr; // @[NutShell.scala 62:22]
  wire [2:0] axi2sb_io_out_req_bits_size; // @[NutShell.scala 62:22]
  wire [3:0] axi2sb_io_out_req_bits_cmd; // @[NutShell.scala 62:22]
  wire [7:0] axi2sb_io_out_req_bits_wmask; // @[NutShell.scala 62:22]
  wire [63:0] axi2sb_io_out_req_bits_wdata; // @[NutShell.scala 62:22]
  wire  axi2sb_io_out_resp_ready; // @[NutShell.scala 62:22]
  wire  axi2sb_io_out_resp_valid; // @[NutShell.scala 62:22]
  wire [3:0] axi2sb_io_out_resp_bits_cmd; // @[NutShell.scala 62:22]
  wire [63:0] axi2sb_io_out_resp_bits_rdata; // @[NutShell.scala 62:22]
  wire  memAddrMap_io_in_req_ready; // @[NutShell.scala 94:26]
  wire  memAddrMap_io_in_req_valid; // @[NutShell.scala 94:26]
  wire [31:0] memAddrMap_io_in_req_bits_addr; // @[NutShell.scala 94:26]
  wire [2:0] memAddrMap_io_in_req_bits_size; // @[NutShell.scala 94:26]
  wire [3:0] memAddrMap_io_in_req_bits_cmd; // @[NutShell.scala 94:26]
  wire [7:0] memAddrMap_io_in_req_bits_wmask; // @[NutShell.scala 94:26]
  wire [63:0] memAddrMap_io_in_req_bits_wdata; // @[NutShell.scala 94:26]
  wire  memAddrMap_io_in_resp_ready; // @[NutShell.scala 94:26]
  wire  memAddrMap_io_in_resp_valid; // @[NutShell.scala 94:26]
  wire [3:0] memAddrMap_io_in_resp_bits_cmd; // @[NutShell.scala 94:26]
  wire [63:0] memAddrMap_io_in_resp_bits_rdata; // @[NutShell.scala 94:26]
  wire  memAddrMap_io_out_req_ready; // @[NutShell.scala 94:26]
  wire  memAddrMap_io_out_req_valid; // @[NutShell.scala 94:26]
  wire [31:0] memAddrMap_io_out_req_bits_addr; // @[NutShell.scala 94:26]
  wire [2:0] memAddrMap_io_out_req_bits_size; // @[NutShell.scala 94:26]
  wire [3:0] memAddrMap_io_out_req_bits_cmd; // @[NutShell.scala 94:26]
  wire [7:0] memAddrMap_io_out_req_bits_wmask; // @[NutShell.scala 94:26]
  wire [63:0] memAddrMap_io_out_req_bits_wdata; // @[NutShell.scala 94:26]
  wire  memAddrMap_io_out_resp_ready; // @[NutShell.scala 94:26]
  wire  memAddrMap_io_out_resp_valid; // @[NutShell.scala 94:26]
  wire [3:0] memAddrMap_io_out_resp_bits_cmd; // @[NutShell.scala 94:26]
  wire [63:0] memAddrMap_io_out_resp_bits_rdata; // @[NutShell.scala 94:26]
  wire  mmioXbar_clock; // @[NutShell.scala 106:24]
  wire  mmioXbar_reset; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_in_req_bits_addr; // @[NutShell.scala 106:24]
  wire [2:0] mmioXbar_io_in_req_bits_size; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_in_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_resp_valid; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_resp_bits_cmd; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_0_req_bits_addr; // @[NutShell.scala 106:24]
  wire [2:0] mmioXbar_io_out_0_req_bits_size; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_0_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_0_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_valid; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_0_resp_bits_cmd; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_1_req_bits_addr; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_1_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_1_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_valid; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_2_req_bits_addr; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_2_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_2_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_valid; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  ReqBlocker_clock; // @[NutShell.scala 120:25]
  wire  ReqBlocker_reset; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_in_0_req_ready; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_in_0_req_valid; // @[NutShell.scala 120:25]
  wire [31:0] ReqBlocker_io_in_0_req_bits_addr; // @[NutShell.scala 120:25]
  wire [2:0] ReqBlocker_io_in_0_req_bits_size; // @[NutShell.scala 120:25]
  wire [3:0] ReqBlocker_io_in_0_req_bits_cmd; // @[NutShell.scala 120:25]
  wire [7:0] ReqBlocker_io_in_0_req_bits_wmask; // @[NutShell.scala 120:25]
  wire [63:0] ReqBlocker_io_in_0_req_bits_wdata; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_in_0_resp_ready; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_in_0_resp_valid; // @[NutShell.scala 120:25]
  wire [3:0] ReqBlocker_io_in_0_resp_bits_cmd; // @[NutShell.scala 120:25]
  wire [63:0] ReqBlocker_io_in_0_resp_bits_rdata; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_in_1_req_ready; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_in_1_req_valid; // @[NutShell.scala 120:25]
  wire [31:0] ReqBlocker_io_in_1_req_bits_addr; // @[NutShell.scala 120:25]
  wire [2:0] ReqBlocker_io_in_1_req_bits_size; // @[NutShell.scala 120:25]
  wire [3:0] ReqBlocker_io_in_1_req_bits_cmd; // @[NutShell.scala 120:25]
  wire [7:0] ReqBlocker_io_in_1_req_bits_wmask; // @[NutShell.scala 120:25]
  wire [63:0] ReqBlocker_io_in_1_req_bits_wdata; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_in_1_resp_ready; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_in_1_resp_valid; // @[NutShell.scala 120:25]
  wire [3:0] ReqBlocker_io_in_1_resp_bits_cmd; // @[NutShell.scala 120:25]
  wire [63:0] ReqBlocker_io_in_1_resp_bits_rdata; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_out_0_req_ready; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_out_0_req_valid; // @[NutShell.scala 120:25]
  wire [31:0] ReqBlocker_io_out_0_req_bits_addr; // @[NutShell.scala 120:25]
  wire [2:0] ReqBlocker_io_out_0_req_bits_size; // @[NutShell.scala 120:25]
  wire [3:0] ReqBlocker_io_out_0_req_bits_cmd; // @[NutShell.scala 120:25]
  wire [7:0] ReqBlocker_io_out_0_req_bits_wmask; // @[NutShell.scala 120:25]
  wire [63:0] ReqBlocker_io_out_0_req_bits_wdata; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_out_0_resp_ready; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_out_0_resp_valid; // @[NutShell.scala 120:25]
  wire [3:0] ReqBlocker_io_out_0_resp_bits_cmd; // @[NutShell.scala 120:25]
  wire [63:0] ReqBlocker_io_out_0_resp_bits_rdata; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_out_1_req_ready; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_out_1_req_valid; // @[NutShell.scala 120:25]
  wire [31:0] ReqBlocker_io_out_1_req_bits_addr; // @[NutShell.scala 120:25]
  wire [2:0] ReqBlocker_io_out_1_req_bits_size; // @[NutShell.scala 120:25]
  wire [3:0] ReqBlocker_io_out_1_req_bits_cmd; // @[NutShell.scala 120:25]
  wire [7:0] ReqBlocker_io_out_1_req_bits_wmask; // @[NutShell.scala 120:25]
  wire [63:0] ReqBlocker_io_out_1_req_bits_wdata; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_out_1_resp_ready; // @[NutShell.scala 120:25]
  wire  ReqBlocker_io_out_1_resp_valid; // @[NutShell.scala 120:25]
  wire [3:0] ReqBlocker_io_out_1_resp_bits_cmd; // @[NutShell.scala 120:25]
  wire [63:0] ReqBlocker_io_out_1_resp_bits_rdata; // @[NutShell.scala 120:25]
  wire  SimpleBusCrossbarNto1_clock; // @[NutShell.scala 121:28]
  wire  SimpleBusCrossbarNto1_reset; // @[NutShell.scala 121:28]
  wire  SimpleBusCrossbarNto1_io_in_0_req_ready; // @[NutShell.scala 121:28]
  wire  SimpleBusCrossbarNto1_io_in_0_req_valid; // @[NutShell.scala 121:28]
  wire [31:0] SimpleBusCrossbarNto1_io_in_0_req_bits_addr; // @[NutShell.scala 121:28]
  wire [2:0] SimpleBusCrossbarNto1_io_in_0_req_bits_size; // @[NutShell.scala 121:28]
  wire [3:0] SimpleBusCrossbarNto1_io_in_0_req_bits_cmd; // @[NutShell.scala 121:28]
  wire [7:0] SimpleBusCrossbarNto1_io_in_0_req_bits_wmask; // @[NutShell.scala 121:28]
  wire [63:0] SimpleBusCrossbarNto1_io_in_0_req_bits_wdata; // @[NutShell.scala 121:28]
  wire  SimpleBusCrossbarNto1_io_in_0_resp_ready; // @[NutShell.scala 121:28]
  wire  SimpleBusCrossbarNto1_io_in_0_resp_valid; // @[NutShell.scala 121:28]
  wire [3:0] SimpleBusCrossbarNto1_io_in_0_resp_bits_cmd; // @[NutShell.scala 121:28]
  wire [63:0] SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata; // @[NutShell.scala 121:28]
  wire  SimpleBusCrossbarNto1_io_in_1_req_ready; // @[NutShell.scala 121:28]
  wire  SimpleBusCrossbarNto1_io_in_1_req_valid; // @[NutShell.scala 121:28]
  wire [31:0] SimpleBusCrossbarNto1_io_in_1_req_bits_addr; // @[NutShell.scala 121:28]
  wire [2:0] SimpleBusCrossbarNto1_io_in_1_req_bits_size; // @[NutShell.scala 121:28]
  wire [3:0] SimpleBusCrossbarNto1_io_in_1_req_bits_cmd; // @[NutShell.scala 121:28]
  wire [7:0] SimpleBusCrossbarNto1_io_in_1_req_bits_wmask; // @[NutShell.scala 121:28]
  wire [63:0] SimpleBusCrossbarNto1_io_in_1_req_bits_wdata; // @[NutShell.scala 121:28]
  wire  SimpleBusCrossbarNto1_io_in_1_resp_ready; // @[NutShell.scala 121:28]
  wire  SimpleBusCrossbarNto1_io_in_1_resp_valid; // @[NutShell.scala 121:28]
  wire [3:0] SimpleBusCrossbarNto1_io_in_1_resp_bits_cmd; // @[NutShell.scala 121:28]
  wire [63:0] SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata; // @[NutShell.scala 121:28]
  wire  SimpleBusCrossbarNto1_io_out_req_ready; // @[NutShell.scala 121:28]
  wire  SimpleBusCrossbarNto1_io_out_req_valid; // @[NutShell.scala 121:28]
  wire [31:0] SimpleBusCrossbarNto1_io_out_req_bits_addr; // @[NutShell.scala 121:28]
  wire [2:0] SimpleBusCrossbarNto1_io_out_req_bits_size; // @[NutShell.scala 121:28]
  wire [3:0] SimpleBusCrossbarNto1_io_out_req_bits_cmd; // @[NutShell.scala 121:28]
  wire [7:0] SimpleBusCrossbarNto1_io_out_req_bits_wmask; // @[NutShell.scala 121:28]
  wire [63:0] SimpleBusCrossbarNto1_io_out_req_bits_wdata; // @[NutShell.scala 121:28]
  wire  SimpleBusCrossbarNto1_io_out_resp_ready; // @[NutShell.scala 121:28]
  wire  SimpleBusCrossbarNto1_io_out_resp_valid; // @[NutShell.scala 121:28]
  wire [3:0] SimpleBusCrossbarNto1_io_out_resp_bits_cmd; // @[NutShell.scala 121:28]
  wire [63:0] SimpleBusCrossbarNto1_io_out_resp_bits_rdata; // @[NutShell.scala 121:28]
  wire  SimpleBus2AXI4Converter_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_in_req_bits_size; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_in_resp_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_out_awid; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_io_out_awlen; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_awsize; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_io_out_awburst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_io_out_wstrb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_wlast; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_bready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_out_arid; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_io_out_arlen; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_arsize; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_io_out_arburst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_rready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_out_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_rlast; // @[ToAXI4.scala 204:24]
  wire  clint_clock; // @[NutShell.scala 129:21]
  wire  clint_reset; // @[NutShell.scala 129:21]
  wire  clint_io__in_awready; // @[NutShell.scala 129:21]
  wire  clint_io__in_awvalid; // @[NutShell.scala 129:21]
  wire [31:0] clint_io__in_awaddr; // @[NutShell.scala 129:21]
  wire  clint_io__in_wready; // @[NutShell.scala 129:21]
  wire  clint_io__in_wvalid; // @[NutShell.scala 129:21]
  wire [63:0] clint_io__in_wdata; // @[NutShell.scala 129:21]
  wire [7:0] clint_io__in_wstrb; // @[NutShell.scala 129:21]
  wire  clint_io__in_bready; // @[NutShell.scala 129:21]
  wire  clint_io__in_bvalid; // @[NutShell.scala 129:21]
  wire  clint_io__in_arready; // @[NutShell.scala 129:21]
  wire  clint_io__in_arvalid; // @[NutShell.scala 129:21]
  wire [31:0] clint_io__in_araddr; // @[NutShell.scala 129:21]
  wire  clint_io__in_rready; // @[NutShell.scala 129:21]
  wire  clint_io__in_rvalid; // @[NutShell.scala 129:21]
  wire [63:0] clint_io__in_rdata; // @[NutShell.scala 129:21]
  wire  clint_io__extra_mtip; // @[NutShell.scala 129:21]
  wire  clint_io__extra_msip; // @[NutShell.scala 129:21]
  wire  clint_io_extra_mtip; // @[NutShell.scala 129:21]
  wire  clint_io_extra_msip; // @[NutShell.scala 129:21]
  wire  SimpleBus2AXI4Converter_1_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_out_wstrb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_bready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_rready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_out_rdata; // @[ToAXI4.scala 204:24]
  wire  plic_clock; // @[NutShell.scala 136:20]
  wire  plic_reset; // @[NutShell.scala 136:20]
  wire  plic_io__in_awready; // @[NutShell.scala 136:20]
  wire  plic_io__in_awvalid; // @[NutShell.scala 136:20]
  wire [31:0] plic_io__in_awaddr; // @[NutShell.scala 136:20]
  wire  plic_io__in_wready; // @[NutShell.scala 136:20]
  wire  plic_io__in_wvalid; // @[NutShell.scala 136:20]
  wire [63:0] plic_io__in_wdata; // @[NutShell.scala 136:20]
  wire [7:0] plic_io__in_wstrb; // @[NutShell.scala 136:20]
  wire  plic_io__in_bready; // @[NutShell.scala 136:20]
  wire  plic_io__in_bvalid; // @[NutShell.scala 136:20]
  wire  plic_io__in_arready; // @[NutShell.scala 136:20]
  wire  plic_io__in_arvalid; // @[NutShell.scala 136:20]
  wire [31:0] plic_io__in_araddr; // @[NutShell.scala 136:20]
  wire  plic_io__in_rready; // @[NutShell.scala 136:20]
  wire  plic_io__in_rvalid; // @[NutShell.scala 136:20]
  wire [63:0] plic_io__in_rdata; // @[NutShell.scala 136:20]
  wire  plic_io__extra_intrVec; // @[NutShell.scala 136:20]
  wire  plic_io__extra_meip_0; // @[NutShell.scala 136:20]
  wire  plic_io_extra_meip_0; // @[NutShell.scala 136:20]
  wire  SimpleBus2AXI4Converter_2_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_2_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_2_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_2_io_out_wstrb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_bready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_rready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_out_rdata; // @[ToAXI4.scala 204:24]
  reg  REG; // @[NutShell.scala 138:47]
  reg  REG_1; // @[NutShell.scala 138:39]
  ysyx_210000_NutCore nutcore ( // @[NutShell.scala 54:23]
    .clock(nutcore_clock),
    .reset(nutcore_reset),
    .io_imem_mem_req_ready(nutcore_io_imem_mem_req_ready),
    .io_imem_mem_req_valid(nutcore_io_imem_mem_req_valid),
    .io_imem_mem_req_bits_addr(nutcore_io_imem_mem_req_bits_addr),
    .io_imem_mem_req_bits_cmd(nutcore_io_imem_mem_req_bits_cmd),
    .io_imem_mem_req_bits_wdata(nutcore_io_imem_mem_req_bits_wdata),
    .io_imem_mem_resp_valid(nutcore_io_imem_mem_resp_valid),
    .io_imem_mem_resp_bits_cmd(nutcore_io_imem_mem_resp_bits_cmd),
    .io_imem_mem_resp_bits_rdata(nutcore_io_imem_mem_resp_bits_rdata),
    .io_dmem_mem_req_ready(nutcore_io_dmem_mem_req_ready),
    .io_dmem_mem_req_valid(nutcore_io_dmem_mem_req_valid),
    .io_dmem_mem_req_bits_addr(nutcore_io_dmem_mem_req_bits_addr),
    .io_dmem_mem_req_bits_cmd(nutcore_io_dmem_mem_req_bits_cmd),
    .io_dmem_mem_req_bits_wdata(nutcore_io_dmem_mem_req_bits_wdata),
    .io_dmem_mem_resp_valid(nutcore_io_dmem_mem_resp_valid),
    .io_dmem_mem_resp_bits_cmd(nutcore_io_dmem_mem_resp_bits_cmd),
    .io_dmem_mem_resp_bits_rdata(nutcore_io_dmem_mem_resp_bits_rdata),
    .io_dmem_coh_req_ready(nutcore_io_dmem_coh_req_ready),
    .io_dmem_coh_req_valid(nutcore_io_dmem_coh_req_valid),
    .io_dmem_coh_req_bits_addr(nutcore_io_dmem_coh_req_bits_addr),
    .io_dmem_coh_req_bits_wdata(nutcore_io_dmem_coh_req_bits_wdata),
    .io_dmem_coh_resp_valid(nutcore_io_dmem_coh_resp_valid),
    .io_dmem_coh_resp_bits_cmd(nutcore_io_dmem_coh_resp_bits_cmd),
    .io_dmem_coh_resp_bits_rdata(nutcore_io_dmem_coh_resp_bits_rdata),
    .io_mmio_req_ready(nutcore_io_mmio_req_ready),
    .io_mmio_req_valid(nutcore_io_mmio_req_valid),
    .io_mmio_req_bits_addr(nutcore_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(nutcore_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(nutcore_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(nutcore_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(nutcore_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(nutcore_io_mmio_resp_ready),
    .io_mmio_resp_valid(nutcore_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(nutcore_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(nutcore_io_mmio_resp_bits_rdata),
    .io_frontend_req_ready(nutcore_io_frontend_req_ready),
    .io_frontend_req_valid(nutcore_io_frontend_req_valid),
    .io_frontend_req_bits_addr(nutcore_io_frontend_req_bits_addr),
    .io_frontend_req_bits_size(nutcore_io_frontend_req_bits_size),
    .io_frontend_req_bits_cmd(nutcore_io_frontend_req_bits_cmd),
    .io_frontend_req_bits_wmask(nutcore_io_frontend_req_bits_wmask),
    .io_frontend_req_bits_wdata(nutcore_io_frontend_req_bits_wdata),
    .io_frontend_resp_ready(nutcore_io_frontend_resp_ready),
    .io_frontend_resp_valid(nutcore_io_frontend_resp_valid),
    .io_frontend_resp_bits_cmd(nutcore_io_frontend_resp_bits_cmd),
    .io_frontend_resp_bits_rdata(nutcore_io_frontend_resp_bits_rdata),
    .io_extra_mtip(nutcore_io_extra_mtip),
    .io_extra_meip_0(nutcore_io_extra_meip_0),
    .io_extra_msip(nutcore_io_extra_msip)
  );
  ysyx_210000_CoherenceManager cohMg ( // @[NutShell.scala 55:21]
    .clock(cohMg_clock),
    .reset(cohMg_reset),
    .io_in_req_ready(cohMg_io_in_req_ready),
    .io_in_req_valid(cohMg_io_in_req_valid),
    .io_in_req_bits_addr(cohMg_io_in_req_bits_addr),
    .io_in_req_bits_cmd(cohMg_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(cohMg_io_in_req_bits_wdata),
    .io_in_resp_valid(cohMg_io_in_resp_valid),
    .io_in_resp_bits_cmd(cohMg_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(cohMg_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(cohMg_io_out_mem_req_ready),
    .io_out_mem_req_valid(cohMg_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(cohMg_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_size(cohMg_io_out_mem_req_bits_size),
    .io_out_mem_req_bits_cmd(cohMg_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wmask(cohMg_io_out_mem_req_bits_wmask),
    .io_out_mem_req_bits_wdata(cohMg_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_ready(cohMg_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(cohMg_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(cohMg_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(cohMg_io_out_mem_resp_bits_rdata),
    .io_out_coh_req_ready(cohMg_io_out_coh_req_ready),
    .io_out_coh_req_valid(cohMg_io_out_coh_req_valid),
    .io_out_coh_req_bits_addr(cohMg_io_out_coh_req_bits_addr),
    .io_out_coh_req_bits_wdata(cohMg_io_out_coh_req_bits_wdata),
    .io_out_coh_resp_ready(cohMg_io_out_coh_resp_ready),
    .io_out_coh_resp_valid(cohMg_io_out_coh_resp_valid),
    .io_out_coh_resp_bits_cmd(cohMg_io_out_coh_resp_bits_cmd),
    .io_out_coh_resp_bits_rdata(cohMg_io_out_coh_resp_bits_rdata)
  );
  ysyx_210000_SimpleBusCrossbarNto1 xbar ( // @[NutShell.scala 56:20]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_in_0_req_ready(xbar_io_in_0_req_ready),
    .io_in_0_req_valid(xbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(xbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(xbar_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(xbar_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(xbar_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(xbar_io_in_0_req_bits_wdata),
    .io_in_0_resp_ready(xbar_io_in_0_resp_ready),
    .io_in_0_resp_valid(xbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(xbar_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(xbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(xbar_io_in_1_req_ready),
    .io_in_1_req_valid(xbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(xbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(xbar_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(xbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(xbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(xbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_ready(xbar_io_in_1_resp_ready),
    .io_in_1_resp_valid(xbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(xbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(xbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(xbar_io_out_req_ready),
    .io_out_req_valid(xbar_io_out_req_valid),
    .io_out_req_bits_addr(xbar_io_out_req_bits_addr),
    .io_out_req_bits_size(xbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(xbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(xbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(xbar_io_out_req_bits_wdata),
    .io_out_resp_ready(xbar_io_out_resp_ready),
    .io_out_resp_valid(xbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(xbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(xbar_io_out_resp_bits_rdata)
  );
  ysyx_210000_AXI42SimpleBusConverter axi2sb ( // @[NutShell.scala 62:22]
    .clock(axi2sb_clock),
    .reset(axi2sb_reset),
    .io_in_awready(axi2sb_io_in_awready),
    .io_in_awvalid(axi2sb_io_in_awvalid),
    .io_in_awaddr(axi2sb_io_in_awaddr),
    .io_in_awid(axi2sb_io_in_awid),
    .io_in_awlen(axi2sb_io_in_awlen),
    .io_in_awsize(axi2sb_io_in_awsize),
    .io_in_wready(axi2sb_io_in_wready),
    .io_in_wvalid(axi2sb_io_in_wvalid),
    .io_in_wdata(axi2sb_io_in_wdata),
    .io_in_wstrb(axi2sb_io_in_wstrb),
    .io_in_wlast(axi2sb_io_in_wlast),
    .io_in_bready(axi2sb_io_in_bready),
    .io_in_bvalid(axi2sb_io_in_bvalid),
    .io_in_arready(axi2sb_io_in_arready),
    .io_in_arvalid(axi2sb_io_in_arvalid),
    .io_in_araddr(axi2sb_io_in_araddr),
    .io_in_arid(axi2sb_io_in_arid),
    .io_in_arlen(axi2sb_io_in_arlen),
    .io_in_arsize(axi2sb_io_in_arsize),
    .io_in_rready(axi2sb_io_in_rready),
    .io_in_rvalid(axi2sb_io_in_rvalid),
    .io_in_rdata(axi2sb_io_in_rdata),
    .io_in_rlast(axi2sb_io_in_rlast),
    .io_in_rid(axi2sb_io_in_rid),
    .io_out_req_ready(axi2sb_io_out_req_ready),
    .io_out_req_valid(axi2sb_io_out_req_valid),
    .io_out_req_bits_addr(axi2sb_io_out_req_bits_addr),
    .io_out_req_bits_size(axi2sb_io_out_req_bits_size),
    .io_out_req_bits_cmd(axi2sb_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(axi2sb_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(axi2sb_io_out_req_bits_wdata),
    .io_out_resp_ready(axi2sb_io_out_resp_ready),
    .io_out_resp_valid(axi2sb_io_out_resp_valid),
    .io_out_resp_bits_cmd(axi2sb_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(axi2sb_io_out_resp_bits_rdata)
  );
  ysyx_210000_SimpleBusAddressMapper memAddrMap ( // @[NutShell.scala 94:26]
    .io_in_req_ready(memAddrMap_io_in_req_ready),
    .io_in_req_valid(memAddrMap_io_in_req_valid),
    .io_in_req_bits_addr(memAddrMap_io_in_req_bits_addr),
    .io_in_req_bits_size(memAddrMap_io_in_req_bits_size),
    .io_in_req_bits_cmd(memAddrMap_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(memAddrMap_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(memAddrMap_io_in_req_bits_wdata),
    .io_in_resp_ready(memAddrMap_io_in_resp_ready),
    .io_in_resp_valid(memAddrMap_io_in_resp_valid),
    .io_in_resp_bits_cmd(memAddrMap_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(memAddrMap_io_in_resp_bits_rdata),
    .io_out_req_ready(memAddrMap_io_out_req_ready),
    .io_out_req_valid(memAddrMap_io_out_req_valid),
    .io_out_req_bits_addr(memAddrMap_io_out_req_bits_addr),
    .io_out_req_bits_size(memAddrMap_io_out_req_bits_size),
    .io_out_req_bits_cmd(memAddrMap_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(memAddrMap_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(memAddrMap_io_out_req_bits_wdata),
    .io_out_resp_ready(memAddrMap_io_out_resp_ready),
    .io_out_resp_valid(memAddrMap_io_out_resp_valid),
    .io_out_resp_bits_cmd(memAddrMap_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(memAddrMap_io_out_resp_bits_rdata)
  );
  ysyx_210000_SimpleBusCrossbar1toN mmioXbar ( // @[NutShell.scala 106:24]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_req_ready(mmioXbar_io_in_req_ready),
    .io_in_req_valid(mmioXbar_io_in_req_valid),
    .io_in_req_bits_addr(mmioXbar_io_in_req_bits_addr),
    .io_in_req_bits_size(mmioXbar_io_in_req_bits_size),
    .io_in_req_bits_cmd(mmioXbar_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(mmioXbar_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(mmioXbar_io_in_req_bits_wdata),
    .io_in_resp_ready(mmioXbar_io_in_resp_ready),
    .io_in_resp_valid(mmioXbar_io_in_resp_valid),
    .io_in_resp_bits_cmd(mmioXbar_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(mmioXbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(mmioXbar_io_out_0_req_ready),
    .io_out_0_req_valid(mmioXbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(mmioXbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_size(mmioXbar_io_out_0_req_bits_size),
    .io_out_0_req_bits_cmd(mmioXbar_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(mmioXbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(mmioXbar_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(mmioXbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(mmioXbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_cmd(mmioXbar_io_out_0_resp_bits_cmd),
    .io_out_0_resp_bits_rdata(mmioXbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(mmioXbar_io_out_1_req_ready),
    .io_out_1_req_valid(mmioXbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(mmioXbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_cmd(mmioXbar_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(mmioXbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(mmioXbar_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(mmioXbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(mmioXbar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(mmioXbar_io_out_1_resp_bits_rdata),
    .io_out_2_req_ready(mmioXbar_io_out_2_req_ready),
    .io_out_2_req_valid(mmioXbar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(mmioXbar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_cmd(mmioXbar_io_out_2_req_bits_cmd),
    .io_out_2_req_bits_wmask(mmioXbar_io_out_2_req_bits_wmask),
    .io_out_2_req_bits_wdata(mmioXbar_io_out_2_req_bits_wdata),
    .io_out_2_resp_ready(mmioXbar_io_out_2_resp_ready),
    .io_out_2_resp_valid(mmioXbar_io_out_2_resp_valid),
    .io_out_2_resp_bits_rdata(mmioXbar_io_out_2_resp_bits_rdata)
  );
  ysyx_210000_ReqBlocker ReqBlocker ( // @[NutShell.scala 120:25]
    .clock(ReqBlocker_clock),
    .reset(ReqBlocker_reset),
    .io_in_0_req_ready(ReqBlocker_io_in_0_req_ready),
    .io_in_0_req_valid(ReqBlocker_io_in_0_req_valid),
    .io_in_0_req_bits_addr(ReqBlocker_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(ReqBlocker_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(ReqBlocker_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(ReqBlocker_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(ReqBlocker_io_in_0_req_bits_wdata),
    .io_in_0_resp_ready(ReqBlocker_io_in_0_resp_ready),
    .io_in_0_resp_valid(ReqBlocker_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(ReqBlocker_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(ReqBlocker_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(ReqBlocker_io_in_1_req_ready),
    .io_in_1_req_valid(ReqBlocker_io_in_1_req_valid),
    .io_in_1_req_bits_addr(ReqBlocker_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(ReqBlocker_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(ReqBlocker_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(ReqBlocker_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(ReqBlocker_io_in_1_req_bits_wdata),
    .io_in_1_resp_ready(ReqBlocker_io_in_1_resp_ready),
    .io_in_1_resp_valid(ReqBlocker_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(ReqBlocker_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(ReqBlocker_io_in_1_resp_bits_rdata),
    .io_out_0_req_ready(ReqBlocker_io_out_0_req_ready),
    .io_out_0_req_valid(ReqBlocker_io_out_0_req_valid),
    .io_out_0_req_bits_addr(ReqBlocker_io_out_0_req_bits_addr),
    .io_out_0_req_bits_size(ReqBlocker_io_out_0_req_bits_size),
    .io_out_0_req_bits_cmd(ReqBlocker_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(ReqBlocker_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(ReqBlocker_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(ReqBlocker_io_out_0_resp_ready),
    .io_out_0_resp_valid(ReqBlocker_io_out_0_resp_valid),
    .io_out_0_resp_bits_cmd(ReqBlocker_io_out_0_resp_bits_cmd),
    .io_out_0_resp_bits_rdata(ReqBlocker_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(ReqBlocker_io_out_1_req_ready),
    .io_out_1_req_valid(ReqBlocker_io_out_1_req_valid),
    .io_out_1_req_bits_addr(ReqBlocker_io_out_1_req_bits_addr),
    .io_out_1_req_bits_size(ReqBlocker_io_out_1_req_bits_size),
    .io_out_1_req_bits_cmd(ReqBlocker_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(ReqBlocker_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(ReqBlocker_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(ReqBlocker_io_out_1_resp_ready),
    .io_out_1_resp_valid(ReqBlocker_io_out_1_resp_valid),
    .io_out_1_resp_bits_cmd(ReqBlocker_io_out_1_resp_bits_cmd),
    .io_out_1_resp_bits_rdata(ReqBlocker_io_out_1_resp_bits_rdata)
  );
  ysyx_210000_SimpleBusCrossbarNto1 SimpleBusCrossbarNto1 ( // @[NutShell.scala 121:28]
    .clock(SimpleBusCrossbarNto1_clock),
    .reset(SimpleBusCrossbarNto1_reset),
    .io_in_0_req_ready(SimpleBusCrossbarNto1_io_in_0_req_ready),
    .io_in_0_req_valid(SimpleBusCrossbarNto1_io_in_0_req_valid),
    .io_in_0_req_bits_addr(SimpleBusCrossbarNto1_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(SimpleBusCrossbarNto1_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(SimpleBusCrossbarNto1_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(SimpleBusCrossbarNto1_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(SimpleBusCrossbarNto1_io_in_0_req_bits_wdata),
    .io_in_0_resp_ready(SimpleBusCrossbarNto1_io_in_0_resp_ready),
    .io_in_0_resp_valid(SimpleBusCrossbarNto1_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(SimpleBusCrossbarNto1_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(SimpleBusCrossbarNto1_io_in_1_req_ready),
    .io_in_1_req_valid(SimpleBusCrossbarNto1_io_in_1_req_valid),
    .io_in_1_req_bits_addr(SimpleBusCrossbarNto1_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(SimpleBusCrossbarNto1_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(SimpleBusCrossbarNto1_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(SimpleBusCrossbarNto1_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(SimpleBusCrossbarNto1_io_in_1_req_bits_wdata),
    .io_in_1_resp_ready(SimpleBusCrossbarNto1_io_in_1_resp_ready),
    .io_in_1_resp_valid(SimpleBusCrossbarNto1_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(SimpleBusCrossbarNto1_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata),
    .io_out_req_ready(SimpleBusCrossbarNto1_io_out_req_ready),
    .io_out_req_valid(SimpleBusCrossbarNto1_io_out_req_valid),
    .io_out_req_bits_addr(SimpleBusCrossbarNto1_io_out_req_bits_addr),
    .io_out_req_bits_size(SimpleBusCrossbarNto1_io_out_req_bits_size),
    .io_out_req_bits_cmd(SimpleBusCrossbarNto1_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(SimpleBusCrossbarNto1_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(SimpleBusCrossbarNto1_io_out_req_bits_wdata),
    .io_out_resp_ready(SimpleBusCrossbarNto1_io_out_resp_ready),
    .io_out_resp_valid(SimpleBusCrossbarNto1_io_out_resp_valid),
    .io_out_resp_bits_cmd(SimpleBusCrossbarNto1_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(SimpleBusCrossbarNto1_io_out_resp_bits_rdata)
  );
  ysyx_210000_SimpleBus2AXI4Converter SimpleBus2AXI4Converter ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_clock),
    .reset(SimpleBus2AXI4Converter_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_io_in_req_bits_addr),
    .io_in_req_bits_size(SimpleBus2AXI4Converter_io_in_req_bits_size),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_io_in_resp_valid),
    .io_in_resp_bits_cmd(SimpleBus2AXI4Converter_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_io_out_awaddr),
    .io_out_awid(SimpleBus2AXI4Converter_io_out_awid),
    .io_out_awlen(SimpleBus2AXI4Converter_io_out_awlen),
    .io_out_awsize(SimpleBus2AXI4Converter_io_out_awsize),
    .io_out_awburst(SimpleBus2AXI4Converter_io_out_awburst),
    .io_out_wready(SimpleBus2AXI4Converter_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_io_out_wdata),
    .io_out_wstrb(SimpleBus2AXI4Converter_io_out_wstrb),
    .io_out_wlast(SimpleBus2AXI4Converter_io_out_wlast),
    .io_out_bready(SimpleBus2AXI4Converter_io_out_bready),
    .io_out_bvalid(SimpleBus2AXI4Converter_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_io_out_araddr),
    .io_out_arid(SimpleBus2AXI4Converter_io_out_arid),
    .io_out_arlen(SimpleBus2AXI4Converter_io_out_arlen),
    .io_out_arsize(SimpleBus2AXI4Converter_io_out_arsize),
    .io_out_arburst(SimpleBus2AXI4Converter_io_out_arburst),
    .io_out_rready(SimpleBus2AXI4Converter_io_out_rready),
    .io_out_rvalid(SimpleBus2AXI4Converter_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_io_out_rdata),
    .io_out_rlast(SimpleBus2AXI4Converter_io_out_rlast)
  );
  ysyx_210000_AXI4CLINT clint ( // @[NutShell.scala 129:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io__in_awready(clint_io__in_awready),
    .io__in_awvalid(clint_io__in_awvalid),
    .io__in_awaddr(clint_io__in_awaddr),
    .io__in_wready(clint_io__in_wready),
    .io__in_wvalid(clint_io__in_wvalid),
    .io__in_wdata(clint_io__in_wdata),
    .io__in_wstrb(clint_io__in_wstrb),
    .io__in_bready(clint_io__in_bready),
    .io__in_bvalid(clint_io__in_bvalid),
    .io__in_arready(clint_io__in_arready),
    .io__in_arvalid(clint_io__in_arvalid),
    .io__in_araddr(clint_io__in_araddr),
    .io__in_rready(clint_io__in_rready),
    .io__in_rvalid(clint_io__in_rvalid),
    .io__in_rdata(clint_io__in_rdata),
    .io__extra_mtip(clint_io__extra_mtip),
    .io__extra_msip(clint_io__extra_msip),
    .io_extra_mtip(clint_io_extra_mtip),
    .io_extra_msip(clint_io_extra_msip)
  );
  ysyx_210000_SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter_1 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_1_clock),
    .reset(SimpleBus2AXI4Converter_1_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_1_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_1_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_1_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_1_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_1_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_1_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_1_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_1_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_1_io_out_awaddr),
    .io_out_wready(SimpleBus2AXI4Converter_1_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_1_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_1_io_out_wdata),
    .io_out_wstrb(SimpleBus2AXI4Converter_1_io_out_wstrb),
    .io_out_bready(SimpleBus2AXI4Converter_1_io_out_bready),
    .io_out_bvalid(SimpleBus2AXI4Converter_1_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_1_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_1_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_1_io_out_araddr),
    .io_out_rready(SimpleBus2AXI4Converter_1_io_out_rready),
    .io_out_rvalid(SimpleBus2AXI4Converter_1_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_1_io_out_rdata)
  );
  ysyx_210000_AXI4PLIC plic ( // @[NutShell.scala 136:20]
    .clock(plic_clock),
    .reset(plic_reset),
    .io__in_awready(plic_io__in_awready),
    .io__in_awvalid(plic_io__in_awvalid),
    .io__in_awaddr(plic_io__in_awaddr),
    .io__in_wready(plic_io__in_wready),
    .io__in_wvalid(plic_io__in_wvalid),
    .io__in_wdata(plic_io__in_wdata),
    .io__in_wstrb(plic_io__in_wstrb),
    .io__in_bready(plic_io__in_bready),
    .io__in_bvalid(plic_io__in_bvalid),
    .io__in_arready(plic_io__in_arready),
    .io__in_arvalid(plic_io__in_arvalid),
    .io__in_araddr(plic_io__in_araddr),
    .io__in_rready(plic_io__in_rready),
    .io__in_rvalid(plic_io__in_rvalid),
    .io__in_rdata(plic_io__in_rdata),
    .io__extra_intrVec(plic_io__extra_intrVec),
    .io__extra_meip_0(plic_io__extra_meip_0),
    .io_extra_meip_0(plic_io_extra_meip_0)
  );
  ysyx_210000_SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter_2 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_2_clock),
    .reset(SimpleBus2AXI4Converter_2_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_2_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_2_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_2_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_2_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_2_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_2_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_2_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_2_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_2_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_2_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_2_io_out_awaddr),
    .io_out_wready(SimpleBus2AXI4Converter_2_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_2_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_2_io_out_wdata),
    .io_out_wstrb(SimpleBus2AXI4Converter_2_io_out_wstrb),
    .io_out_bready(SimpleBus2AXI4Converter_2_io_out_bready),
    .io_out_bvalid(SimpleBus2AXI4Converter_2_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_2_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_2_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_2_io_out_araddr),
    .io_out_rready(SimpleBus2AXI4Converter_2_io_out_rready),
    .io_out_rvalid(SimpleBus2AXI4Converter_2_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_2_io_out_rdata)
  );
  assign io_master_awvalid = SimpleBus2AXI4Converter_io_out_awvalid; // @[NutShell.scala 126:15]
  assign io_master_awaddr = SimpleBus2AXI4Converter_io_out_awaddr; // @[NutShell.scala 126:15]
  assign io_master_awid = SimpleBus2AXI4Converter_io_out_awid; // @[NutShell.scala 126:15]
  assign io_master_awlen = SimpleBus2AXI4Converter_io_out_awlen; // @[NutShell.scala 126:15]
  assign io_master_awsize = SimpleBus2AXI4Converter_io_out_awsize; // @[NutShell.scala 126:15]
  assign io_master_awburst = SimpleBus2AXI4Converter_io_out_awburst; // @[NutShell.scala 126:15]
  assign io_master_wvalid = SimpleBus2AXI4Converter_io_out_wvalid; // @[NutShell.scala 126:15]
  assign io_master_wdata = SimpleBus2AXI4Converter_io_out_wdata; // @[NutShell.scala 126:15]
  assign io_master_wstrb = SimpleBus2AXI4Converter_io_out_wstrb; // @[NutShell.scala 126:15]
  assign io_master_wlast = SimpleBus2AXI4Converter_io_out_wlast; // @[NutShell.scala 126:15]
  assign io_master_bready = SimpleBus2AXI4Converter_io_out_bready; // @[NutShell.scala 126:15]
  assign io_master_arvalid = SimpleBus2AXI4Converter_io_out_arvalid; // @[NutShell.scala 126:15]
  assign io_master_araddr = SimpleBus2AXI4Converter_io_out_araddr; // @[NutShell.scala 126:15]
  assign io_master_arid = 4'h0; // @[NutShell.scala 126:15]
  assign io_master_arlen = SimpleBus2AXI4Converter_io_out_arlen; // @[NutShell.scala 126:15]
  assign io_master_arsize = SimpleBus2AXI4Converter_io_out_arsize; // @[NutShell.scala 126:15]
  assign io_master_arburst = 2'h2; // @[NutShell.scala 126:15]
  assign io_master_rready = SimpleBus2AXI4Converter_io_out_rready; // @[NutShell.scala 126:15]
  assign io_slave_awready = axi2sb_io_in_awready; // @[NutShell.scala 63:16]
  assign io_slave_wready = axi2sb_io_in_wready; // @[NutShell.scala 63:16]
  assign io_slave_bvalid = axi2sb_io_in_bvalid; // @[NutShell.scala 63:16]
  assign io_slave_bresp = 2'h0; // @[NutShell.scala 63:16]
  assign io_slave_bid = 4'h0; // @[NutShell.scala 63:16]
  assign io_slave_arready = axi2sb_io_in_arready; // @[NutShell.scala 63:16]
  assign io_slave_rvalid = axi2sb_io_in_rvalid; // @[NutShell.scala 63:16]
  assign io_slave_rresp = 2'h0; // @[NutShell.scala 63:16]
  assign io_slave_rdata = axi2sb_io_in_rdata; // @[NutShell.scala 63:16]
  assign io_slave_rlast = axi2sb_io_in_rlast; // @[NutShell.scala 63:16]
  assign io_slave_rid = axi2sb_io_in_rid[3:0]; // @[NutShell.scala 63:16]
  assign nutcore_clock = clock;
  assign nutcore_reset = reset;
  assign nutcore_io_imem_mem_req_ready = cohMg_io_in_req_ready; // @[NutShell.scala 57:15]
  assign nutcore_io_imem_mem_resp_valid = cohMg_io_in_resp_valid; // @[NutShell.scala 57:15]
  assign nutcore_io_imem_mem_resp_bits_cmd = cohMg_io_in_resp_bits_cmd; // @[NutShell.scala 57:15]
  assign nutcore_io_imem_mem_resp_bits_rdata = cohMg_io_in_resp_bits_rdata; // @[NutShell.scala 57:15]
  assign nutcore_io_dmem_mem_req_ready = xbar_io_in_1_req_ready; // @[NutShell.scala 60:17]
  assign nutcore_io_dmem_mem_resp_valid = xbar_io_in_1_resp_valid; // @[NutShell.scala 60:17]
  assign nutcore_io_dmem_mem_resp_bits_cmd = xbar_io_in_1_resp_bits_cmd; // @[NutShell.scala 60:17]
  assign nutcore_io_dmem_mem_resp_bits_rdata = xbar_io_in_1_resp_bits_rdata; // @[NutShell.scala 60:17]
  assign nutcore_io_dmem_coh_req_valid = cohMg_io_out_coh_req_valid; // @[NutShell.scala 58:23]
  assign nutcore_io_dmem_coh_req_bits_addr = cohMg_io_out_coh_req_bits_addr; // @[NutShell.scala 58:23]
  assign nutcore_io_dmem_coh_req_bits_wdata = cohMg_io_out_coh_req_bits_wdata; // @[NutShell.scala 58:23]
  assign nutcore_io_mmio_req_ready = mmioXbar_io_in_req_ready; // @[NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_valid = mmioXbar_io_in_resp_valid; // @[NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_cmd = mmioXbar_io_in_resp_bits_cmd; // @[NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_rdata = mmioXbar_io_in_resp_bits_rdata; // @[NutShell.scala 107:18]
  assign nutcore_io_frontend_req_valid = axi2sb_io_out_req_valid; // @[NutShell.scala 64:23]
  assign nutcore_io_frontend_req_bits_addr = axi2sb_io_out_req_bits_addr; // @[NutShell.scala 64:23]
  assign nutcore_io_frontend_req_bits_size = axi2sb_io_out_req_bits_size; // @[NutShell.scala 64:23]
  assign nutcore_io_frontend_req_bits_cmd = axi2sb_io_out_req_bits_cmd; // @[NutShell.scala 64:23]
  assign nutcore_io_frontend_req_bits_wmask = axi2sb_io_out_req_bits_wmask; // @[NutShell.scala 64:23]
  assign nutcore_io_frontend_req_bits_wdata = axi2sb_io_out_req_bits_wdata; // @[NutShell.scala 64:23]
  assign nutcore_io_frontend_resp_ready = axi2sb_io_out_resp_ready; // @[NutShell.scala 64:23]
  assign nutcore_io_extra_mtip = clint_io_extra_mtip;
  assign nutcore_io_extra_meip_0 = plic_io_extra_meip_0;
  assign nutcore_io_extra_msip = clint_io_extra_msip;
  assign cohMg_clock = clock;
  assign cohMg_reset = reset;
  assign cohMg_io_in_req_valid = nutcore_io_imem_mem_req_valid; // @[NutShell.scala 57:15]
  assign cohMg_io_in_req_bits_addr = nutcore_io_imem_mem_req_bits_addr; // @[NutShell.scala 57:15]
  assign cohMg_io_in_req_bits_cmd = nutcore_io_imem_mem_req_bits_cmd; // @[NutShell.scala 57:15]
  assign cohMg_io_in_req_bits_wdata = nutcore_io_imem_mem_req_bits_wdata; // @[NutShell.scala 57:15]
  assign cohMg_io_out_mem_req_ready = xbar_io_in_0_req_ready; // @[NutShell.scala 59:17]
  assign cohMg_io_out_mem_resp_valid = xbar_io_in_0_resp_valid; // @[NutShell.scala 59:17]
  assign cohMg_io_out_mem_resp_bits_cmd = xbar_io_in_0_resp_bits_cmd; // @[NutShell.scala 59:17]
  assign cohMg_io_out_mem_resp_bits_rdata = xbar_io_in_0_resp_bits_rdata; // @[NutShell.scala 59:17]
  assign cohMg_io_out_coh_req_ready = nutcore_io_dmem_coh_req_ready; // @[NutShell.scala 58:23]
  assign cohMg_io_out_coh_resp_valid = nutcore_io_dmem_coh_resp_valid; // @[NutShell.scala 58:23]
  assign cohMg_io_out_coh_resp_bits_cmd = nutcore_io_dmem_coh_resp_bits_cmd; // @[NutShell.scala 58:23]
  assign cohMg_io_out_coh_resp_bits_rdata = nutcore_io_dmem_coh_resp_bits_rdata; // @[NutShell.scala 58:23]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_in_0_req_valid = cohMg_io_out_mem_req_valid; // @[NutShell.scala 59:17]
  assign xbar_io_in_0_req_bits_addr = cohMg_io_out_mem_req_bits_addr; // @[NutShell.scala 59:17]
  assign xbar_io_in_0_req_bits_size = cohMg_io_out_mem_req_bits_size; // @[NutShell.scala 59:17]
  assign xbar_io_in_0_req_bits_cmd = cohMg_io_out_mem_req_bits_cmd; // @[NutShell.scala 59:17]
  assign xbar_io_in_0_req_bits_wmask = cohMg_io_out_mem_req_bits_wmask; // @[NutShell.scala 59:17]
  assign xbar_io_in_0_req_bits_wdata = cohMg_io_out_mem_req_bits_wdata; // @[NutShell.scala 59:17]
  assign xbar_io_in_0_resp_ready = 1'h1; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_valid = nutcore_io_dmem_mem_req_valid; // @[NutShell.scala 60:17]
  assign xbar_io_in_1_req_bits_addr = nutcore_io_dmem_mem_req_bits_addr; // @[NutShell.scala 60:17]
  assign xbar_io_in_1_req_bits_size = 3'h3; // @[NutShell.scala 60:17]
  assign xbar_io_in_1_req_bits_cmd = nutcore_io_dmem_mem_req_bits_cmd; // @[NutShell.scala 60:17]
  assign xbar_io_in_1_req_bits_wmask = 8'hff; // @[NutShell.scala 60:17]
  assign xbar_io_in_1_req_bits_wdata = nutcore_io_dmem_mem_req_bits_wdata; // @[NutShell.scala 60:17]
  assign xbar_io_in_1_resp_ready = 1'h1; // @[NutShell.scala 60:17]
  assign xbar_io_out_req_ready = memAddrMap_io_in_req_ready; // @[NutShell.scala 95:20]
  assign xbar_io_out_resp_valid = memAddrMap_io_in_resp_valid; // @[NutShell.scala 95:20]
  assign xbar_io_out_resp_bits_cmd = memAddrMap_io_in_resp_bits_cmd; // @[NutShell.scala 95:20]
  assign xbar_io_out_resp_bits_rdata = memAddrMap_io_in_resp_bits_rdata; // @[NutShell.scala 95:20]
  assign axi2sb_clock = clock;
  assign axi2sb_reset = reset;
  assign axi2sb_io_in_awvalid = io_slave_awvalid; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_awaddr = io_slave_awaddr; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_awid = {{14'd0}, io_slave_awid}; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_awlen = io_slave_awlen; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_awsize = io_slave_awsize; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_wvalid = io_slave_wvalid; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_wdata = io_slave_wdata; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_wstrb = io_slave_wstrb; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_wlast = io_slave_wlast; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_bready = io_slave_bready; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_arvalid = io_slave_arvalid; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_araddr = io_slave_araddr; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_arid = {{14'd0}, io_slave_arid}; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_arlen = io_slave_arlen; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_arsize = io_slave_arsize; // @[NutShell.scala 63:16]
  assign axi2sb_io_in_rready = io_slave_rready; // @[NutShell.scala 63:16]
  assign axi2sb_io_out_req_ready = nutcore_io_frontend_req_ready; // @[NutShell.scala 64:23]
  assign axi2sb_io_out_resp_valid = nutcore_io_frontend_resp_valid; // @[NutShell.scala 64:23]
  assign axi2sb_io_out_resp_bits_cmd = nutcore_io_frontend_resp_bits_cmd; // @[NutShell.scala 64:23]
  assign axi2sb_io_out_resp_bits_rdata = nutcore_io_frontend_resp_bits_rdata; // @[NutShell.scala 64:23]
  assign memAddrMap_io_in_req_valid = xbar_io_out_req_valid; // @[NutShell.scala 95:20]
  assign memAddrMap_io_in_req_bits_addr = xbar_io_out_req_bits_addr; // @[NutShell.scala 95:20]
  assign memAddrMap_io_in_req_bits_size = xbar_io_out_req_bits_size; // @[NutShell.scala 95:20]
  assign memAddrMap_io_in_req_bits_cmd = xbar_io_out_req_bits_cmd; // @[NutShell.scala 95:20]
  assign memAddrMap_io_in_req_bits_wmask = xbar_io_out_req_bits_wmask; // @[NutShell.scala 95:20]
  assign memAddrMap_io_in_req_bits_wdata = xbar_io_out_req_bits_wdata; // @[NutShell.scala 95:20]
  assign memAddrMap_io_in_resp_ready = xbar_io_out_resp_ready; // @[NutShell.scala 95:20]
  assign memAddrMap_io_out_req_ready = ReqBlocker_io_in_0_req_ready; // @[NutShell.scala 122:22]
  assign memAddrMap_io_out_resp_valid = ReqBlocker_io_in_0_resp_valid; // @[NutShell.scala 122:22]
  assign memAddrMap_io_out_resp_bits_cmd = ReqBlocker_io_in_0_resp_bits_cmd; // @[NutShell.scala 122:22]
  assign memAddrMap_io_out_resp_bits_rdata = ReqBlocker_io_in_0_resp_bits_rdata; // @[NutShell.scala 122:22]
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_req_valid = nutcore_io_mmio_req_valid; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_addr = nutcore_io_mmio_req_bits_addr; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_size = nutcore_io_mmio_req_bits_size; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_cmd = nutcore_io_mmio_req_bits_cmd; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wmask = nutcore_io_mmio_req_bits_wmask; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wdata = nutcore_io_mmio_req_bits_wdata; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_resp_ready = nutcore_io_mmio_resp_ready; // @[NutShell.scala 107:18]
  assign mmioXbar_io_out_0_req_ready = ReqBlocker_io_in_1_req_ready; // @[NutShell.scala 123:22]
  assign mmioXbar_io_out_0_resp_valid = ReqBlocker_io_in_1_resp_valid; // @[NutShell.scala 123:22]
  assign mmioXbar_io_out_0_resp_bits_cmd = ReqBlocker_io_in_1_resp_bits_cmd; // @[NutShell.scala 123:22]
  assign mmioXbar_io_out_0_resp_bits_rdata = ReqBlocker_io_in_1_resp_bits_rdata; // @[NutShell.scala 123:22]
  assign mmioXbar_io_out_1_req_ready = SimpleBus2AXI4Converter_1_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_valid = SimpleBus2AXI4Converter_1_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_bits_rdata = SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_req_ready = SimpleBus2AXI4Converter_2_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_resp_valid = SimpleBus2AXI4Converter_2_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_resp_bits_rdata = SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign ReqBlocker_clock = clock;
  assign ReqBlocker_reset = reset;
  assign ReqBlocker_io_in_0_req_valid = memAddrMap_io_out_req_valid; // @[NutShell.scala 122:22]
  assign ReqBlocker_io_in_0_req_bits_addr = memAddrMap_io_out_req_bits_addr; // @[NutShell.scala 122:22]
  assign ReqBlocker_io_in_0_req_bits_size = memAddrMap_io_out_req_bits_size; // @[NutShell.scala 122:22]
  assign ReqBlocker_io_in_0_req_bits_cmd = memAddrMap_io_out_req_bits_cmd; // @[NutShell.scala 122:22]
  assign ReqBlocker_io_in_0_req_bits_wmask = memAddrMap_io_out_req_bits_wmask; // @[NutShell.scala 122:22]
  assign ReqBlocker_io_in_0_req_bits_wdata = memAddrMap_io_out_req_bits_wdata; // @[NutShell.scala 122:22]
  assign ReqBlocker_io_in_0_resp_ready = memAddrMap_io_out_resp_ready; // @[NutShell.scala 122:22]
  assign ReqBlocker_io_in_1_req_valid = mmioXbar_io_out_0_req_valid; // @[NutShell.scala 123:22]
  assign ReqBlocker_io_in_1_req_bits_addr = mmioXbar_io_out_0_req_bits_addr; // @[NutShell.scala 123:22]
  assign ReqBlocker_io_in_1_req_bits_size = mmioXbar_io_out_0_req_bits_size; // @[NutShell.scala 123:22]
  assign ReqBlocker_io_in_1_req_bits_cmd = mmioXbar_io_out_0_req_bits_cmd; // @[NutShell.scala 123:22]
  assign ReqBlocker_io_in_1_req_bits_wmask = mmioXbar_io_out_0_req_bits_wmask; // @[NutShell.scala 123:22]
  assign ReqBlocker_io_in_1_req_bits_wdata = mmioXbar_io_out_0_req_bits_wdata; // @[NutShell.scala 123:22]
  assign ReqBlocker_io_in_1_resp_ready = mmioXbar_io_out_0_resp_ready; // @[NutShell.scala 123:22]
  assign ReqBlocker_io_out_0_req_ready = SimpleBusCrossbarNto1_io_in_0_req_ready; // @[NutShell.scala 124:25]
  assign ReqBlocker_io_out_0_resp_valid = SimpleBusCrossbarNto1_io_in_0_resp_valid; // @[NutShell.scala 124:25]
  assign ReqBlocker_io_out_0_resp_bits_cmd = SimpleBusCrossbarNto1_io_in_0_resp_bits_cmd; // @[NutShell.scala 124:25]
  assign ReqBlocker_io_out_0_resp_bits_rdata = SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata; // @[NutShell.scala 124:25]
  assign ReqBlocker_io_out_1_req_ready = SimpleBusCrossbarNto1_io_in_1_req_ready; // @[NutShell.scala 125:25]
  assign ReqBlocker_io_out_1_resp_valid = SimpleBusCrossbarNto1_io_in_1_resp_valid; // @[NutShell.scala 125:25]
  assign ReqBlocker_io_out_1_resp_bits_cmd = SimpleBusCrossbarNto1_io_in_1_resp_bits_cmd; // @[NutShell.scala 125:25]
  assign ReqBlocker_io_out_1_resp_bits_rdata = SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata; // @[NutShell.scala 125:25]
  assign SimpleBusCrossbarNto1_clock = clock;
  assign SimpleBusCrossbarNto1_reset = reset;
  assign SimpleBusCrossbarNto1_io_in_0_req_valid = ReqBlocker_io_out_0_req_valid; // @[NutShell.scala 124:25]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_addr = ReqBlocker_io_out_0_req_bits_addr; // @[NutShell.scala 124:25]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_size = ReqBlocker_io_out_0_req_bits_size; // @[NutShell.scala 124:25]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_cmd = ReqBlocker_io_out_0_req_bits_cmd; // @[NutShell.scala 124:25]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_wmask = ReqBlocker_io_out_0_req_bits_wmask; // @[NutShell.scala 124:25]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_wdata = ReqBlocker_io_out_0_req_bits_wdata; // @[NutShell.scala 124:25]
  assign SimpleBusCrossbarNto1_io_in_0_resp_ready = ReqBlocker_io_out_0_resp_ready; // @[NutShell.scala 124:25]
  assign SimpleBusCrossbarNto1_io_in_1_req_valid = ReqBlocker_io_out_1_req_valid; // @[NutShell.scala 125:25]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_addr = ReqBlocker_io_out_1_req_bits_addr; // @[NutShell.scala 125:25]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_size = ReqBlocker_io_out_1_req_bits_size; // @[NutShell.scala 125:25]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_cmd = ReqBlocker_io_out_1_req_bits_cmd; // @[NutShell.scala 125:25]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_wmask = ReqBlocker_io_out_1_req_bits_wmask; // @[NutShell.scala 125:25]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_wdata = ReqBlocker_io_out_1_req_bits_wdata; // @[NutShell.scala 125:25]
  assign SimpleBusCrossbarNto1_io_in_1_resp_ready = ReqBlocker_io_out_1_resp_ready; // @[NutShell.scala 125:25]
  assign SimpleBusCrossbarNto1_io_out_req_ready = SimpleBus2AXI4Converter_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBusCrossbarNto1_io_out_resp_valid = SimpleBus2AXI4Converter_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBusCrossbarNto1_io_out_resp_bits_cmd = SimpleBus2AXI4Converter_io_in_resp_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBusCrossbarNto1_io_out_resp_bits_rdata = SimpleBus2AXI4Converter_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_clock = clock;
  assign SimpleBus2AXI4Converter_reset = reset;
  assign SimpleBus2AXI4Converter_io_in_req_valid = SimpleBusCrossbarNto1_io_out_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_addr = SimpleBusCrossbarNto1_io_out_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_size = SimpleBusCrossbarNto1_io_out_req_bits_size; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_cmd = SimpleBusCrossbarNto1_io_out_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_wmask = SimpleBusCrossbarNto1_io_out_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_wdata = SimpleBusCrossbarNto1_io_out_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_resp_ready = SimpleBusCrossbarNto1_io_out_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_out_awready = io_master_awready; // @[NutShell.scala 126:15]
  assign SimpleBus2AXI4Converter_io_out_wready = io_master_wready; // @[NutShell.scala 126:15]
  assign SimpleBus2AXI4Converter_io_out_bvalid = io_master_bvalid; // @[NutShell.scala 126:15]
  assign SimpleBus2AXI4Converter_io_out_arready = io_master_arready; // @[NutShell.scala 126:15]
  assign SimpleBus2AXI4Converter_io_out_rvalid = io_master_rvalid; // @[NutShell.scala 126:15]
  assign SimpleBus2AXI4Converter_io_out_rdata = io_master_rdata; // @[NutShell.scala 126:15]
  assign SimpleBus2AXI4Converter_io_out_rlast = io_master_rlast; // @[NutShell.scala 126:15]
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io__in_awvalid = SimpleBus2AXI4Converter_1_io_out_awvalid; // @[NutShell.scala 130:15]
  assign clint_io__in_awaddr = SimpleBus2AXI4Converter_1_io_out_awaddr; // @[NutShell.scala 130:15]
  assign clint_io__in_wvalid = SimpleBus2AXI4Converter_1_io_out_wvalid; // @[NutShell.scala 130:15]
  assign clint_io__in_wdata = SimpleBus2AXI4Converter_1_io_out_wdata; // @[NutShell.scala 130:15]
  assign clint_io__in_wstrb = SimpleBus2AXI4Converter_1_io_out_wstrb; // @[NutShell.scala 130:15]
  assign clint_io__in_bready = SimpleBus2AXI4Converter_1_io_out_bready; // @[NutShell.scala 130:15]
  assign clint_io__in_arvalid = SimpleBus2AXI4Converter_1_io_out_arvalid; // @[NutShell.scala 130:15]
  assign clint_io__in_araddr = SimpleBus2AXI4Converter_1_io_out_araddr; // @[NutShell.scala 130:15]
  assign clint_io__in_rready = SimpleBus2AXI4Converter_1_io_out_rready; // @[NutShell.scala 130:15]
  assign SimpleBus2AXI4Converter_1_clock = clock;
  assign SimpleBus2AXI4Converter_1_reset = reset;
  assign SimpleBus2AXI4Converter_1_io_in_req_valid = mmioXbar_io_out_1_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_addr = mmioXbar_io_out_1_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_cmd = mmioXbar_io_out_1_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_wmask = mmioXbar_io_out_1_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_wdata = mmioXbar_io_out_1_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_resp_ready = mmioXbar_io_out_1_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_out_awready = clint_io__in_awready; // @[NutShell.scala 130:15]
  assign SimpleBus2AXI4Converter_1_io_out_wready = clint_io__in_wready; // @[NutShell.scala 130:15]
  assign SimpleBus2AXI4Converter_1_io_out_bvalid = clint_io__in_bvalid; // @[NutShell.scala 130:15]
  assign SimpleBus2AXI4Converter_1_io_out_arready = clint_io__in_arready; // @[NutShell.scala 130:15]
  assign SimpleBus2AXI4Converter_1_io_out_rvalid = clint_io__in_rvalid; // @[NutShell.scala 130:15]
  assign SimpleBus2AXI4Converter_1_io_out_rdata = clint_io__in_rdata; // @[NutShell.scala 130:15]
  assign plic_clock = clock;
  assign plic_reset = reset;
  assign plic_io__in_awvalid = SimpleBus2AXI4Converter_2_io_out_awvalid; // @[NutShell.scala 137:14]
  assign plic_io__in_awaddr = SimpleBus2AXI4Converter_2_io_out_awaddr; // @[NutShell.scala 137:14]
  assign plic_io__in_wvalid = SimpleBus2AXI4Converter_2_io_out_wvalid; // @[NutShell.scala 137:14]
  assign plic_io__in_wdata = SimpleBus2AXI4Converter_2_io_out_wdata; // @[NutShell.scala 137:14]
  assign plic_io__in_wstrb = SimpleBus2AXI4Converter_2_io_out_wstrb; // @[NutShell.scala 137:14]
  assign plic_io__in_bready = SimpleBus2AXI4Converter_2_io_out_bready; // @[NutShell.scala 137:14]
  assign plic_io__in_arvalid = SimpleBus2AXI4Converter_2_io_out_arvalid; // @[NutShell.scala 137:14]
  assign plic_io__in_araddr = SimpleBus2AXI4Converter_2_io_out_araddr; // @[NutShell.scala 137:14]
  assign plic_io__in_rready = SimpleBus2AXI4Converter_2_io_out_rready; // @[NutShell.scala 137:14]
  assign plic_io__extra_intrVec = REG_1; // @[NutShell.scala 138:29]
  assign SimpleBus2AXI4Converter_2_clock = clock;
  assign SimpleBus2AXI4Converter_2_reset = reset;
  assign SimpleBus2AXI4Converter_2_io_in_req_valid = mmioXbar_io_out_2_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_addr = mmioXbar_io_out_2_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_cmd = mmioXbar_io_out_2_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_wmask = mmioXbar_io_out_2_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_wdata = mmioXbar_io_out_2_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_resp_ready = mmioXbar_io_out_2_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_out_awready = plic_io__in_awready; // @[NutShell.scala 137:14]
  assign SimpleBus2AXI4Converter_2_io_out_wready = plic_io__in_wready; // @[NutShell.scala 137:14]
  assign SimpleBus2AXI4Converter_2_io_out_bvalid = plic_io__in_bvalid; // @[NutShell.scala 137:14]
  assign SimpleBus2AXI4Converter_2_io_out_arready = plic_io__in_arready; // @[NutShell.scala 137:14]
  assign SimpleBus2AXI4Converter_2_io_out_rvalid = plic_io__in_rvalid; // @[NutShell.scala 137:14]
  assign SimpleBus2AXI4Converter_2_io_out_rdata = plic_io__in_rdata; // @[NutShell.scala 137:14]
  always @(posedge clock) begin
    if (reset) begin // @[NutShell.scala 138:47]
      REG <= 1'h0; // @[NutShell.scala 138:47]
    end else begin
      REG <= io_interrupt; // @[NutShell.scala 138:47]
    end
    if (reset) begin // @[NutShell.scala 138:39]
      REG_1 <= 1'h0; // @[NutShell.scala 138:39]
    end else begin
      REG_1 <= REG; // @[NutShell.scala 138:39]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210000_Top(
  input   clock,
  input   reset
);
  wire  nutshell_clock; // @[TopMain.scala 28:24]
  wire  nutshell_reset; // @[TopMain.scala 28:24]
  wire  nutshell_io_master_awready; // @[TopMain.scala 28:24]
  wire  nutshell_io_master_awvalid; // @[TopMain.scala 28:24]
  wire [31:0] nutshell_io_master_awaddr; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_master_awid; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_master_awlen; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_master_awsize; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_master_awburst; // @[TopMain.scala 28:24]
  wire  nutshell_io_master_wready; // @[TopMain.scala 28:24]
  wire  nutshell_io_master_wvalid; // @[TopMain.scala 28:24]
  wire [63:0] nutshell_io_master_wdata; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_master_wstrb; // @[TopMain.scala 28:24]
  wire  nutshell_io_master_wlast; // @[TopMain.scala 28:24]
  wire  nutshell_io_master_bready; // @[TopMain.scala 28:24]
  wire  nutshell_io_master_bvalid; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_master_bresp; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_master_bid; // @[TopMain.scala 28:24]
  wire  nutshell_io_master_arready; // @[TopMain.scala 28:24]
  wire  nutshell_io_master_arvalid; // @[TopMain.scala 28:24]
  wire [31:0] nutshell_io_master_araddr; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_master_arid; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_master_arlen; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_master_arsize; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_master_arburst; // @[TopMain.scala 28:24]
  wire  nutshell_io_master_rready; // @[TopMain.scala 28:24]
  wire  nutshell_io_master_rvalid; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_master_rresp; // @[TopMain.scala 28:24]
  wire [63:0] nutshell_io_master_rdata; // @[TopMain.scala 28:24]
  wire  nutshell_io_master_rlast; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_master_rid; // @[TopMain.scala 28:24]
  wire  nutshell_io_slave_awready; // @[TopMain.scala 28:24]
  wire  nutshell_io_slave_awvalid; // @[TopMain.scala 28:24]
  wire [31:0] nutshell_io_slave_awaddr; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_slave_awid; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_slave_awlen; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_slave_awsize; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_slave_awburst; // @[TopMain.scala 28:24]
  wire  nutshell_io_slave_wready; // @[TopMain.scala 28:24]
  wire  nutshell_io_slave_wvalid; // @[TopMain.scala 28:24]
  wire [63:0] nutshell_io_slave_wdata; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_slave_wstrb; // @[TopMain.scala 28:24]
  wire  nutshell_io_slave_wlast; // @[TopMain.scala 28:24]
  wire  nutshell_io_slave_bready; // @[TopMain.scala 28:24]
  wire  nutshell_io_slave_bvalid; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_slave_bresp; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_slave_bid; // @[TopMain.scala 28:24]
  wire  nutshell_io_slave_arready; // @[TopMain.scala 28:24]
  wire  nutshell_io_slave_arvalid; // @[TopMain.scala 28:24]
  wire [31:0] nutshell_io_slave_araddr; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_slave_arid; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_slave_arlen; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_slave_arsize; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_slave_arburst; // @[TopMain.scala 28:24]
  wire  nutshell_io_slave_rready; // @[TopMain.scala 28:24]
  wire  nutshell_io_slave_rvalid; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_slave_rresp; // @[TopMain.scala 28:24]
  wire [63:0] nutshell_io_slave_rdata; // @[TopMain.scala 28:24]
  wire  nutshell_io_slave_rlast; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_slave_rid; // @[TopMain.scala 28:24]
  wire  nutshell_io_interrupt; // @[TopMain.scala 28:24]
  ysyx_210000 nutshell ( // @[TopMain.scala 28:24]
    .clock(nutshell_clock),
    .reset(nutshell_reset),
    .io_master_awready(nutshell_io_master_awready),
    .io_master_awvalid(nutshell_io_master_awvalid),
    .io_master_awaddr(nutshell_io_master_awaddr),
    .io_master_awid(nutshell_io_master_awid),
    .io_master_awlen(nutshell_io_master_awlen),
    .io_master_awsize(nutshell_io_master_awsize),
    .io_master_awburst(nutshell_io_master_awburst),
    .io_master_wready(nutshell_io_master_wready),
    .io_master_wvalid(nutshell_io_master_wvalid),
    .io_master_wdata(nutshell_io_master_wdata),
    .io_master_wstrb(nutshell_io_master_wstrb),
    .io_master_wlast(nutshell_io_master_wlast),
    .io_master_bready(nutshell_io_master_bready),
    .io_master_bvalid(nutshell_io_master_bvalid),
    .io_master_bresp(nutshell_io_master_bresp),
    .io_master_bid(nutshell_io_master_bid),
    .io_master_arready(nutshell_io_master_arready),
    .io_master_arvalid(nutshell_io_master_arvalid),
    .io_master_araddr(nutshell_io_master_araddr),
    .io_master_arid(nutshell_io_master_arid),
    .io_master_arlen(nutshell_io_master_arlen),
    .io_master_arsize(nutshell_io_master_arsize),
    .io_master_arburst(nutshell_io_master_arburst),
    .io_master_rready(nutshell_io_master_rready),
    .io_master_rvalid(nutshell_io_master_rvalid),
    .io_master_rresp(nutshell_io_master_rresp),
    .io_master_rdata(nutshell_io_master_rdata),
    .io_master_rlast(nutshell_io_master_rlast),
    .io_master_rid(nutshell_io_master_rid),
    .io_slave_awready(nutshell_io_slave_awready),
    .io_slave_awvalid(nutshell_io_slave_awvalid),
    .io_slave_awaddr(nutshell_io_slave_awaddr),
    .io_slave_awid(nutshell_io_slave_awid),
    .io_slave_awlen(nutshell_io_slave_awlen),
    .io_slave_awsize(nutshell_io_slave_awsize),
    .io_slave_awburst(nutshell_io_slave_awburst),
    .io_slave_wready(nutshell_io_slave_wready),
    .io_slave_wvalid(nutshell_io_slave_wvalid),
    .io_slave_wdata(nutshell_io_slave_wdata),
    .io_slave_wstrb(nutshell_io_slave_wstrb),
    .io_slave_wlast(nutshell_io_slave_wlast),
    .io_slave_bready(nutshell_io_slave_bready),
    .io_slave_bvalid(nutshell_io_slave_bvalid),
    .io_slave_bresp(nutshell_io_slave_bresp),
    .io_slave_bid(nutshell_io_slave_bid),
    .io_slave_arready(nutshell_io_slave_arready),
    .io_slave_arvalid(nutshell_io_slave_arvalid),
    .io_slave_araddr(nutshell_io_slave_araddr),
    .io_slave_arid(nutshell_io_slave_arid),
    .io_slave_arlen(nutshell_io_slave_arlen),
    .io_slave_arsize(nutshell_io_slave_arsize),
    .io_slave_arburst(nutshell_io_slave_arburst),
    .io_slave_rready(nutshell_io_slave_rready),
    .io_slave_rvalid(nutshell_io_slave_rvalid),
    .io_slave_rresp(nutshell_io_slave_rresp),
    .io_slave_rdata(nutshell_io_slave_rdata),
    .io_slave_rlast(nutshell_io_slave_rlast),
    .io_slave_rid(nutshell_io_slave_rid),
    .io_interrupt(nutshell_io_interrupt)
  );
  assign nutshell_clock = clock;
  assign nutshell_reset = reset;
  assign nutshell_io_master_awready = 1'h0;
  assign nutshell_io_master_wready = 1'h0;
  assign nutshell_io_master_bvalid = 1'h0;
  assign nutshell_io_master_bresp = 2'h0;
  assign nutshell_io_master_bid = 4'h0;
  assign nutshell_io_master_arready = 1'h0;
  assign nutshell_io_master_rvalid = 1'h0;
  assign nutshell_io_master_rresp = 2'h0;
  assign nutshell_io_master_rdata = 64'h0;
  assign nutshell_io_master_rlast = 1'h0;
  assign nutshell_io_master_rid = 4'h0;
  assign nutshell_io_slave_awvalid = 1'h0;
  assign nutshell_io_slave_awaddr = 32'h0;
  assign nutshell_io_slave_awid = 4'h0;
  assign nutshell_io_slave_awlen = 8'h0;
  assign nutshell_io_slave_awsize = 3'h0;
  assign nutshell_io_slave_awburst = 2'h0;
  assign nutshell_io_slave_wvalid = 1'h0;
  assign nutshell_io_slave_wdata = 64'h0;
  assign nutshell_io_slave_wstrb = 8'h0;
  assign nutshell_io_slave_wlast = 1'h0;
  assign nutshell_io_slave_bready = 1'h0;
  assign nutshell_io_slave_arvalid = 1'h0;
  assign nutshell_io_slave_araddr = 32'h0;
  assign nutshell_io_slave_arid = 4'h0;
  assign nutshell_io_slave_arlen = 8'h0;
  assign nutshell_io_slave_arsize = 3'h0;
  assign nutshell_io_slave_arburst = 2'h0;
  assign nutshell_io_slave_rready = 1'h0;
  assign nutshell_io_interrupt = 1'h0;
endmodule
module ysyx_210000_array(
  input  [4:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [76:0] RW0_wdata_0,
  output [76:0] RW0_rdata_0
);
  wire [4:0] array_ext_RW0_addr;
  wire  array_ext_RW0_en;
  wire  array_ext_RW0_clk;
  wire  array_ext_RW0_wmode;
  wire [76:0] array_ext_RW0_wdata;
  wire [76:0] array_ext_RW0_rdata;
  array_ext array_ext (
    .RW0_addr(array_ext_RW0_addr),
    .RW0_en(array_ext_RW0_en),
    .RW0_clk(array_ext_RW0_clk),
    .RW0_wmode(array_ext_RW0_wmode),
    .RW0_wdata(array_ext_RW0_wdata),
    .RW0_rdata(array_ext_RW0_rdata)
  );
  assign array_ext_RW0_clk = RW0_clk;
  assign array_ext_RW0_en = RW0_en;
  assign array_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_ext_RW0_rdata;
  assign array_ext_RW0_wmode = RW0_wmode;
  assign array_ext_RW0_wdata = RW0_wdata_0;
endmodule
module ysyx_210000_array_0(
  input  [3:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [23:0] RW0_wdata_0,
  input  [23:0] RW0_wdata_1,
  input  [23:0] RW0_wdata_2,
  input  [23:0] RW0_wdata_3,
  output [23:0] RW0_rdata_0,
  output [23:0] RW0_rdata_1,
  output [23:0] RW0_rdata_2,
  output [23:0] RW0_rdata_3,
  input         RW0_wmask_0,
  input         RW0_wmask_1,
  input         RW0_wmask_2,
  input         RW0_wmask_3
);
  wire [3:0] array_0_ext_RW0_addr;
  wire  array_0_ext_RW0_en;
  wire  array_0_ext_RW0_clk;
  wire  array_0_ext_RW0_wmode;
  wire [95:0] array_0_ext_RW0_wdata;
  wire [95:0] array_0_ext_RW0_rdata;
  wire [3:0] array_0_ext_RW0_wmask;
  wire [47:0] _GEN_0 = {RW0_wdata_3,RW0_wdata_2};
  wire [47:0] _GEN_1 = {RW0_wdata_1,RW0_wdata_0};
  wire [1:0] _GEN_2 = {RW0_wmask_3,RW0_wmask_2};
  wire [1:0] _GEN_3 = {RW0_wmask_1,RW0_wmask_0};
  array_0_ext array_0_ext (
    .RW0_addr(array_0_ext_RW0_addr),
    .RW0_en(array_0_ext_RW0_en),
    .RW0_clk(array_0_ext_RW0_clk),
    .RW0_wmode(array_0_ext_RW0_wmode),
    .RW0_wdata(array_0_ext_RW0_wdata),
    .RW0_rdata(array_0_ext_RW0_rdata),
    .RW0_wmask(array_0_ext_RW0_wmask)
  );
  assign array_0_ext_RW0_clk = RW0_clk;
  assign array_0_ext_RW0_en = RW0_en;
  assign array_0_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_0_ext_RW0_rdata[23:0];
  assign RW0_rdata_1 = array_0_ext_RW0_rdata[47:24];
  assign RW0_rdata_2 = array_0_ext_RW0_rdata[71:48];
  assign RW0_rdata_3 = array_0_ext_RW0_rdata[95:72];
  assign array_0_ext_RW0_wmode = RW0_wmode;
  assign array_0_ext_RW0_wdata = {_GEN_0,_GEN_1};
  assign array_0_ext_RW0_wmask = {_GEN_2,_GEN_3};
endmodule

module array_ext(
  input RW0_clk,
  input [4:0] RW0_addr,
  input RW0_en,
  input RW0_wmode,
  input [76:0] RW0_wdata,
  output [76:0] RW0_rdata
);

  reg reg_RW0_ren;
  reg [4:0] reg_RW0_addr;
  reg [76:0] ram [31:0];
  `ifdef RANDOMIZE_MEM_INIT
    integer initvar;
    initial begin
      #`RANDOMIZE_DELAY begin end
      for (initvar = 0; initvar < 32; initvar = initvar+1)
        ram[initvar] = {3 {$random}};
      reg_RW0_addr = {1 {$random}};
    end
  `endif
  integer i;
  always @(posedge RW0_clk)
    reg_RW0_ren <= RW0_en && !RW0_wmode;
  always @(posedge RW0_clk)
    if (RW0_en && !RW0_wmode) reg_RW0_addr <= RW0_addr;
  always @(posedge RW0_clk)
    if (RW0_en && RW0_wmode) begin
      for(i=0;i<1;i=i+1) begin
        ram[RW0_addr][i*77 +: 77] <= RW0_wdata[i*77 +: 77];
      end
    end
  `ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [95:0] RW0_random;
  `ifdef RANDOMIZE_MEM_INIT
    initial begin
      #`RANDOMIZE_DELAY begin end
      RW0_random = {$random, $random, $random};
      reg_RW0_ren = RW0_random[0];
    end
  `endif
  always @(posedge RW0_clk) RW0_random <= {$random, $random, $random};
  assign RW0_rdata = reg_RW0_ren ? ram[reg_RW0_addr] : RW0_random[76:0];
  `else
  assign RW0_rdata = ram[reg_RW0_addr];
  `endif

endmodule

module array_0_ext(
  input RW0_clk,
  input [3:0] RW0_addr,
  input RW0_en,
  input RW0_wmode,
  input [3:0] RW0_wmask,
  input [95:0] RW0_wdata,
  output [95:0] RW0_rdata
);

  reg reg_RW0_ren;
  reg [3:0] reg_RW0_addr;
  reg [95:0] ram [15:0];
  `ifdef RANDOMIZE_MEM_INIT
    integer initvar;
    initial begin
      #`RANDOMIZE_DELAY begin end
      for (initvar = 0; initvar < 16; initvar = initvar+1)
        ram[initvar] = {3 {$random}};
      reg_RW0_addr = {1 {$random}};
    end
  `endif
  integer i;
  always @(posedge RW0_clk)
    reg_RW0_ren <= RW0_en && !RW0_wmode;
  always @(posedge RW0_clk)
    if (RW0_en && !RW0_wmode) reg_RW0_addr <= RW0_addr;
  always @(posedge RW0_clk)
    if (RW0_en && RW0_wmode) begin
      for(i=0;i<4;i=i+1) begin
        if(RW0_wmask[i]) begin
          ram[RW0_addr][i*24 +: 24] <= RW0_wdata[i*24 +: 24];
        end
      end
    end
  `ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [95:0] RW0_random;
  `ifdef RANDOMIZE_MEM_INIT
    initial begin
      #`RANDOMIZE_DELAY begin end
      RW0_random = {$random, $random, $random};
      reg_RW0_ren = RW0_random[0];
    end
  `endif
  always @(posedge RW0_clk) RW0_random <= {$random, $random, $random};
  assign RW0_rdata = reg_RW0_ren ? ram[reg_RW0_addr] : RW0_random[95:0];
  `else
  assign RW0_rdata = ram[reg_RW0_addr];
  `endif

endmodule
