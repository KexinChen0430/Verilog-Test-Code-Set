module page352;

`define first_half "start of string
$display(`first_half end of string");

`define max(a,b)((a) > (b) ? (a) : (b))
n = `max(p+q, r+s) ;

endmodule