module constmod ;

input

a1=8'b10101100,  //λ��Ϊ8�����Ķ����Ʊ�ʾ, 'b��ʾ������
a2=8'ha2,        //λ��Ϊ8������ʮ�����ƣ�'h��ʾʮ�����ơ�

b1=4'b10x0, //λ��Ϊ4�Ķ��������ӵ�λ����ڶ�λΪ����ֵ
b2=4'b101z, //λ��Ϊ4�Ķ��������ӵ�λ�����һλΪ����ֵ
b3=12'dz,   //λ��Ϊ12��ʮ��������ֵΪ����ֵ(��һ�ֱ�﷽ʽ)
b4=12'd?,   //λ��Ϊ12��ʮ��������ֵΪ����ֵ(�ڶ��ֱ�﷽ʽ)
b5=8'h4x,   //λ��Ϊ8��ʮ�������������λֵΪ����ֵ

c1=-8'd5,   //������ʽ����5�Ĳ������ð�λ����������ʾ)
c2=16'b1010_1011_1111_1010,
c3=1,
c4=-1,
c5='BX
;

parameter  msb=7;       //�������msbΪ����7
parameter  e=25, f=29;  //��������������� 
parameter  r=5.7;       //����rΪһ��ʵ�Ͳ��� 
parameter  byte_size=8, byte_msb=byte_size-1; //�ó������ʽ��ֵ 
parameter  average_delay = (r+f)/2;           //�ó������ʽ��ֵ 

endmodule