`define xxx a^b
module aaa(a,b,out);
input a, b;
output `out;
`define yyy out =
wire out;
assign  `yyy `xxx;
endmodule 