module XbarCircuit_2(
  input          clock,
  input          reset,
  output         io_in_1_a_ready,
  input          io_in_1_a_valid,
  input  [2:0]   io_in_1_a_bits_opcode,
  input  [2:0]   io_in_1_a_bits_size,
  input  [5:0]   io_in_1_a_bits_source,
  input  [35:0]  io_in_1_a_bits_address,
  input  [31:0]  io_in_1_a_bits_mask,
  input  [255:0] io_in_1_a_bits_data,
  input          io_in_1_d_ready,
  output         io_in_1_d_valid,
  output [2:0]   io_in_1_d_bits_opcode,
  output [1:0]   io_in_1_d_bits_param,
  output [2:0]   io_in_1_d_bits_size,
  output [5:0]   io_in_1_d_bits_source,
  output         io_in_1_d_bits_denied,
  output [255:0] io_in_1_d_bits_data,
  output         io_in_0_a_ready,
  input          io_in_0_a_valid,
  input  [2:0]   io_in_0_a_bits_opcode,
  input  [2:0]   io_in_0_a_bits_size,
  input  [5:0]   io_in_0_a_bits_source,
  input  [35:0]  io_in_0_a_bits_address,
  input  [31:0]  io_in_0_a_bits_mask,
  input  [255:0] io_in_0_a_bits_data,
  input          io_in_0_d_ready,
  output         io_in_0_d_valid,
  output [2:0]   io_in_0_d_bits_opcode,
  output [1:0]   io_in_0_d_bits_param,
  output [2:0]   io_in_0_d_bits_size,
  output [5:0]   io_in_0_d_bits_source,
  output         io_in_0_d_bits_denied,
  output [255:0] io_in_0_d_bits_data,
  input          io_out_0_a_ready,
  output         io_out_0_a_valid,
  output [2:0]   io_out_0_a_bits_opcode,
  output [2:0]   io_out_0_a_bits_size,
  output [6:0]   io_out_0_a_bits_source,
  output [35:0]  io_out_0_a_bits_address,
  output [31:0]  io_out_0_a_bits_mask,
  output [255:0] io_out_0_a_bits_data,
  output         io_out_0_d_ready,
  input          io_out_0_d_valid,
  input  [2:0]   io_out_0_d_bits_opcode,
  input  [1:0]   io_out_0_d_bits_param,
  input  [2:0]   io_out_0_d_bits_size,
  input  [6:0]   io_out_0_d_bits_source,
  input          io_out_0_d_bits_denied,
  input  [255:0] io_out_0_d_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] _GEN_1 = {{1'd0}, io_in_0_a_bits_source}; // @[Xbar.scala 237:55]
  wire [6:0] _T = _GEN_1 | 7'h40; // @[Xbar.scala 237:55]
  wire  _T_56 = ~io_out_0_d_bits_source[6]; // @[Parameters.scala 54:32]
  wire [12:0] _T_62 = 13'h3f << io_in_0_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _T_64 = ~_T_62[5:0]; // @[package.scala 234:46]
  wire  _T_67 = ~io_in_0_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire  _T_68 = _T_67 & _T_64[5]; // @[Edges.scala 220:14]
  wire [12:0] _T_70 = 13'h3f << io_in_1_a_bits_size; // @[package.scala 234:77]
  wire [5:0] _T_72 = ~_T_70[5:0]; // @[package.scala 234:46]
  wire  _T_75 = ~io_in_1_a_bits_opcode[2]; // @[Edges.scala 91:28]
  wire  _T_76 = _T_75 & _T_72[5]; // @[Edges.scala 220:14]
  reg  REG; // @[Arbiter.scala 87:30]
  wire  _T_132 = ~REG; // @[Arbiter.scala 88:28]
  wire  _T_133 = _T_132 & io_out_0_a_ready; // @[Arbiter.scala 89:24]
  wire [1:0] _T_138 = {io_in_1_a_valid,io_in_0_a_valid}; // @[Cat.scala 30:58]
  reg [1:0] REG_1; // @[Arbiter.scala 23:23]
  wire [1:0] _T_144 = ~REG_1; // @[Arbiter.scala 24:30]
  wire [1:0] _T_145 = _T_138 & _T_144; // @[Arbiter.scala 24:28]
  wire [3:0] _T_146 = {_T_145,io_in_1_a_valid,io_in_0_a_valid}; // @[Cat.scala 30:58]
  wire [3:0] _GEN_2 = {{1'd0}, _T_146[3:1]}; // @[package.scala 253:43]
  wire [3:0] _T_148 = _T_146 | _GEN_2; // @[package.scala 253:43]
  wire [3:0] _T_151 = {REG_1, 2'h0}; // @[Arbiter.scala 25:66]
  wire [3:0] _GEN_3 = {{1'd0}, _T_148[3:1]}; // @[Arbiter.scala 25:58]
  wire [3:0] _T_152 = _GEN_3 | _T_151; // @[Arbiter.scala 25:58]
  wire [1:0] _T_155 = _T_152[3:2] & _T_152[1:0]; // @[Arbiter.scala 26:39]
  wire [1:0] _T_156 = ~_T_155; // @[Arbiter.scala 26:18]
  wire [1:0] _T_159 = _T_156 & _T_138; // @[Arbiter.scala 28:29]
  wire [2:0] _T_160 = {_T_159, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _T_162 = _T_159 | _T_160[1:0]; // @[package.scala 244:43]
  wire  _T_167 = _T_156[0] & io_in_0_a_valid; // @[Arbiter.scala 97:79]
  wire  _T_168 = _T_156[1] & io_in_1_a_valid; // @[Arbiter.scala 97:79]
  wire  _T_183 = io_in_0_a_valid | io_in_1_a_valid; // @[Arbiter.scala 107:36]
  wire  _T_197 = _T_167 & _T_68; // @[Arbiter.scala 111:73]
  wire  _T_198 = _T_168 & _T_76; // @[Arbiter.scala 111:73]
  wire  _T_199 = _T_197 | _T_198; // @[Arbiter.scala 112:44]
  reg  REG_2_0; // @[Arbiter.scala 116:26]
  wire  _T_206_0 = _T_132 ? _T_167 : REG_2_0; // @[Arbiter.scala 117:30]
  reg  REG_2_1; // @[Arbiter.scala 116:26]
  wire  _T_206_1 = _T_132 ? _T_168 : REG_2_1; // @[Arbiter.scala 117:30]
  wire  _T_214 = REG_2_0 & io_in_0_a_valid | REG_2_1 & io_in_1_a_valid; // @[Mux.scala 27:72]
  wire  _T_215 = _T_132 ? _T_183 : _T_214; // @[Arbiter.scala 125:29]
  wire  _T_202 = io_out_0_a_ready & _T_215; // @[ReadyValidCancel.scala 50:33]
  wire  _T_208_0 = _T_132 ? _T_156[0] : REG_2_0; // @[Arbiter.scala 121:24]
  wire  _T_208_1 = _T_132 ? _T_156[1] : REG_2_1; // @[Arbiter.scala 121:24]
  wire [255:0] _T_222 = _T_206_0 ? io_in_0_a_bits_data : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_223 = _T_206_1 ? io_in_1_a_bits_data : 256'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_225 = _T_206_0 ? io_in_0_a_bits_mask : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_226 = _T_206_1 ? io_in_1_a_bits_mask : 32'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_228 = _T_206_0 ? io_in_0_a_bits_address : 36'h0; // @[Mux.scala 27:72]
  wire [35:0] _T_229 = _T_206_1 ? io_in_1_a_bits_address : 36'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_231 = _T_206_0 ? _T : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _WIRE_9_1_a_bits_source = {{1'd0}, io_in_1_a_bits_source}; // @[Xbar.scala 231:18 237:29]
  wire [6:0] _T_232 = _T_206_1 ? _WIRE_9_1_a_bits_source : 7'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_234 = _T_206_0 ? io_in_0_a_bits_size : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_235 = _T_206_1 ? io_in_1_a_bits_size : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_240 = _T_206_0 ? io_in_0_a_bits_opcode : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_241 = _T_206_1 ? io_in_1_a_bits_opcode : 3'h0; // @[Mux.scala 27:72]
  assign io_in_1_a_ready = io_out_0_a_ready & _T_208_1; // @[Arbiter.scala 123:31]
  assign io_in_1_d_valid = io_out_0_d_valid & _T_56; // @[Xbar.scala 179:40]
  assign io_in_1_d_bits_opcode = io_out_0_d_bits_opcode; // @[Bundle_ACancel.scala 23:19 Xbar.scala 136:12]
  assign io_in_1_d_bits_param = io_out_0_d_bits_param; // @[Bundle_ACancel.scala 23:19 Xbar.scala 136:12]
  assign io_in_1_d_bits_size = io_out_0_d_bits_size; // @[Bundle_ACancel.scala 23:19 Xbar.scala 136:12]
  assign io_in_1_d_bits_source = io_out_0_d_bits_source[5:0]; // @[Xbar.scala 228:69]
  assign io_in_1_d_bits_denied = io_out_0_d_bits_denied; // @[Bundle_ACancel.scala 23:19 Xbar.scala 136:12]
  assign io_in_1_d_bits_data = io_out_0_d_bits_data; // @[Bundle_ACancel.scala 23:19 Xbar.scala 136:12]
  assign io_in_0_a_ready = io_out_0_a_ready & _T_208_0; // @[Arbiter.scala 123:31]
  assign io_in_0_d_valid = io_out_0_d_valid & io_out_0_d_bits_source[6]; // @[Xbar.scala 179:40]
  assign io_in_0_d_bits_opcode = io_out_0_d_bits_opcode; // @[Bundle_ACancel.scala 23:19 Xbar.scala 136:12]
  assign io_in_0_d_bits_param = io_out_0_d_bits_param; // @[Bundle_ACancel.scala 23:19 Xbar.scala 136:12]
  assign io_in_0_d_bits_size = io_out_0_d_bits_size; // @[Bundle_ACancel.scala 23:19 Xbar.scala 136:12]
  assign io_in_0_d_bits_source = io_out_0_d_bits_source[5:0]; // @[Xbar.scala 228:69]
  assign io_in_0_d_bits_denied = io_out_0_d_bits_denied; // @[Bundle_ACancel.scala 23:19 Xbar.scala 136:12]
  assign io_in_0_d_bits_data = io_out_0_d_bits_data; // @[Bundle_ACancel.scala 23:19 Xbar.scala 136:12]
  assign io_out_0_a_valid = _T_132 ? _T_183 : _T_214; // @[Arbiter.scala 125:29]
  assign io_out_0_a_bits_opcode = _T_240 | _T_241; // @[Mux.scala 27:72]
  assign io_out_0_a_bits_size = _T_234 | _T_235; // @[Mux.scala 27:72]
  assign io_out_0_a_bits_source = _T_231 | _T_232; // @[Mux.scala 27:72]
  assign io_out_0_a_bits_address = _T_228 | _T_229; // @[Mux.scala 27:72]
  assign io_out_0_a_bits_mask = _T_225 | _T_226; // @[Mux.scala 27:72]
  assign io_out_0_a_bits_data = _T_222 | _T_223; // @[Mux.scala 27:72]
  assign io_out_0_d_ready = io_out_0_d_bits_source[6] & io_in_0_d_ready | _T_56 & io_in_1_d_ready; // @[Mux.scala 27:72]
  always @(posedge clock) begin
    if (reset) begin // @[Arbiter.scala 87:30]
      REG <= 1'h0; // @[Arbiter.scala 87:30]
    end else if (_T_133) begin // @[Arbiter.scala 113:23]
      REG <= _T_199;
    end else begin
      REG <= REG - _T_202;
    end
    if (reset) begin // @[Arbiter.scala 23:23]
      REG_1 <= 2'h3; // @[Arbiter.scala 23:23]
    end else if (_T_133 & |_T_138) begin // @[Arbiter.scala 27:32]
      REG_1 <= _T_162; // @[Arbiter.scala 28:12]
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      REG_2_0 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (_T_132) begin // @[Arbiter.scala 117:30]
      REG_2_0 <= _T_167;
    end
    if (reset) begin // @[Arbiter.scala 116:26]
      REG_2_1 <= 1'h0; // @[Arbiter.scala 116:26]
    end else if (_T_132) begin // @[Arbiter.scala 117:30]
      REG_2_1 <= _T_168;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  REG_2_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  REG_2_1 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule