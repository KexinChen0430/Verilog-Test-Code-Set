// module add(x, y ,out);
//   input [1:0] x;
//   input [1:0] y;
//   output [1:0] out;

//   assign out = x + y;

// endmodule

module add(x, y ,out);
  input x;
  input y;
  output out;

  assign out = x + y;

endmodule