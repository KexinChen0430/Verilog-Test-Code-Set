
`timescale 1ns/1ns 
 
module t; 
 
reg a = 1;

reg [7:0]      data_buf[8:0];

endmodule