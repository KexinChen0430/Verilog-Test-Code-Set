module ysyx_210128_PatternHistoryTableLocal(
  input        clock,
  input        reset,
  input  [2:0] io_rindex_0,
  input  [2:0] io_rindex_1,
  input  [5:0] io_raddr_0,
  input  [5:0] io_raddr_1,
  output       io_rdirect_0,
  output       io_rdirect_1,
  input  [2:0] io_windex,
  input  [5:0] io_waddr,
  input        io_wen,
  input        io_wjmp
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_77;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
`endif // RANDOMIZE_REG_INIT
  reg  pht_1_0 [0:63]; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_0_MPORT_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_0_MPORT_8_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_8_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_8_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_0_MPORT_16_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_16_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_16_data; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_32_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_32_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_32_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_32_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_48_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_48_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_48_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_48_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_50_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_50_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_50_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_50_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_52_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_52_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_52_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_52_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_54_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_54_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_54_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_54_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_56_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_56_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_56_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_56_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_58_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_58_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_58_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_58_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_60_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_60_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_60_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_60_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_62_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_62_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_62_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_62_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_64_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_64_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_64_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_64_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_66_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_66_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_66_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_66_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_68_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_68_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_68_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_68_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_70_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_70_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_70_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_70_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_72_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_72_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_72_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_72_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_74_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_74_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_74_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_74_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_76_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_76_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_76_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_76_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_78_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_78_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_78_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_78_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_80_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_80_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_80_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_80_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_82_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_82_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_82_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_82_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_84_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_84_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_84_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_84_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_86_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_86_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_86_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_86_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_88_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_88_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_88_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_88_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_90_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_90_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_90_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_90_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_92_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_92_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_92_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_92_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_94_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_94_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_94_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_94_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_96_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_96_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_96_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_96_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_98_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_98_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_98_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_98_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_100_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_100_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_100_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_100_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_102_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_102_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_102_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_102_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_104_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_104_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_104_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_104_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_106_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_106_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_106_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_106_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_108_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_108_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_108_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_108_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_110_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_110_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_110_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_110_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_112_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_112_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_112_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_112_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_114_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_114_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_114_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_114_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_116_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_116_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_116_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_116_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_118_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_118_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_118_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_118_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_120_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_120_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_120_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_120_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_122_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_122_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_122_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_122_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_124_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_124_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_124_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_124_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_126_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_126_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_126_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_126_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_128_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_128_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_128_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_128_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_130_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_130_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_130_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_130_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_132_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_132_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_132_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_132_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_134_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_134_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_134_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_134_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_136_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_136_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_136_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_136_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_138_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_138_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_138_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_138_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_140_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_140_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_140_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_140_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_142_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_142_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_142_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_142_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_144_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_144_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_144_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_144_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_146_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_146_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_146_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_146_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_148_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_148_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_148_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_148_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_150_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_150_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_150_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_150_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_152_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_152_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_152_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_152_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_154_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_154_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_154_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_154_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_156_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_156_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_156_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_156_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_158_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_158_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_158_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_158_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_160_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_160_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_160_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_160_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_162_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_162_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_162_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_162_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_164_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_164_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_164_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_164_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_166_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_166_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_166_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_166_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_168_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_168_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_168_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_168_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_170_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_170_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_170_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_170_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_172_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_172_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_172_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_172_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_174_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_0_MPORT_174_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_174_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_0_MPORT_174_en; // @[PatternHistoryTable.scala 21:28]
//   reg  pht_1_0_MPORT_en_pipe_0;
  reg [5:0] pht_1_0_MPORT_addr_pipe_0;
//   reg  pht_1_0_MPORT_8_en_pipe_0;
  reg [5:0] pht_1_0_MPORT_8_addr_pipe_0;
//   reg  pht_1_0_MPORT_16_en_pipe_0;
  reg [5:0] pht_1_0_MPORT_16_addr_pipe_0;
  reg  pht_1_1 [0:63]; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_1_MPORT_1_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_1_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_1_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_1_MPORT_9_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_9_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_9_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_1_MPORT_18_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_18_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_18_data; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_34_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_34_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_34_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_34_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_176_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_176_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_176_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_176_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_178_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_178_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_178_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_178_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_180_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_180_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_180_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_180_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_182_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_182_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_182_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_182_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_184_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_184_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_184_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_184_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_186_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_186_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_186_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_186_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_188_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_188_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_188_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_188_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_190_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_190_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_190_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_190_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_192_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_192_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_192_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_192_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_194_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_194_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_194_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_194_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_196_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_196_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_196_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_196_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_198_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_198_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_198_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_198_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_200_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_200_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_200_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_200_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_202_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_202_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_202_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_202_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_204_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_204_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_204_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_204_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_206_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_206_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_206_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_206_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_208_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_208_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_208_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_208_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_210_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_210_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_210_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_210_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_212_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_212_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_212_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_212_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_214_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_214_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_214_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_214_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_216_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_216_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_216_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_216_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_218_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_218_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_218_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_218_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_220_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_220_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_220_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_220_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_222_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_222_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_222_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_222_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_224_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_224_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_224_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_224_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_226_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_226_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_226_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_226_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_228_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_228_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_228_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_228_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_230_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_230_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_230_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_230_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_232_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_232_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_232_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_232_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_234_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_234_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_234_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_234_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_236_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_236_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_236_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_236_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_238_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_238_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_238_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_238_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_240_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_240_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_240_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_240_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_242_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_242_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_242_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_242_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_244_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_244_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_244_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_244_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_246_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_246_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_246_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_246_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_248_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_248_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_248_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_248_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_250_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_250_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_250_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_250_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_252_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_252_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_252_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_252_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_254_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_254_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_254_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_254_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_256_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_256_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_256_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_256_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_258_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_258_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_258_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_258_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_260_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_260_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_260_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_260_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_262_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_262_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_262_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_262_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_264_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_264_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_264_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_264_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_266_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_266_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_266_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_266_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_268_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_268_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_268_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_268_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_270_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_270_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_270_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_270_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_272_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_272_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_272_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_272_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_274_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_274_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_274_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_274_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_276_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_276_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_276_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_276_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_278_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_278_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_278_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_278_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_280_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_280_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_280_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_280_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_282_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_282_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_282_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_282_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_284_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_284_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_284_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_284_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_286_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_286_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_286_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_286_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_288_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_288_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_288_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_288_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_290_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_290_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_290_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_290_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_292_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_292_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_292_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_292_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_294_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_294_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_294_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_294_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_296_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_296_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_296_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_296_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_298_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_298_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_298_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_298_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_300_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_300_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_300_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_300_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_302_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_1_MPORT_302_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_302_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_1_MPORT_302_en; // @[PatternHistoryTable.scala 21:28]
//   reg  pht_1_1_MPORT_1_en_pipe_0;
  reg [5:0] pht_1_1_MPORT_1_addr_pipe_0;
//   reg  pht_1_1_MPORT_9_en_pipe_0;
  reg [5:0] pht_1_1_MPORT_9_addr_pipe_0;
//   reg  pht_1_1_MPORT_18_en_pipe_0;
  reg [5:0] pht_1_1_MPORT_18_addr_pipe_0;
  reg  pht_1_2 [0:63]; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_2_MPORT_2_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_2_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_2_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_2_MPORT_10_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_10_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_10_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_2_MPORT_20_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_20_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_20_data; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_36_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_36_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_36_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_36_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_304_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_304_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_304_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_304_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_306_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_306_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_306_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_306_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_308_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_308_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_308_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_308_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_310_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_310_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_310_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_310_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_312_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_312_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_312_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_312_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_314_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_314_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_314_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_314_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_316_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_316_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_316_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_316_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_318_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_318_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_318_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_318_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_320_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_320_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_320_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_320_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_322_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_322_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_322_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_322_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_324_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_324_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_324_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_324_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_326_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_326_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_326_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_326_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_328_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_328_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_328_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_328_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_330_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_330_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_330_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_330_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_332_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_332_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_332_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_332_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_334_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_334_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_334_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_334_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_336_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_336_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_336_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_336_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_338_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_338_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_338_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_338_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_340_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_340_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_340_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_340_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_342_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_342_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_342_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_342_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_344_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_344_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_344_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_344_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_346_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_346_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_346_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_346_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_348_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_348_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_348_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_348_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_350_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_350_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_350_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_350_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_352_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_352_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_352_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_352_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_354_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_354_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_354_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_354_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_356_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_356_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_356_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_356_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_358_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_358_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_358_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_358_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_360_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_360_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_360_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_360_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_362_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_362_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_362_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_362_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_364_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_364_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_364_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_364_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_366_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_366_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_366_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_366_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_368_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_368_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_368_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_368_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_370_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_370_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_370_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_370_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_372_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_372_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_372_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_372_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_374_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_374_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_374_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_374_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_376_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_376_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_376_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_376_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_378_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_378_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_378_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_378_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_380_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_380_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_380_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_380_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_382_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_382_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_382_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_382_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_384_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_384_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_384_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_384_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_386_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_386_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_386_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_386_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_388_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_388_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_388_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_388_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_390_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_390_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_390_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_390_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_392_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_392_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_392_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_392_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_394_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_394_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_394_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_394_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_396_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_396_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_396_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_396_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_398_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_398_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_398_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_398_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_400_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_400_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_400_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_400_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_402_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_402_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_402_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_402_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_404_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_404_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_404_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_404_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_406_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_406_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_406_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_406_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_408_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_408_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_408_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_408_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_410_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_410_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_410_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_410_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_412_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_412_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_412_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_412_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_414_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_414_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_414_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_414_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_416_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_416_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_416_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_416_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_418_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_418_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_418_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_418_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_420_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_420_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_420_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_420_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_422_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_422_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_422_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_422_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_424_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_424_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_424_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_424_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_426_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_426_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_426_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_426_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_428_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_428_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_428_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_428_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_430_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_2_MPORT_430_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_430_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_2_MPORT_430_en; // @[PatternHistoryTable.scala 21:28]
//   reg  pht_1_2_MPORT_2_en_pipe_0;
  reg [5:0] pht_1_2_MPORT_2_addr_pipe_0;
//   reg  pht_1_2_MPORT_10_en_pipe_0;
  reg [5:0] pht_1_2_MPORT_10_addr_pipe_0;
//   reg  pht_1_2_MPORT_20_en_pipe_0;
  reg [5:0] pht_1_2_MPORT_20_addr_pipe_0;
  reg  pht_1_3 [0:63]; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_3_MPORT_3_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_3_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_3_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_3_MPORT_11_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_11_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_11_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_3_MPORT_22_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_22_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_22_data; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_38_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_38_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_38_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_38_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_432_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_432_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_432_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_432_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_434_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_434_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_434_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_434_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_436_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_436_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_436_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_436_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_438_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_438_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_438_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_438_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_440_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_440_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_440_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_440_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_442_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_442_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_442_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_442_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_444_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_444_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_444_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_444_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_446_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_446_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_446_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_446_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_448_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_448_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_448_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_448_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_450_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_450_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_450_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_450_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_452_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_452_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_452_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_452_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_454_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_454_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_454_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_454_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_456_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_456_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_456_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_456_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_458_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_458_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_458_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_458_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_460_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_460_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_460_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_460_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_462_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_462_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_462_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_462_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_464_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_464_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_464_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_464_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_466_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_466_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_466_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_466_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_468_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_468_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_468_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_468_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_470_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_470_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_470_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_470_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_472_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_472_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_472_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_472_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_474_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_474_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_474_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_474_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_476_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_476_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_476_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_476_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_478_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_478_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_478_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_478_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_480_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_480_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_480_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_480_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_482_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_482_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_482_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_482_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_484_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_484_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_484_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_484_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_486_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_486_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_486_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_486_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_488_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_488_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_488_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_488_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_490_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_490_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_490_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_490_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_492_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_492_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_492_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_492_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_494_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_494_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_494_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_494_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_496_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_496_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_496_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_496_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_498_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_498_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_498_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_498_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_500_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_500_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_500_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_500_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_502_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_502_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_502_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_502_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_504_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_504_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_504_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_504_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_506_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_506_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_506_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_506_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_508_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_508_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_508_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_508_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_510_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_510_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_510_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_510_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_512_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_512_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_512_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_512_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_514_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_514_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_514_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_514_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_516_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_516_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_516_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_516_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_518_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_518_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_518_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_518_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_520_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_520_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_520_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_520_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_522_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_522_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_522_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_522_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_524_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_524_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_524_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_524_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_526_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_526_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_526_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_526_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_528_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_528_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_528_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_528_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_530_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_530_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_530_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_530_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_532_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_532_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_532_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_532_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_534_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_534_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_534_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_534_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_536_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_536_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_536_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_536_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_538_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_538_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_538_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_538_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_540_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_540_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_540_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_540_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_542_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_542_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_542_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_542_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_544_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_544_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_544_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_544_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_546_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_546_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_546_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_546_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_548_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_548_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_548_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_548_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_550_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_550_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_550_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_550_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_552_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_552_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_552_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_552_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_554_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_554_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_554_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_554_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_556_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_556_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_556_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_556_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_558_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_3_MPORT_558_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_558_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_3_MPORT_558_en; // @[PatternHistoryTable.scala 21:28]
//   reg  pht_1_3_MPORT_3_en_pipe_0;
  reg [5:0] pht_1_3_MPORT_3_addr_pipe_0;
//   reg  pht_1_3_MPORT_11_en_pipe_0;
  reg [5:0] pht_1_3_MPORT_11_addr_pipe_0;
//   reg  pht_1_3_MPORT_22_en_pipe_0;
  reg [5:0] pht_1_3_MPORT_22_addr_pipe_0;
  reg  pht_1_4 [0:63]; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_4_MPORT_4_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_4_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_4_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_4_MPORT_12_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_12_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_12_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_4_MPORT_24_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_24_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_24_data; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_40_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_40_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_40_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_40_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_560_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_560_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_560_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_560_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_562_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_562_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_562_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_562_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_564_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_564_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_564_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_564_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_566_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_566_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_566_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_566_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_568_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_568_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_568_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_568_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_570_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_570_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_570_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_570_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_572_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_572_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_572_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_572_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_574_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_574_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_574_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_574_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_576_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_576_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_576_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_576_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_578_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_578_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_578_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_578_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_580_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_580_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_580_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_580_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_582_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_582_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_582_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_582_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_584_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_584_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_584_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_584_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_586_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_586_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_586_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_586_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_588_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_588_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_588_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_588_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_590_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_590_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_590_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_590_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_592_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_592_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_592_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_592_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_594_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_594_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_594_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_594_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_596_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_596_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_596_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_596_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_598_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_598_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_598_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_598_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_600_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_600_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_600_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_600_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_602_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_602_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_602_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_602_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_604_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_604_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_604_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_604_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_606_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_606_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_606_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_606_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_608_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_608_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_608_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_608_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_610_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_610_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_610_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_610_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_612_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_612_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_612_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_612_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_614_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_614_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_614_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_614_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_616_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_616_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_616_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_616_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_618_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_618_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_618_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_618_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_620_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_620_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_620_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_620_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_622_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_622_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_622_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_622_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_624_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_624_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_624_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_624_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_626_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_626_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_626_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_626_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_628_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_628_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_628_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_628_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_630_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_630_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_630_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_630_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_632_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_632_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_632_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_632_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_634_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_634_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_634_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_634_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_636_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_636_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_636_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_636_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_638_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_638_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_638_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_638_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_640_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_640_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_640_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_640_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_642_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_642_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_642_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_642_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_644_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_644_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_644_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_644_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_646_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_646_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_646_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_646_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_648_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_648_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_648_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_648_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_650_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_650_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_650_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_650_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_652_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_652_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_652_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_652_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_654_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_654_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_654_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_654_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_656_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_656_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_656_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_656_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_658_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_658_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_658_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_658_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_660_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_660_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_660_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_660_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_662_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_662_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_662_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_662_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_664_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_664_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_664_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_664_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_666_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_666_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_666_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_666_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_668_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_668_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_668_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_668_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_670_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_670_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_670_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_670_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_672_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_672_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_672_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_672_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_674_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_674_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_674_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_674_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_676_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_676_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_676_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_676_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_678_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_678_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_678_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_678_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_680_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_680_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_680_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_680_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_682_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_682_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_682_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_682_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_684_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_684_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_684_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_684_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_686_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_4_MPORT_686_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_686_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_4_MPORT_686_en; // @[PatternHistoryTable.scala 21:28]
//   reg  pht_1_4_MPORT_4_en_pipe_0;
  reg [5:0] pht_1_4_MPORT_4_addr_pipe_0;
//   reg  pht_1_4_MPORT_12_en_pipe_0;
  reg [5:0] pht_1_4_MPORT_12_addr_pipe_0;
//   reg  pht_1_4_MPORT_24_en_pipe_0;
  reg [5:0] pht_1_4_MPORT_24_addr_pipe_0;
  reg  pht_1_5 [0:63]; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_5_MPORT_5_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_5_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_5_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_5_MPORT_13_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_13_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_13_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_5_MPORT_26_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_26_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_26_data; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_42_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_42_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_42_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_42_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_688_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_688_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_688_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_688_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_690_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_690_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_690_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_690_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_692_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_692_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_692_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_692_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_694_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_694_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_694_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_694_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_696_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_696_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_696_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_696_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_698_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_698_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_698_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_698_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_700_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_700_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_700_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_700_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_702_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_702_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_702_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_702_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_704_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_704_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_704_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_704_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_706_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_706_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_706_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_706_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_708_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_708_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_708_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_708_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_710_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_710_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_710_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_710_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_712_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_712_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_712_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_712_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_714_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_714_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_714_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_714_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_716_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_716_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_716_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_716_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_718_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_718_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_718_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_718_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_720_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_720_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_720_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_720_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_722_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_722_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_722_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_722_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_724_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_724_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_724_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_724_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_726_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_726_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_726_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_726_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_728_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_728_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_728_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_728_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_730_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_730_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_730_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_730_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_732_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_732_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_732_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_732_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_734_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_734_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_734_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_734_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_736_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_736_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_736_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_736_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_738_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_738_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_738_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_738_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_740_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_740_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_740_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_740_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_742_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_742_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_742_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_742_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_744_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_744_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_744_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_744_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_746_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_746_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_746_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_746_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_748_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_748_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_748_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_748_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_750_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_750_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_750_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_750_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_752_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_752_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_752_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_752_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_754_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_754_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_754_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_754_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_756_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_756_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_756_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_756_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_758_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_758_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_758_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_758_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_760_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_760_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_760_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_760_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_762_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_762_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_762_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_762_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_764_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_764_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_764_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_764_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_766_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_766_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_766_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_766_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_768_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_768_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_768_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_768_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_770_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_770_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_770_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_770_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_772_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_772_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_772_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_772_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_774_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_774_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_774_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_774_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_776_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_776_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_776_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_776_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_778_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_778_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_778_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_778_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_780_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_780_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_780_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_780_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_782_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_782_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_782_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_782_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_784_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_784_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_784_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_784_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_786_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_786_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_786_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_786_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_788_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_788_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_788_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_788_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_790_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_790_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_790_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_790_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_792_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_792_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_792_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_792_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_794_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_794_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_794_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_794_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_796_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_796_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_796_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_796_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_798_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_798_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_798_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_798_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_800_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_800_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_800_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_800_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_802_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_802_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_802_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_802_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_804_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_804_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_804_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_804_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_806_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_806_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_806_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_806_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_808_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_808_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_808_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_808_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_810_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_810_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_810_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_810_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_812_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_812_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_812_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_812_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_814_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_5_MPORT_814_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_814_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_5_MPORT_814_en; // @[PatternHistoryTable.scala 21:28]
//   reg  pht_1_5_MPORT_5_en_pipe_0;
  reg [5:0] pht_1_5_MPORT_5_addr_pipe_0;
//   reg  pht_1_5_MPORT_13_en_pipe_0;
  reg [5:0] pht_1_5_MPORT_13_addr_pipe_0;
//   reg  pht_1_5_MPORT_26_en_pipe_0;
  reg [5:0] pht_1_5_MPORT_26_addr_pipe_0;
  reg  pht_1_6 [0:63]; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_6_MPORT_6_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_6_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_6_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_6_MPORT_14_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_14_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_14_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_6_MPORT_28_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_28_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_28_data; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_44_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_44_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_44_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_44_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_816_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_816_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_816_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_816_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_818_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_818_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_818_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_818_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_820_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_820_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_820_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_820_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_822_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_822_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_822_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_822_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_824_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_824_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_824_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_824_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_826_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_826_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_826_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_826_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_828_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_828_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_828_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_828_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_830_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_830_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_830_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_830_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_832_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_832_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_832_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_832_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_834_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_834_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_834_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_834_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_836_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_836_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_836_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_836_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_838_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_838_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_838_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_838_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_840_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_840_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_840_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_840_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_842_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_842_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_842_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_842_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_844_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_844_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_844_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_844_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_846_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_846_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_846_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_846_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_848_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_848_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_848_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_848_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_850_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_850_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_850_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_850_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_852_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_852_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_852_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_852_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_854_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_854_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_854_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_854_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_856_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_856_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_856_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_856_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_858_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_858_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_858_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_858_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_860_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_860_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_860_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_860_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_862_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_862_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_862_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_862_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_864_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_864_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_864_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_864_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_866_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_866_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_866_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_866_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_868_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_868_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_868_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_868_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_870_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_870_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_870_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_870_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_872_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_872_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_872_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_872_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_874_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_874_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_874_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_874_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_876_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_876_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_876_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_876_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_878_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_878_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_878_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_878_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_880_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_880_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_880_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_880_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_882_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_882_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_882_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_882_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_884_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_884_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_884_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_884_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_886_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_886_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_886_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_886_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_888_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_888_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_888_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_888_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_890_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_890_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_890_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_890_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_892_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_892_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_892_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_892_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_894_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_894_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_894_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_894_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_896_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_896_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_896_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_896_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_898_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_898_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_898_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_898_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_900_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_900_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_900_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_900_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_902_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_902_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_902_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_902_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_904_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_904_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_904_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_904_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_906_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_906_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_906_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_906_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_908_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_908_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_908_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_908_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_910_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_910_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_910_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_910_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_912_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_912_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_912_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_912_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_914_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_914_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_914_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_914_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_916_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_916_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_916_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_916_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_918_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_918_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_918_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_918_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_920_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_920_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_920_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_920_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_922_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_922_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_922_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_922_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_924_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_924_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_924_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_924_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_926_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_926_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_926_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_926_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_928_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_928_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_928_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_928_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_930_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_930_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_930_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_930_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_932_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_932_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_932_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_932_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_934_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_934_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_934_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_934_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_936_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_936_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_936_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_936_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_938_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_938_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_938_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_938_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_940_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_940_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_940_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_940_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_942_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_6_MPORT_942_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_942_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_6_MPORT_942_en; // @[PatternHistoryTable.scala 21:28]
//   reg  pht_1_6_MPORT_6_en_pipe_0;
  reg [5:0] pht_1_6_MPORT_6_addr_pipe_0;
//   reg  pht_1_6_MPORT_14_en_pipe_0;
  reg [5:0] pht_1_6_MPORT_14_addr_pipe_0;
//   reg  pht_1_6_MPORT_28_en_pipe_0;
  reg [5:0] pht_1_6_MPORT_28_addr_pipe_0;
  reg  pht_1_7 [0:63]; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_7_MPORT_7_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_7_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_7_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_7_MPORT_15_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_15_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_15_data; // @[PatternHistoryTable.scala 21:28]
//   wire  pht_1_7_MPORT_30_en; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_30_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_30_data; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_46_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_46_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_46_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_46_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_944_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_944_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_944_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_944_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_946_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_946_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_946_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_946_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_948_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_948_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_948_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_948_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_950_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_950_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_950_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_950_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_952_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_952_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_952_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_952_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_954_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_954_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_954_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_954_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_956_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_956_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_956_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_956_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_958_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_958_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_958_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_958_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_960_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_960_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_960_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_960_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_962_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_962_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_962_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_962_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_964_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_964_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_964_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_964_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_966_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_966_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_966_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_966_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_968_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_968_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_968_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_968_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_970_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_970_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_970_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_970_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_972_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_972_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_972_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_972_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_974_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_974_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_974_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_974_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_976_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_976_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_976_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_976_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_978_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_978_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_978_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_978_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_980_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_980_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_980_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_980_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_982_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_982_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_982_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_982_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_984_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_984_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_984_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_984_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_986_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_986_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_986_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_986_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_988_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_988_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_988_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_988_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_990_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_990_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_990_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_990_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_992_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_992_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_992_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_992_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_994_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_994_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_994_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_994_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_996_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_996_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_996_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_996_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_998_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_998_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_998_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_998_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1000_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1000_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1000_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1000_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1002_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1002_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1002_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1002_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1004_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1004_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1004_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1004_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1006_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1006_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1006_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1006_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1008_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1008_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1008_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1008_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1010_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1010_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1010_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1010_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1012_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1012_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1012_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1012_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1014_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1014_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1014_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1014_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1016_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1016_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1016_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1016_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1018_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1018_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1018_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1018_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1020_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1020_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1020_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1020_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1022_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1022_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1022_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1022_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1024_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1024_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1024_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1024_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1026_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1026_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1026_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1026_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1028_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1028_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1028_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1028_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1030_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1030_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1030_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1030_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1032_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1032_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1032_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1032_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1034_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1034_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1034_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1034_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1036_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1036_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1036_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1036_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1038_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1038_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1038_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1038_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1040_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1040_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1040_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1040_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1042_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1042_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1042_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1042_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1044_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1044_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1044_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1044_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1046_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1046_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1046_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1046_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1048_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1048_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1048_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1048_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1050_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1050_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1050_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1050_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1052_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1052_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1052_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1052_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1054_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1054_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1054_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1054_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1056_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1056_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1056_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1056_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1058_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1058_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1058_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1058_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1060_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1060_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1060_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1060_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1062_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1062_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1062_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1062_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1064_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1064_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1064_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1064_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1066_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1066_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1066_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1066_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1068_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1068_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1068_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1068_en; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1070_data; // @[PatternHistoryTable.scala 21:28]
  wire [5:0] pht_1_7_MPORT_1070_addr; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1070_mask; // @[PatternHistoryTable.scala 21:28]
  wire  pht_1_7_MPORT_1070_en; // @[PatternHistoryTable.scala 21:28]
//   reg  pht_1_7_MPORT_7_en_pipe_0;
  reg [5:0] pht_1_7_MPORT_7_addr_pipe_0;
//   reg  pht_1_7_MPORT_15_en_pipe_0;
  reg [5:0] pht_1_7_MPORT_15_addr_pipe_0;
//   reg  pht_1_7_MPORT_30_en_pipe_0;
  reg [5:0] pht_1_7_MPORT_30_addr_pipe_0;
  reg  pht_0_0 [0:63]; // @[PatternHistoryTable.scala 26:28]
//   wire  pht_0_0_MPORT_17_en; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_17_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_17_data; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_33_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_33_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_33_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_33_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_49_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_49_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_49_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_49_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_51_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_51_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_51_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_51_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_53_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_53_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_53_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_53_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_55_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_55_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_55_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_55_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_57_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_57_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_57_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_57_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_59_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_59_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_59_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_59_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_61_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_61_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_61_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_61_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_63_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_63_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_63_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_63_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_65_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_65_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_65_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_65_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_67_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_67_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_67_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_67_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_69_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_69_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_69_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_69_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_71_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_71_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_71_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_71_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_73_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_73_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_73_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_73_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_75_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_75_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_75_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_75_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_77_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_77_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_77_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_77_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_79_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_79_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_79_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_79_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_81_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_81_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_81_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_81_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_83_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_83_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_83_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_83_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_85_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_85_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_85_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_85_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_87_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_87_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_87_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_87_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_89_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_89_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_89_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_89_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_91_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_91_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_91_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_91_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_93_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_93_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_93_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_93_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_95_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_95_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_95_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_95_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_97_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_97_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_97_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_97_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_99_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_99_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_99_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_99_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_101_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_101_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_101_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_101_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_103_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_103_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_103_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_103_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_105_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_105_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_105_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_105_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_107_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_107_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_107_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_107_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_109_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_109_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_109_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_109_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_111_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_111_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_111_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_111_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_113_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_113_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_113_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_113_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_115_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_115_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_115_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_115_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_117_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_117_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_117_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_117_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_119_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_119_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_119_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_119_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_121_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_121_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_121_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_121_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_123_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_123_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_123_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_123_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_125_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_125_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_125_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_125_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_127_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_127_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_127_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_127_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_129_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_129_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_129_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_129_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_131_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_131_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_131_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_131_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_133_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_133_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_133_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_133_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_135_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_135_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_135_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_135_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_137_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_137_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_137_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_137_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_139_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_139_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_139_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_139_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_141_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_141_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_141_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_141_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_143_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_143_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_143_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_143_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_145_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_145_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_145_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_145_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_147_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_147_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_147_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_147_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_149_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_149_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_149_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_149_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_151_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_151_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_151_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_151_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_153_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_153_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_153_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_153_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_155_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_155_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_155_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_155_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_157_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_157_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_157_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_157_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_159_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_159_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_159_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_159_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_161_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_161_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_161_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_161_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_163_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_163_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_163_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_163_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_165_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_165_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_165_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_165_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_167_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_167_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_167_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_167_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_169_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_169_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_169_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_169_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_171_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_171_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_171_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_171_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_173_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_173_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_173_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_173_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_175_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_0_MPORT_175_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_175_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_0_MPORT_175_en; // @[PatternHistoryTable.scala 26:28]
//   reg  pht_0_0_MPORT_17_en_pipe_0;
  reg [5:0] pht_0_0_MPORT_17_addr_pipe_0;
  reg  pht_0_1 [0:63]; // @[PatternHistoryTable.scala 26:28]
//   wire  pht_0_1_MPORT_19_en; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_19_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_19_data; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_35_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_35_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_35_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_35_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_177_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_177_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_177_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_177_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_179_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_179_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_179_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_179_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_181_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_181_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_181_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_181_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_183_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_183_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_183_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_183_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_185_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_185_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_185_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_185_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_187_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_187_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_187_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_187_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_189_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_189_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_189_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_189_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_191_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_191_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_191_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_191_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_193_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_193_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_193_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_193_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_195_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_195_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_195_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_195_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_197_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_197_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_197_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_197_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_199_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_199_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_199_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_199_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_201_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_201_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_201_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_201_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_203_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_203_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_203_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_203_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_205_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_205_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_205_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_205_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_207_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_207_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_207_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_207_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_209_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_209_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_209_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_209_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_211_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_211_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_211_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_211_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_213_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_213_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_213_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_213_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_215_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_215_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_215_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_215_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_217_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_217_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_217_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_217_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_219_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_219_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_219_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_219_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_221_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_221_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_221_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_221_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_223_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_223_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_223_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_223_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_225_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_225_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_225_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_225_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_227_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_227_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_227_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_227_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_229_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_229_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_229_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_229_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_231_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_231_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_231_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_231_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_233_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_233_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_233_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_233_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_235_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_235_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_235_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_235_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_237_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_237_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_237_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_237_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_239_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_239_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_239_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_239_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_241_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_241_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_241_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_241_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_243_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_243_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_243_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_243_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_245_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_245_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_245_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_245_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_247_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_247_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_247_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_247_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_249_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_249_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_249_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_249_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_251_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_251_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_251_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_251_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_253_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_253_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_253_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_253_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_255_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_255_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_255_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_255_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_257_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_257_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_257_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_257_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_259_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_259_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_259_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_259_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_261_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_261_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_261_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_261_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_263_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_263_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_263_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_263_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_265_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_265_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_265_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_265_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_267_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_267_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_267_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_267_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_269_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_269_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_269_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_269_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_271_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_271_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_271_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_271_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_273_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_273_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_273_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_273_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_275_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_275_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_275_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_275_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_277_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_277_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_277_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_277_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_279_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_279_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_279_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_279_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_281_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_281_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_281_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_281_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_283_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_283_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_283_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_283_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_285_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_285_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_285_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_285_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_287_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_287_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_287_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_287_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_289_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_289_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_289_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_289_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_291_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_291_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_291_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_291_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_293_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_293_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_293_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_293_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_295_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_295_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_295_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_295_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_297_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_297_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_297_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_297_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_299_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_299_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_299_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_299_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_301_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_301_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_301_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_301_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_303_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_1_MPORT_303_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_303_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_1_MPORT_303_en; // @[PatternHistoryTable.scala 26:28]
//   reg  pht_0_1_MPORT_19_en_pipe_0;
  reg [5:0] pht_0_1_MPORT_19_addr_pipe_0;
  reg  pht_0_2 [0:63]; // @[PatternHistoryTable.scala 26:28]
//   wire  pht_0_2_MPORT_21_en; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_21_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_21_data; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_37_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_37_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_37_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_37_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_305_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_305_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_305_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_305_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_307_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_307_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_307_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_307_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_309_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_309_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_309_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_309_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_311_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_311_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_311_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_311_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_313_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_313_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_313_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_313_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_315_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_315_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_315_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_315_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_317_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_317_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_317_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_317_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_319_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_319_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_319_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_319_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_321_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_321_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_321_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_321_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_323_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_323_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_323_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_323_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_325_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_325_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_325_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_325_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_327_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_327_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_327_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_327_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_329_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_329_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_329_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_329_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_331_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_331_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_331_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_331_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_333_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_333_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_333_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_333_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_335_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_335_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_335_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_335_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_337_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_337_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_337_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_337_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_339_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_339_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_339_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_339_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_341_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_341_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_341_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_341_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_343_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_343_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_343_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_343_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_345_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_345_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_345_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_345_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_347_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_347_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_347_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_347_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_349_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_349_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_349_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_349_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_351_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_351_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_351_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_351_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_353_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_353_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_353_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_353_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_355_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_355_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_355_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_355_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_357_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_357_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_357_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_357_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_359_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_359_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_359_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_359_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_361_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_361_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_361_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_361_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_363_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_363_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_363_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_363_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_365_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_365_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_365_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_365_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_367_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_367_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_367_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_367_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_369_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_369_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_369_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_369_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_371_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_371_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_371_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_371_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_373_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_373_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_373_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_373_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_375_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_375_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_375_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_375_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_377_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_377_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_377_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_377_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_379_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_379_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_379_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_379_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_381_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_381_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_381_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_381_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_383_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_383_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_383_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_383_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_385_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_385_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_385_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_385_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_387_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_387_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_387_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_387_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_389_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_389_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_389_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_389_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_391_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_391_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_391_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_391_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_393_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_393_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_393_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_393_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_395_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_395_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_395_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_395_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_397_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_397_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_397_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_397_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_399_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_399_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_399_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_399_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_401_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_401_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_401_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_401_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_403_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_403_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_403_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_403_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_405_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_405_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_405_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_405_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_407_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_407_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_407_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_407_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_409_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_409_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_409_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_409_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_411_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_411_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_411_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_411_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_413_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_413_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_413_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_413_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_415_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_415_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_415_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_415_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_417_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_417_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_417_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_417_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_419_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_419_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_419_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_419_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_421_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_421_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_421_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_421_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_423_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_423_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_423_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_423_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_425_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_425_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_425_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_425_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_427_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_427_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_427_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_427_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_429_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_429_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_429_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_429_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_431_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_2_MPORT_431_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_431_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_2_MPORT_431_en; // @[PatternHistoryTable.scala 26:28]
//   reg  pht_0_2_MPORT_21_en_pipe_0;
  reg [5:0] pht_0_2_MPORT_21_addr_pipe_0;
  reg  pht_0_3 [0:63]; // @[PatternHistoryTable.scala 26:28]
//   wire  pht_0_3_MPORT_23_en; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_23_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_23_data; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_39_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_39_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_39_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_39_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_433_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_433_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_433_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_433_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_435_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_435_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_435_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_435_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_437_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_437_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_437_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_437_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_439_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_439_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_439_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_439_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_441_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_441_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_441_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_441_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_443_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_443_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_443_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_443_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_445_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_445_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_445_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_445_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_447_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_447_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_447_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_447_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_449_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_449_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_449_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_449_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_451_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_451_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_451_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_451_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_453_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_453_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_453_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_453_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_455_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_455_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_455_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_455_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_457_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_457_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_457_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_457_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_459_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_459_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_459_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_459_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_461_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_461_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_461_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_461_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_463_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_463_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_463_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_463_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_465_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_465_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_465_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_465_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_467_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_467_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_467_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_467_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_469_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_469_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_469_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_469_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_471_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_471_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_471_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_471_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_473_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_473_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_473_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_473_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_475_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_475_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_475_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_475_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_477_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_477_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_477_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_477_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_479_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_479_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_479_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_479_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_481_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_481_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_481_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_481_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_483_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_483_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_483_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_483_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_485_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_485_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_485_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_485_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_487_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_487_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_487_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_487_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_489_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_489_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_489_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_489_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_491_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_491_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_491_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_491_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_493_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_493_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_493_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_493_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_495_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_495_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_495_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_495_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_497_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_497_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_497_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_497_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_499_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_499_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_499_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_499_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_501_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_501_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_501_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_501_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_503_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_503_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_503_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_503_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_505_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_505_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_505_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_505_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_507_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_507_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_507_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_507_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_509_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_509_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_509_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_509_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_511_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_511_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_511_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_511_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_513_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_513_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_513_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_513_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_515_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_515_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_515_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_515_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_517_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_517_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_517_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_517_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_519_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_519_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_519_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_519_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_521_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_521_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_521_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_521_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_523_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_523_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_523_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_523_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_525_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_525_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_525_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_525_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_527_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_527_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_527_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_527_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_529_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_529_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_529_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_529_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_531_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_531_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_531_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_531_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_533_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_533_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_533_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_533_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_535_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_535_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_535_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_535_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_537_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_537_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_537_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_537_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_539_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_539_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_539_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_539_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_541_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_541_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_541_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_541_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_543_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_543_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_543_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_543_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_545_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_545_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_545_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_545_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_547_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_547_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_547_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_547_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_549_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_549_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_549_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_549_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_551_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_551_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_551_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_551_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_553_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_553_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_553_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_553_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_555_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_555_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_555_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_555_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_557_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_557_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_557_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_557_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_559_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_3_MPORT_559_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_559_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_3_MPORT_559_en; // @[PatternHistoryTable.scala 26:28]
//   reg  pht_0_3_MPORT_23_en_pipe_0;
  reg [5:0] pht_0_3_MPORT_23_addr_pipe_0;
  reg  pht_0_4 [0:63]; // @[PatternHistoryTable.scala 26:28]
//   wire  pht_0_4_MPORT_25_en; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_25_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_25_data; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_41_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_41_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_41_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_41_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_561_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_561_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_561_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_561_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_563_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_563_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_563_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_563_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_565_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_565_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_565_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_565_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_567_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_567_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_567_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_567_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_569_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_569_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_569_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_569_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_571_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_571_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_571_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_571_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_573_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_573_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_573_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_573_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_575_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_575_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_575_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_575_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_577_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_577_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_577_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_577_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_579_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_579_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_579_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_579_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_581_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_581_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_581_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_581_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_583_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_583_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_583_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_583_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_585_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_585_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_585_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_585_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_587_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_587_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_587_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_587_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_589_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_589_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_589_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_589_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_591_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_591_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_591_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_591_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_593_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_593_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_593_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_593_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_595_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_595_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_595_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_595_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_597_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_597_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_597_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_597_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_599_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_599_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_599_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_599_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_601_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_601_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_601_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_601_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_603_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_603_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_603_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_603_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_605_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_605_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_605_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_605_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_607_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_607_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_607_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_607_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_609_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_609_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_609_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_609_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_611_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_611_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_611_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_611_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_613_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_613_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_613_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_613_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_615_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_615_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_615_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_615_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_617_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_617_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_617_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_617_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_619_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_619_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_619_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_619_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_621_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_621_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_621_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_621_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_623_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_623_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_623_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_623_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_625_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_625_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_625_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_625_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_627_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_627_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_627_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_627_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_629_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_629_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_629_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_629_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_631_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_631_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_631_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_631_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_633_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_633_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_633_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_633_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_635_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_635_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_635_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_635_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_637_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_637_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_637_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_637_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_639_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_639_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_639_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_639_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_641_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_641_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_641_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_641_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_643_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_643_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_643_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_643_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_645_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_645_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_645_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_645_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_647_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_647_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_647_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_647_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_649_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_649_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_649_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_649_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_651_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_651_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_651_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_651_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_653_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_653_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_653_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_653_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_655_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_655_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_655_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_655_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_657_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_657_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_657_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_657_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_659_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_659_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_659_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_659_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_661_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_661_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_661_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_661_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_663_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_663_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_663_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_663_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_665_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_665_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_665_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_665_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_667_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_667_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_667_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_667_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_669_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_669_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_669_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_669_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_671_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_671_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_671_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_671_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_673_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_673_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_673_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_673_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_675_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_675_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_675_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_675_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_677_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_677_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_677_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_677_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_679_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_679_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_679_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_679_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_681_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_681_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_681_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_681_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_683_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_683_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_683_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_683_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_685_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_685_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_685_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_685_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_687_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_4_MPORT_687_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_687_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_4_MPORT_687_en; // @[PatternHistoryTable.scala 26:28]
//   reg  pht_0_4_MPORT_25_en_pipe_0;
  reg [5:0] pht_0_4_MPORT_25_addr_pipe_0;
  reg  pht_0_5 [0:63]; // @[PatternHistoryTable.scala 26:28]
//   wire  pht_0_5_MPORT_27_en; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_27_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_27_data; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_43_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_43_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_43_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_43_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_689_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_689_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_689_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_689_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_691_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_691_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_691_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_691_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_693_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_693_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_693_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_693_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_695_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_695_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_695_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_695_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_697_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_697_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_697_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_697_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_699_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_699_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_699_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_699_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_701_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_701_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_701_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_701_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_703_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_703_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_703_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_703_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_705_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_705_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_705_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_705_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_707_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_707_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_707_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_707_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_709_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_709_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_709_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_709_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_711_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_711_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_711_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_711_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_713_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_713_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_713_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_713_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_715_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_715_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_715_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_715_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_717_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_717_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_717_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_717_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_719_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_719_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_719_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_719_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_721_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_721_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_721_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_721_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_723_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_723_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_723_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_723_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_725_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_725_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_725_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_725_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_727_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_727_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_727_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_727_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_729_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_729_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_729_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_729_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_731_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_731_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_731_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_731_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_733_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_733_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_733_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_733_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_735_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_735_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_735_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_735_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_737_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_737_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_737_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_737_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_739_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_739_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_739_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_739_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_741_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_741_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_741_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_741_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_743_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_743_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_743_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_743_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_745_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_745_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_745_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_745_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_747_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_747_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_747_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_747_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_749_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_749_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_749_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_749_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_751_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_751_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_751_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_751_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_753_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_753_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_753_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_753_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_755_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_755_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_755_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_755_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_757_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_757_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_757_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_757_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_759_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_759_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_759_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_759_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_761_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_761_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_761_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_761_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_763_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_763_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_763_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_763_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_765_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_765_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_765_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_765_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_767_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_767_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_767_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_767_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_769_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_769_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_769_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_769_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_771_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_771_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_771_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_771_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_773_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_773_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_773_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_773_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_775_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_775_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_775_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_775_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_777_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_777_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_777_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_777_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_779_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_779_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_779_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_779_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_781_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_781_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_781_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_781_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_783_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_783_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_783_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_783_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_785_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_785_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_785_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_785_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_787_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_787_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_787_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_787_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_789_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_789_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_789_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_789_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_791_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_791_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_791_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_791_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_793_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_793_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_793_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_793_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_795_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_795_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_795_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_795_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_797_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_797_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_797_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_797_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_799_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_799_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_799_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_799_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_801_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_801_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_801_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_801_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_803_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_803_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_803_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_803_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_805_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_805_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_805_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_805_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_807_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_807_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_807_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_807_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_809_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_809_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_809_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_809_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_811_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_811_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_811_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_811_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_813_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_813_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_813_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_813_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_815_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_5_MPORT_815_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_815_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_5_MPORT_815_en; // @[PatternHistoryTable.scala 26:28]
//   reg  pht_0_5_MPORT_27_en_pipe_0;
  reg [5:0] pht_0_5_MPORT_27_addr_pipe_0;
  reg  pht_0_6 [0:63]; // @[PatternHistoryTable.scala 26:28]
//   wire  pht_0_6_MPORT_29_en; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_29_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_29_data; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_45_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_45_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_45_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_45_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_817_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_817_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_817_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_817_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_819_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_819_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_819_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_819_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_821_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_821_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_821_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_821_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_823_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_823_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_823_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_823_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_825_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_825_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_825_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_825_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_827_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_827_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_827_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_827_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_829_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_829_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_829_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_829_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_831_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_831_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_831_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_831_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_833_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_833_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_833_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_833_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_835_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_835_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_835_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_835_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_837_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_837_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_837_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_837_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_839_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_839_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_839_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_839_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_841_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_841_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_841_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_841_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_843_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_843_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_843_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_843_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_845_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_845_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_845_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_845_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_847_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_847_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_847_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_847_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_849_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_849_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_849_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_849_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_851_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_851_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_851_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_851_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_853_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_853_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_853_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_853_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_855_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_855_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_855_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_855_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_857_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_857_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_857_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_857_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_859_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_859_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_859_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_859_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_861_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_861_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_861_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_861_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_863_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_863_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_863_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_863_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_865_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_865_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_865_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_865_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_867_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_867_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_867_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_867_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_869_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_869_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_869_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_869_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_871_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_871_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_871_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_871_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_873_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_873_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_873_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_873_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_875_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_875_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_875_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_875_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_877_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_877_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_877_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_877_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_879_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_879_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_879_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_879_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_881_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_881_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_881_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_881_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_883_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_883_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_883_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_883_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_885_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_885_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_885_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_885_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_887_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_887_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_887_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_887_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_889_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_889_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_889_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_889_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_891_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_891_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_891_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_891_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_893_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_893_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_893_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_893_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_895_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_895_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_895_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_895_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_897_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_897_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_897_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_897_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_899_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_899_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_899_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_899_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_901_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_901_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_901_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_901_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_903_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_903_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_903_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_903_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_905_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_905_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_905_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_905_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_907_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_907_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_907_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_907_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_909_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_909_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_909_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_909_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_911_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_911_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_911_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_911_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_913_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_913_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_913_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_913_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_915_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_915_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_915_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_915_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_917_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_917_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_917_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_917_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_919_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_919_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_919_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_919_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_921_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_921_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_921_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_921_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_923_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_923_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_923_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_923_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_925_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_925_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_925_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_925_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_927_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_927_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_927_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_927_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_929_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_929_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_929_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_929_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_931_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_931_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_931_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_931_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_933_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_933_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_933_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_933_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_935_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_935_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_935_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_935_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_937_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_937_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_937_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_937_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_939_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_939_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_939_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_939_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_941_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_941_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_941_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_941_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_943_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_6_MPORT_943_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_943_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_6_MPORT_943_en; // @[PatternHistoryTable.scala 26:28]
//   reg  pht_0_6_MPORT_29_en_pipe_0;
  reg [5:0] pht_0_6_MPORT_29_addr_pipe_0;
  reg  pht_0_7 [0:63]; // @[PatternHistoryTable.scala 26:28]
//   wire  pht_0_7_MPORT_31_en; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_31_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_31_data; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_47_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_47_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_47_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_47_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_945_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_945_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_945_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_945_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_947_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_947_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_947_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_947_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_949_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_949_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_949_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_949_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_951_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_951_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_951_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_951_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_953_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_953_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_953_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_953_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_955_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_955_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_955_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_955_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_957_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_957_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_957_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_957_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_959_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_959_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_959_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_959_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_961_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_961_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_961_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_961_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_963_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_963_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_963_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_963_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_965_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_965_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_965_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_965_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_967_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_967_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_967_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_967_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_969_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_969_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_969_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_969_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_971_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_971_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_971_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_971_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_973_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_973_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_973_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_973_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_975_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_975_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_975_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_975_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_977_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_977_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_977_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_977_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_979_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_979_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_979_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_979_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_981_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_981_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_981_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_981_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_983_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_983_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_983_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_983_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_985_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_985_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_985_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_985_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_987_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_987_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_987_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_987_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_989_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_989_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_989_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_989_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_991_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_991_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_991_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_991_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_993_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_993_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_993_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_993_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_995_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_995_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_995_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_995_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_997_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_997_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_997_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_997_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_999_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_999_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_999_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_999_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1001_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1001_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1001_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1001_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1003_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1003_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1003_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1003_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1005_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1005_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1005_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1005_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1007_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1007_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1007_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1007_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1009_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1009_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1009_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1009_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1011_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1011_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1011_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1011_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1013_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1013_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1013_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1013_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1015_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1015_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1015_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1015_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1017_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1017_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1017_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1017_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1019_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1019_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1019_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1019_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1021_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1021_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1021_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1021_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1023_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1023_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1023_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1023_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1025_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1025_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1025_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1025_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1027_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1027_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1027_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1027_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1029_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1029_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1029_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1029_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1031_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1031_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1031_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1031_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1033_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1033_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1033_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1033_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1035_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1035_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1035_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1035_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1037_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1037_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1037_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1037_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1039_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1039_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1039_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1039_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1041_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1041_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1041_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1041_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1043_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1043_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1043_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1043_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1045_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1045_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1045_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1045_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1047_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1047_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1047_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1047_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1049_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1049_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1049_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1049_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1051_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1051_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1051_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1051_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1053_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1053_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1053_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1053_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1055_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1055_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1055_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1055_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1057_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1057_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1057_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1057_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1059_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1059_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1059_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1059_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1061_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1061_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1061_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1061_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1063_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1063_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1063_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1063_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1065_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1065_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1065_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1065_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1067_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1067_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1067_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1067_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1069_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1069_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1069_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1069_en; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1071_data; // @[PatternHistoryTable.scala 26:28]
  wire [5:0] pht_0_7_MPORT_1071_addr; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1071_mask; // @[PatternHistoryTable.scala 26:28]
  wire  pht_0_7_MPORT_1071_en; // @[PatternHistoryTable.scala 26:28]
//   reg  pht_0_7_MPORT_31_en_pipe_0;
  reg [5:0] pht_0_7_MPORT_31_addr_pipe_0;
  reg [2:0] REG; // @[PatternHistoryTable.scala 42:20]
  wire  _GEN_11 = REG == 3'h0 & pht_1_0_MPORT_data; // @[PatternHistoryTable.scala 40:19 42:44 43:23]
  reg [2:0] REG_1; // @[PatternHistoryTable.scala 42:20]
  wire  _GEN_12 = REG_1 == 3'h1 ? pht_1_1_MPORT_1_data : _GEN_11; // @[PatternHistoryTable.scala 42:44 43:23]
  reg [2:0] REG_2; // @[PatternHistoryTable.scala 42:20]
  wire  _GEN_13 = REG_2 == 3'h2 ? pht_1_2_MPORT_2_data : _GEN_12; // @[PatternHistoryTable.scala 42:44 43:23]
  reg [2:0] REG_3; // @[PatternHistoryTable.scala 42:20]
  wire  _GEN_14 = REG_3 == 3'h3 ? pht_1_3_MPORT_3_data : _GEN_13; // @[PatternHistoryTable.scala 42:44 43:23]
  reg [2:0] REG_4; // @[PatternHistoryTable.scala 42:20]
  wire  _GEN_15 = REG_4 == 3'h4 ? pht_1_4_MPORT_4_data : _GEN_14; // @[PatternHistoryTable.scala 42:44 43:23]
  reg [2:0] REG_5; // @[PatternHistoryTable.scala 42:20]
  wire  _GEN_16 = REG_5 == 3'h5 ? pht_1_5_MPORT_5_data : _GEN_15; // @[PatternHistoryTable.scala 42:44 43:23]
  reg [2:0] REG_6; // @[PatternHistoryTable.scala 42:20]
  wire  _GEN_17 = REG_6 == 3'h6 ? pht_1_6_MPORT_6_data : _GEN_16; // @[PatternHistoryTable.scala 42:44 43:23]
  reg [2:0] REG_7; // @[PatternHistoryTable.scala 42:20]
  reg [2:0] REG_8; // @[PatternHistoryTable.scala 42:20]
  wire  _GEN_28 = REG_8 == 3'h0 & pht_1_0_MPORT_8_data; // @[PatternHistoryTable.scala 40:19 42:44 43:23]
  reg [2:0] REG_9; // @[PatternHistoryTable.scala 42:20]
  wire  _GEN_29 = REG_9 == 3'h1 ? pht_1_1_MPORT_9_data : _GEN_28; // @[PatternHistoryTable.scala 42:44 43:23]
  reg [2:0] REG_10; // @[PatternHistoryTable.scala 42:20]
  wire  _GEN_30 = REG_10 == 3'h2 ? pht_1_2_MPORT_10_data : _GEN_29; // @[PatternHistoryTable.scala 42:44 43:23]
  reg [2:0] REG_11; // @[PatternHistoryTable.scala 42:20]
  wire  _GEN_31 = REG_11 == 3'h3 ? pht_1_3_MPORT_11_data : _GEN_30; // @[PatternHistoryTable.scala 42:44 43:23]
  reg [2:0] REG_12; // @[PatternHistoryTable.scala 42:20]
  wire  _GEN_32 = REG_12 == 3'h4 ? pht_1_4_MPORT_12_data : _GEN_31; // @[PatternHistoryTable.scala 42:44 43:23]
  reg [2:0] REG_13; // @[PatternHistoryTable.scala 42:20]
  wire  _GEN_33 = REG_13 == 3'h5 ? pht_1_5_MPORT_13_data : _GEN_32; // @[PatternHistoryTable.scala 42:44 43:23]
  reg [2:0] REG_14; // @[PatternHistoryTable.scala 42:20]
  wire  _GEN_34 = REG_14 == 3'h6 ? pht_1_6_MPORT_14_data : _GEN_33; // @[PatternHistoryTable.scala 42:44 43:23]
  reg [2:0] REG_15; // @[PatternHistoryTable.scala 42:20]
  wire [1:0] pht_wdata_0 = {pht_1_0_MPORT_16_data,pht_0_0_MPORT_17_data}; // @[Cat.scala 30:58]
  wire [1:0] pht_wdata_1 = {pht_1_1_MPORT_18_data,pht_0_1_MPORT_19_data}; // @[Cat.scala 30:58]
  wire [1:0] pht_wdata_2 = {pht_1_2_MPORT_20_data,pht_0_2_MPORT_21_data}; // @[Cat.scala 30:58]
  wire [1:0] pht_wdata_3 = {pht_1_3_MPORT_22_data,pht_0_3_MPORT_23_data}; // @[Cat.scala 30:58]
  wire [1:0] pht_wdata_4 = {pht_1_4_MPORT_24_data,pht_0_4_MPORT_25_data}; // @[Cat.scala 30:58]
  wire [1:0] pht_wdata_5 = {pht_1_5_MPORT_26_data,pht_0_5_MPORT_27_data}; // @[Cat.scala 30:58]
  wire [1:0] pht_wdata_6 = {pht_1_6_MPORT_28_data,pht_0_6_MPORT_29_data}; // @[Cat.scala 30:58]
  wire [1:0] pht_wdata_7 = {pht_1_7_MPORT_30_data,pht_0_7_MPORT_31_data}; // @[Cat.scala 30:58]
  reg  REG_16; // @[PatternHistoryTable.scala 59:16]
  reg [2:0] REG_17; // @[PatternHistoryTable.scala 61:20]
  wire [1:0] _GEN_53 = REG_17 == 3'h0 ? pht_wdata_0 : 2'h0; // @[PatternHistoryTable.scala 61:41 62:21]
  reg [2:0] REG_18; // @[PatternHistoryTable.scala 61:20]
  wire [1:0] _GEN_54 = REG_18 == 3'h1 ? pht_wdata_1 : _GEN_53; // @[PatternHistoryTable.scala 61:41 62:21]
  reg [2:0] REG_19; // @[PatternHistoryTable.scala 61:20]
  wire [1:0] _GEN_55 = REG_19 == 3'h2 ? pht_wdata_2 : _GEN_54; // @[PatternHistoryTable.scala 61:41 62:21]
  reg [2:0] REG_20; // @[PatternHistoryTable.scala 61:20]
  wire [1:0] _GEN_56 = REG_20 == 3'h3 ? pht_wdata_3 : _GEN_55; // @[PatternHistoryTable.scala 61:41 62:21]
  reg [2:0] REG_21; // @[PatternHistoryTable.scala 61:20]
  wire [1:0] _GEN_57 = REG_21 == 3'h4 ? pht_wdata_4 : _GEN_56; // @[PatternHistoryTable.scala 61:41 62:21]
  reg [2:0] REG_22; // @[PatternHistoryTable.scala 61:20]
  wire [1:0] _GEN_58 = REG_22 == 3'h5 ? pht_wdata_5 : _GEN_57; // @[PatternHistoryTable.scala 61:41 62:21]
  reg [2:0] REG_23; // @[PatternHistoryTable.scala 61:20]
  wire [1:0] _GEN_59 = REG_23 == 3'h6 ? pht_wdata_6 : _GEN_58; // @[PatternHistoryTable.scala 61:41 62:21]
  reg [2:0] REG_24; // @[PatternHistoryTable.scala 61:20]
  wire [1:0] _GEN_60 = REG_24 == 3'h7 ? pht_wdata_7 : _GEN_59; // @[PatternHistoryTable.scala 61:41 62:21]
  wire [1:0] pht_wdata_r = REG_16 ? _GEN_60 : 2'h0; // @[PatternHistoryTable.scala 59:26]
  reg  REG_25; // @[PatternHistoryTable.scala 67:23]
  reg  REG_26; // @[PatternHistoryTable.scala 68:23]
  wire [1:0] _T_113 = REG_26 ? 2'h2 : 2'h0; // @[PatternHistoryTable.scala 68:15]
  reg  REG_27; // @[PatternHistoryTable.scala 69:23]
  wire [1:0] _T_114 = REG_27 ? 2'h3 : 2'h1; // @[PatternHistoryTable.scala 69:15]
  reg  REG_28; // @[PatternHistoryTable.scala 70:23]
  wire [1:0] _T_115 = REG_28 ? 2'h3 : 2'h2; // @[PatternHistoryTable.scala 70:15]
  wire [1:0] _T_117 = 2'h1 == pht_wdata_r ? _T_113 : {{1'd0}, REG_25}; // @[Mux.scala 80:57]
  wire [1:0] _T_119 = 2'h2 == pht_wdata_r ? _T_114 : _T_117; // @[Mux.scala 80:57]
  wire [1:0] pht_wdata_w = 2'h3 == pht_wdata_r ? _T_115 : _T_119; // @[Mux.scala 80:57]
  reg  REG_29; // @[PatternHistoryTable.scala 72:16]
  reg  REG_30; // @[PatternHistoryTable.scala 74:20]
  reg [5:0] REG_31; // @[PatternHistoryTable.scala 75:31]
  reg [5:0] REG_32; // @[PatternHistoryTable.scala 76:31]
  reg  REG_33; // @[PatternHistoryTable.scala 74:20]
  reg [5:0] REG_34; // @[PatternHistoryTable.scala 75:31]
  reg [5:0] REG_35; // @[PatternHistoryTable.scala 76:31]
  reg  REG_36; // @[PatternHistoryTable.scala 74:20]
  reg [5:0] REG_37; // @[PatternHistoryTable.scala 75:31]
  reg [5:0] REG_38; // @[PatternHistoryTable.scala 76:31]
  reg  REG_39; // @[PatternHistoryTable.scala 74:20]
  reg [5:0] REG_40; // @[PatternHistoryTable.scala 75:31]
  reg [5:0] REG_41; // @[PatternHistoryTable.scala 76:31]
  reg  REG_42; // @[PatternHistoryTable.scala 74:20]
  reg [5:0] REG_43; // @[PatternHistoryTable.scala 75:31]
  reg [5:0] REG_44; // @[PatternHistoryTable.scala 76:31]
  reg  REG_45; // @[PatternHistoryTable.scala 74:20]
  reg [5:0] REG_46; // @[PatternHistoryTable.scala 75:31]
  reg [5:0] REG_47; // @[PatternHistoryTable.scala 76:31]
  reg  REG_48; // @[PatternHistoryTable.scala 74:20]
  reg [5:0] REG_49; // @[PatternHistoryTable.scala 75:31]
  reg [5:0] REG_50; // @[PatternHistoryTable.scala 76:31]
  reg  REG_51; // @[PatternHistoryTable.scala 74:20]
  reg [5:0] REG_52; // @[PatternHistoryTable.scala 75:31]
  reg [5:0] REG_53; // @[PatternHistoryTable.scala 76:31]
//   assign pht_1_0_MPORT_en = pht_1_0_MPORT_en_pipe_0;
  assign pht_1_0_MPORT_addr = pht_1_0_MPORT_addr_pipe_0;
  assign pht_1_0_MPORT_data = pht_1_0[pht_1_0_MPORT_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_0_MPORT_8_en = pht_1_0_MPORT_8_en_pipe_0;
  assign pht_1_0_MPORT_8_addr = pht_1_0_MPORT_8_addr_pipe_0;
  assign pht_1_0_MPORT_8_data = pht_1_0[pht_1_0_MPORT_8_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_0_MPORT_16_en = pht_1_0_MPORT_16_en_pipe_0;
  assign pht_1_0_MPORT_16_addr = pht_1_0_MPORT_16_addr_pipe_0;
  assign pht_1_0_MPORT_16_data = pht_1_0[pht_1_0_MPORT_16_addr]; // @[PatternHistoryTable.scala 21:28]
  assign pht_1_0_MPORT_32_data = pht_wdata_w[1];
  assign pht_1_0_MPORT_32_addr = REG_31;
  assign pht_1_0_MPORT_32_mask = 1'h1;
  assign pht_1_0_MPORT_32_en = REG_29 & REG_30;
  assign pht_1_0_MPORT_48_data = 1'h0;
  assign pht_1_0_MPORT_48_addr = 6'h0;
  assign pht_1_0_MPORT_48_mask = 1'h1;
  assign pht_1_0_MPORT_48_en = reset;
  assign pht_1_0_MPORT_50_data = 1'h0;
  assign pht_1_0_MPORT_50_addr = 6'h1;
  assign pht_1_0_MPORT_50_mask = 1'h1;
  assign pht_1_0_MPORT_50_en = reset;
  assign pht_1_0_MPORT_52_data = 1'h0;
  assign pht_1_0_MPORT_52_addr = 6'h2;
  assign pht_1_0_MPORT_52_mask = 1'h1;
  assign pht_1_0_MPORT_52_en = reset;
  assign pht_1_0_MPORT_54_data = 1'h0;
  assign pht_1_0_MPORT_54_addr = 6'h3;
  assign pht_1_0_MPORT_54_mask = 1'h1;
  assign pht_1_0_MPORT_54_en = reset;
  assign pht_1_0_MPORT_56_data = 1'h0;
  assign pht_1_0_MPORT_56_addr = 6'h4;
  assign pht_1_0_MPORT_56_mask = 1'h1;
  assign pht_1_0_MPORT_56_en = reset;
  assign pht_1_0_MPORT_58_data = 1'h0;
  assign pht_1_0_MPORT_58_addr = 6'h5;
  assign pht_1_0_MPORT_58_mask = 1'h1;
  assign pht_1_0_MPORT_58_en = reset;
  assign pht_1_0_MPORT_60_data = 1'h0;
  assign pht_1_0_MPORT_60_addr = 6'h6;
  assign pht_1_0_MPORT_60_mask = 1'h1;
  assign pht_1_0_MPORT_60_en = reset;
  assign pht_1_0_MPORT_62_data = 1'h0;
  assign pht_1_0_MPORT_62_addr = 6'h7;
  assign pht_1_0_MPORT_62_mask = 1'h1;
  assign pht_1_0_MPORT_62_en = reset;
  assign pht_1_0_MPORT_64_data = 1'h0;
  assign pht_1_0_MPORT_64_addr = 6'h8;
  assign pht_1_0_MPORT_64_mask = 1'h1;
  assign pht_1_0_MPORT_64_en = reset;
  assign pht_1_0_MPORT_66_data = 1'h0;
  assign pht_1_0_MPORT_66_addr = 6'h9;
  assign pht_1_0_MPORT_66_mask = 1'h1;
  assign pht_1_0_MPORT_66_en = reset;
  assign pht_1_0_MPORT_68_data = 1'h0;
  assign pht_1_0_MPORT_68_addr = 6'ha;
  assign pht_1_0_MPORT_68_mask = 1'h1;
  assign pht_1_0_MPORT_68_en = reset;
  assign pht_1_0_MPORT_70_data = 1'h0;
  assign pht_1_0_MPORT_70_addr = 6'hb;
  assign pht_1_0_MPORT_70_mask = 1'h1;
  assign pht_1_0_MPORT_70_en = reset;
  assign pht_1_0_MPORT_72_data = 1'h0;
  assign pht_1_0_MPORT_72_addr = 6'hc;
  assign pht_1_0_MPORT_72_mask = 1'h1;
  assign pht_1_0_MPORT_72_en = reset;
  assign pht_1_0_MPORT_74_data = 1'h0;
  assign pht_1_0_MPORT_74_addr = 6'hd;
  assign pht_1_0_MPORT_74_mask = 1'h1;
  assign pht_1_0_MPORT_74_en = reset;
  assign pht_1_0_MPORT_76_data = 1'h0;
  assign pht_1_0_MPORT_76_addr = 6'he;
  assign pht_1_0_MPORT_76_mask = 1'h1;
  assign pht_1_0_MPORT_76_en = reset;
  assign pht_1_0_MPORT_78_data = 1'h0;
  assign pht_1_0_MPORT_78_addr = 6'hf;
  assign pht_1_0_MPORT_78_mask = 1'h1;
  assign pht_1_0_MPORT_78_en = reset;
  assign pht_1_0_MPORT_80_data = 1'h0;
  assign pht_1_0_MPORT_80_addr = 6'h10;
  assign pht_1_0_MPORT_80_mask = 1'h1;
  assign pht_1_0_MPORT_80_en = reset;
  assign pht_1_0_MPORT_82_data = 1'h0;
  assign pht_1_0_MPORT_82_addr = 6'h11;
  assign pht_1_0_MPORT_82_mask = 1'h1;
  assign pht_1_0_MPORT_82_en = reset;
  assign pht_1_0_MPORT_84_data = 1'h0;
  assign pht_1_0_MPORT_84_addr = 6'h12;
  assign pht_1_0_MPORT_84_mask = 1'h1;
  assign pht_1_0_MPORT_84_en = reset;
  assign pht_1_0_MPORT_86_data = 1'h0;
  assign pht_1_0_MPORT_86_addr = 6'h13;
  assign pht_1_0_MPORT_86_mask = 1'h1;
  assign pht_1_0_MPORT_86_en = reset;
  assign pht_1_0_MPORT_88_data = 1'h0;
  assign pht_1_0_MPORT_88_addr = 6'h14;
  assign pht_1_0_MPORT_88_mask = 1'h1;
  assign pht_1_0_MPORT_88_en = reset;
  assign pht_1_0_MPORT_90_data = 1'h0;
  assign pht_1_0_MPORT_90_addr = 6'h15;
  assign pht_1_0_MPORT_90_mask = 1'h1;
  assign pht_1_0_MPORT_90_en = reset;
  assign pht_1_0_MPORT_92_data = 1'h0;
  assign pht_1_0_MPORT_92_addr = 6'h16;
  assign pht_1_0_MPORT_92_mask = 1'h1;
  assign pht_1_0_MPORT_92_en = reset;
  assign pht_1_0_MPORT_94_data = 1'h0;
  assign pht_1_0_MPORT_94_addr = 6'h17;
  assign pht_1_0_MPORT_94_mask = 1'h1;
  assign pht_1_0_MPORT_94_en = reset;
  assign pht_1_0_MPORT_96_data = 1'h0;
  assign pht_1_0_MPORT_96_addr = 6'h18;
  assign pht_1_0_MPORT_96_mask = 1'h1;
  assign pht_1_0_MPORT_96_en = reset;
  assign pht_1_0_MPORT_98_data = 1'h0;
  assign pht_1_0_MPORT_98_addr = 6'h19;
  assign pht_1_0_MPORT_98_mask = 1'h1;
  assign pht_1_0_MPORT_98_en = reset;
  assign pht_1_0_MPORT_100_data = 1'h0;
  assign pht_1_0_MPORT_100_addr = 6'h1a;
  assign pht_1_0_MPORT_100_mask = 1'h1;
  assign pht_1_0_MPORT_100_en = reset;
  assign pht_1_0_MPORT_102_data = 1'h0;
  assign pht_1_0_MPORT_102_addr = 6'h1b;
  assign pht_1_0_MPORT_102_mask = 1'h1;
  assign pht_1_0_MPORT_102_en = reset;
  assign pht_1_0_MPORT_104_data = 1'h0;
  assign pht_1_0_MPORT_104_addr = 6'h1c;
  assign pht_1_0_MPORT_104_mask = 1'h1;
  assign pht_1_0_MPORT_104_en = reset;
  assign pht_1_0_MPORT_106_data = 1'h0;
  assign pht_1_0_MPORT_106_addr = 6'h1d;
  assign pht_1_0_MPORT_106_mask = 1'h1;
  assign pht_1_0_MPORT_106_en = reset;
  assign pht_1_0_MPORT_108_data = 1'h0;
  assign pht_1_0_MPORT_108_addr = 6'h1e;
  assign pht_1_0_MPORT_108_mask = 1'h1;
  assign pht_1_0_MPORT_108_en = reset;
  assign pht_1_0_MPORT_110_data = 1'h0;
  assign pht_1_0_MPORT_110_addr = 6'h1f;
  assign pht_1_0_MPORT_110_mask = 1'h1;
  assign pht_1_0_MPORT_110_en = reset;
  assign pht_1_0_MPORT_112_data = 1'h0;
  assign pht_1_0_MPORT_112_addr = 6'h20;
  assign pht_1_0_MPORT_112_mask = 1'h1;
  assign pht_1_0_MPORT_112_en = reset;
  assign pht_1_0_MPORT_114_data = 1'h0;
  assign pht_1_0_MPORT_114_addr = 6'h21;
  assign pht_1_0_MPORT_114_mask = 1'h1;
  assign pht_1_0_MPORT_114_en = reset;
  assign pht_1_0_MPORT_116_data = 1'h0;
  assign pht_1_0_MPORT_116_addr = 6'h22;
  assign pht_1_0_MPORT_116_mask = 1'h1;
  assign pht_1_0_MPORT_116_en = reset;
  assign pht_1_0_MPORT_118_data = 1'h0;
  assign pht_1_0_MPORT_118_addr = 6'h23;
  assign pht_1_0_MPORT_118_mask = 1'h1;
  assign pht_1_0_MPORT_118_en = reset;
  assign pht_1_0_MPORT_120_data = 1'h0;
  assign pht_1_0_MPORT_120_addr = 6'h24;
  assign pht_1_0_MPORT_120_mask = 1'h1;
  assign pht_1_0_MPORT_120_en = reset;
  assign pht_1_0_MPORT_122_data = 1'h0;
  assign pht_1_0_MPORT_122_addr = 6'h25;
  assign pht_1_0_MPORT_122_mask = 1'h1;
  assign pht_1_0_MPORT_122_en = reset;
  assign pht_1_0_MPORT_124_data = 1'h0;
  assign pht_1_0_MPORT_124_addr = 6'h26;
  assign pht_1_0_MPORT_124_mask = 1'h1;
  assign pht_1_0_MPORT_124_en = reset;
  assign pht_1_0_MPORT_126_data = 1'h0;
  assign pht_1_0_MPORT_126_addr = 6'h27;
  assign pht_1_0_MPORT_126_mask = 1'h1;
  assign pht_1_0_MPORT_126_en = reset;
  assign pht_1_0_MPORT_128_data = 1'h0;
  assign pht_1_0_MPORT_128_addr = 6'h28;
  assign pht_1_0_MPORT_128_mask = 1'h1;
  assign pht_1_0_MPORT_128_en = reset;
  assign pht_1_0_MPORT_130_data = 1'h0;
  assign pht_1_0_MPORT_130_addr = 6'h29;
  assign pht_1_0_MPORT_130_mask = 1'h1;
  assign pht_1_0_MPORT_130_en = reset;
  assign pht_1_0_MPORT_132_data = 1'h0;
  assign pht_1_0_MPORT_132_addr = 6'h2a;
  assign pht_1_0_MPORT_132_mask = 1'h1;
  assign pht_1_0_MPORT_132_en = reset;
  assign pht_1_0_MPORT_134_data = 1'h0;
  assign pht_1_0_MPORT_134_addr = 6'h2b;
  assign pht_1_0_MPORT_134_mask = 1'h1;
  assign pht_1_0_MPORT_134_en = reset;
  assign pht_1_0_MPORT_136_data = 1'h0;
  assign pht_1_0_MPORT_136_addr = 6'h2c;
  assign pht_1_0_MPORT_136_mask = 1'h1;
  assign pht_1_0_MPORT_136_en = reset;
  assign pht_1_0_MPORT_138_data = 1'h0;
  assign pht_1_0_MPORT_138_addr = 6'h2d;
  assign pht_1_0_MPORT_138_mask = 1'h1;
  assign pht_1_0_MPORT_138_en = reset;
  assign pht_1_0_MPORT_140_data = 1'h0;
  assign pht_1_0_MPORT_140_addr = 6'h2e;
  assign pht_1_0_MPORT_140_mask = 1'h1;
  assign pht_1_0_MPORT_140_en = reset;
  assign pht_1_0_MPORT_142_data = 1'h0;
  assign pht_1_0_MPORT_142_addr = 6'h2f;
  assign pht_1_0_MPORT_142_mask = 1'h1;
  assign pht_1_0_MPORT_142_en = reset;
  assign pht_1_0_MPORT_144_data = 1'h0;
  assign pht_1_0_MPORT_144_addr = 6'h30;
  assign pht_1_0_MPORT_144_mask = 1'h1;
  assign pht_1_0_MPORT_144_en = reset;
  assign pht_1_0_MPORT_146_data = 1'h0;
  assign pht_1_0_MPORT_146_addr = 6'h31;
  assign pht_1_0_MPORT_146_mask = 1'h1;
  assign pht_1_0_MPORT_146_en = reset;
  assign pht_1_0_MPORT_148_data = 1'h0;
  assign pht_1_0_MPORT_148_addr = 6'h32;
  assign pht_1_0_MPORT_148_mask = 1'h1;
  assign pht_1_0_MPORT_148_en = reset;
  assign pht_1_0_MPORT_150_data = 1'h0;
  assign pht_1_0_MPORT_150_addr = 6'h33;
  assign pht_1_0_MPORT_150_mask = 1'h1;
  assign pht_1_0_MPORT_150_en = reset;
  assign pht_1_0_MPORT_152_data = 1'h0;
  assign pht_1_0_MPORT_152_addr = 6'h34;
  assign pht_1_0_MPORT_152_mask = 1'h1;
  assign pht_1_0_MPORT_152_en = reset;
  assign pht_1_0_MPORT_154_data = 1'h0;
  assign pht_1_0_MPORT_154_addr = 6'h35;
  assign pht_1_0_MPORT_154_mask = 1'h1;
  assign pht_1_0_MPORT_154_en = reset;
  assign pht_1_0_MPORT_156_data = 1'h0;
  assign pht_1_0_MPORT_156_addr = 6'h36;
  assign pht_1_0_MPORT_156_mask = 1'h1;
  assign pht_1_0_MPORT_156_en = reset;
  assign pht_1_0_MPORT_158_data = 1'h0;
  assign pht_1_0_MPORT_158_addr = 6'h37;
  assign pht_1_0_MPORT_158_mask = 1'h1;
  assign pht_1_0_MPORT_158_en = reset;
  assign pht_1_0_MPORT_160_data = 1'h0;
  assign pht_1_0_MPORT_160_addr = 6'h38;
  assign pht_1_0_MPORT_160_mask = 1'h1;
  assign pht_1_0_MPORT_160_en = reset;
  assign pht_1_0_MPORT_162_data = 1'h0;
  assign pht_1_0_MPORT_162_addr = 6'h39;
  assign pht_1_0_MPORT_162_mask = 1'h1;
  assign pht_1_0_MPORT_162_en = reset;
  assign pht_1_0_MPORT_164_data = 1'h0;
  assign pht_1_0_MPORT_164_addr = 6'h3a;
  assign pht_1_0_MPORT_164_mask = 1'h1;
  assign pht_1_0_MPORT_164_en = reset;
  assign pht_1_0_MPORT_166_data = 1'h0;
  assign pht_1_0_MPORT_166_addr = 6'h3b;
  assign pht_1_0_MPORT_166_mask = 1'h1;
  assign pht_1_0_MPORT_166_en = reset;
  assign pht_1_0_MPORT_168_data = 1'h0;
  assign pht_1_0_MPORT_168_addr = 6'h3c;
  assign pht_1_0_MPORT_168_mask = 1'h1;
  assign pht_1_0_MPORT_168_en = reset;
  assign pht_1_0_MPORT_170_data = 1'h0;
  assign pht_1_0_MPORT_170_addr = 6'h3d;
  assign pht_1_0_MPORT_170_mask = 1'h1;
  assign pht_1_0_MPORT_170_en = reset;
  assign pht_1_0_MPORT_172_data = 1'h0;
  assign pht_1_0_MPORT_172_addr = 6'h3e;
  assign pht_1_0_MPORT_172_mask = 1'h1;
  assign pht_1_0_MPORT_172_en = reset;
  assign pht_1_0_MPORT_174_data = 1'h0;
  assign pht_1_0_MPORT_174_addr = 6'h3f;
  assign pht_1_0_MPORT_174_mask = 1'h1;
  assign pht_1_0_MPORT_174_en = reset;
//   assign pht_1_1_MPORT_1_en = pht_1_1_MPORT_1_en_pipe_0;
  assign pht_1_1_MPORT_1_addr = pht_1_1_MPORT_1_addr_pipe_0;
  assign pht_1_1_MPORT_1_data = pht_1_1[pht_1_1_MPORT_1_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_1_MPORT_9_en = pht_1_1_MPORT_9_en_pipe_0;
  assign pht_1_1_MPORT_9_addr = pht_1_1_MPORT_9_addr_pipe_0;
  assign pht_1_1_MPORT_9_data = pht_1_1[pht_1_1_MPORT_9_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_1_MPORT_18_en = pht_1_1_MPORT_18_en_pipe_0;
  assign pht_1_1_MPORT_18_addr = pht_1_1_MPORT_18_addr_pipe_0;
  assign pht_1_1_MPORT_18_data = pht_1_1[pht_1_1_MPORT_18_addr]; // @[PatternHistoryTable.scala 21:28]
  assign pht_1_1_MPORT_34_data = pht_wdata_w[1];
  assign pht_1_1_MPORT_34_addr = REG_34;
  assign pht_1_1_MPORT_34_mask = 1'h1;
  assign pht_1_1_MPORT_34_en = REG_29 & REG_33;
  assign pht_1_1_MPORT_176_data = 1'h0;
  assign pht_1_1_MPORT_176_addr = 6'h0;
  assign pht_1_1_MPORT_176_mask = 1'h1;
  assign pht_1_1_MPORT_176_en = reset;
  assign pht_1_1_MPORT_178_data = 1'h0;
  assign pht_1_1_MPORT_178_addr = 6'h1;
  assign pht_1_1_MPORT_178_mask = 1'h1;
  assign pht_1_1_MPORT_178_en = reset;
  assign pht_1_1_MPORT_180_data = 1'h0;
  assign pht_1_1_MPORT_180_addr = 6'h2;
  assign pht_1_1_MPORT_180_mask = 1'h1;
  assign pht_1_1_MPORT_180_en = reset;
  assign pht_1_1_MPORT_182_data = 1'h0;
  assign pht_1_1_MPORT_182_addr = 6'h3;
  assign pht_1_1_MPORT_182_mask = 1'h1;
  assign pht_1_1_MPORT_182_en = reset;
  assign pht_1_1_MPORT_184_data = 1'h0;
  assign pht_1_1_MPORT_184_addr = 6'h4;
  assign pht_1_1_MPORT_184_mask = 1'h1;
  assign pht_1_1_MPORT_184_en = reset;
  assign pht_1_1_MPORT_186_data = 1'h0;
  assign pht_1_1_MPORT_186_addr = 6'h5;
  assign pht_1_1_MPORT_186_mask = 1'h1;
  assign pht_1_1_MPORT_186_en = reset;
  assign pht_1_1_MPORT_188_data = 1'h0;
  assign pht_1_1_MPORT_188_addr = 6'h6;
  assign pht_1_1_MPORT_188_mask = 1'h1;
  assign pht_1_1_MPORT_188_en = reset;
  assign pht_1_1_MPORT_190_data = 1'h0;
  assign pht_1_1_MPORT_190_addr = 6'h7;
  assign pht_1_1_MPORT_190_mask = 1'h1;
  assign pht_1_1_MPORT_190_en = reset;
  assign pht_1_1_MPORT_192_data = 1'h0;
  assign pht_1_1_MPORT_192_addr = 6'h8;
  assign pht_1_1_MPORT_192_mask = 1'h1;
  assign pht_1_1_MPORT_192_en = reset;
  assign pht_1_1_MPORT_194_data = 1'h0;
  assign pht_1_1_MPORT_194_addr = 6'h9;
  assign pht_1_1_MPORT_194_mask = 1'h1;
  assign pht_1_1_MPORT_194_en = reset;
  assign pht_1_1_MPORT_196_data = 1'h0;
  assign pht_1_1_MPORT_196_addr = 6'ha;
  assign pht_1_1_MPORT_196_mask = 1'h1;
  assign pht_1_1_MPORT_196_en = reset;
  assign pht_1_1_MPORT_198_data = 1'h0;
  assign pht_1_1_MPORT_198_addr = 6'hb;
  assign pht_1_1_MPORT_198_mask = 1'h1;
  assign pht_1_1_MPORT_198_en = reset;
  assign pht_1_1_MPORT_200_data = 1'h0;
  assign pht_1_1_MPORT_200_addr = 6'hc;
  assign pht_1_1_MPORT_200_mask = 1'h1;
  assign pht_1_1_MPORT_200_en = reset;
  assign pht_1_1_MPORT_202_data = 1'h0;
  assign pht_1_1_MPORT_202_addr = 6'hd;
  assign pht_1_1_MPORT_202_mask = 1'h1;
  assign pht_1_1_MPORT_202_en = reset;
  assign pht_1_1_MPORT_204_data = 1'h0;
  assign pht_1_1_MPORT_204_addr = 6'he;
  assign pht_1_1_MPORT_204_mask = 1'h1;
  assign pht_1_1_MPORT_204_en = reset;
  assign pht_1_1_MPORT_206_data = 1'h0;
  assign pht_1_1_MPORT_206_addr = 6'hf;
  assign pht_1_1_MPORT_206_mask = 1'h1;
  assign pht_1_1_MPORT_206_en = reset;
  assign pht_1_1_MPORT_208_data = 1'h0;
  assign pht_1_1_MPORT_208_addr = 6'h10;
  assign pht_1_1_MPORT_208_mask = 1'h1;
  assign pht_1_1_MPORT_208_en = reset;
  assign pht_1_1_MPORT_210_data = 1'h0;
  assign pht_1_1_MPORT_210_addr = 6'h11;
  assign pht_1_1_MPORT_210_mask = 1'h1;
  assign pht_1_1_MPORT_210_en = reset;
  assign pht_1_1_MPORT_212_data = 1'h0;
  assign pht_1_1_MPORT_212_addr = 6'h12;
  assign pht_1_1_MPORT_212_mask = 1'h1;
  assign pht_1_1_MPORT_212_en = reset;
  assign pht_1_1_MPORT_214_data = 1'h0;
  assign pht_1_1_MPORT_214_addr = 6'h13;
  assign pht_1_1_MPORT_214_mask = 1'h1;
  assign pht_1_1_MPORT_214_en = reset;
  assign pht_1_1_MPORT_216_data = 1'h0;
  assign pht_1_1_MPORT_216_addr = 6'h14;
  assign pht_1_1_MPORT_216_mask = 1'h1;
  assign pht_1_1_MPORT_216_en = reset;
  assign pht_1_1_MPORT_218_data = 1'h0;
  assign pht_1_1_MPORT_218_addr = 6'h15;
  assign pht_1_1_MPORT_218_mask = 1'h1;
  assign pht_1_1_MPORT_218_en = reset;
  assign pht_1_1_MPORT_220_data = 1'h0;
  assign pht_1_1_MPORT_220_addr = 6'h16;
  assign pht_1_1_MPORT_220_mask = 1'h1;
  assign pht_1_1_MPORT_220_en = reset;
  assign pht_1_1_MPORT_222_data = 1'h0;
  assign pht_1_1_MPORT_222_addr = 6'h17;
  assign pht_1_1_MPORT_222_mask = 1'h1;
  assign pht_1_1_MPORT_222_en = reset;
  assign pht_1_1_MPORT_224_data = 1'h0;
  assign pht_1_1_MPORT_224_addr = 6'h18;
  assign pht_1_1_MPORT_224_mask = 1'h1;
  assign pht_1_1_MPORT_224_en = reset;
  assign pht_1_1_MPORT_226_data = 1'h0;
  assign pht_1_1_MPORT_226_addr = 6'h19;
  assign pht_1_1_MPORT_226_mask = 1'h1;
  assign pht_1_1_MPORT_226_en = reset;
  assign pht_1_1_MPORT_228_data = 1'h0;
  assign pht_1_1_MPORT_228_addr = 6'h1a;
  assign pht_1_1_MPORT_228_mask = 1'h1;
  assign pht_1_1_MPORT_228_en = reset;
  assign pht_1_1_MPORT_230_data = 1'h0;
  assign pht_1_1_MPORT_230_addr = 6'h1b;
  assign pht_1_1_MPORT_230_mask = 1'h1;
  assign pht_1_1_MPORT_230_en = reset;
  assign pht_1_1_MPORT_232_data = 1'h0;
  assign pht_1_1_MPORT_232_addr = 6'h1c;
  assign pht_1_1_MPORT_232_mask = 1'h1;
  assign pht_1_1_MPORT_232_en = reset;
  assign pht_1_1_MPORT_234_data = 1'h0;
  assign pht_1_1_MPORT_234_addr = 6'h1d;
  assign pht_1_1_MPORT_234_mask = 1'h1;
  assign pht_1_1_MPORT_234_en = reset;
  assign pht_1_1_MPORT_236_data = 1'h0;
  assign pht_1_1_MPORT_236_addr = 6'h1e;
  assign pht_1_1_MPORT_236_mask = 1'h1;
  assign pht_1_1_MPORT_236_en = reset;
  assign pht_1_1_MPORT_238_data = 1'h0;
  assign pht_1_1_MPORT_238_addr = 6'h1f;
  assign pht_1_1_MPORT_238_mask = 1'h1;
  assign pht_1_1_MPORT_238_en = reset;
  assign pht_1_1_MPORT_240_data = 1'h0;
  assign pht_1_1_MPORT_240_addr = 6'h20;
  assign pht_1_1_MPORT_240_mask = 1'h1;
  assign pht_1_1_MPORT_240_en = reset;
  assign pht_1_1_MPORT_242_data = 1'h0;
  assign pht_1_1_MPORT_242_addr = 6'h21;
  assign pht_1_1_MPORT_242_mask = 1'h1;
  assign pht_1_1_MPORT_242_en = reset;
  assign pht_1_1_MPORT_244_data = 1'h0;
  assign pht_1_1_MPORT_244_addr = 6'h22;
  assign pht_1_1_MPORT_244_mask = 1'h1;
  assign pht_1_1_MPORT_244_en = reset;
  assign pht_1_1_MPORT_246_data = 1'h0;
  assign pht_1_1_MPORT_246_addr = 6'h23;
  assign pht_1_1_MPORT_246_mask = 1'h1;
  assign pht_1_1_MPORT_246_en = reset;
  assign pht_1_1_MPORT_248_data = 1'h0;
  assign pht_1_1_MPORT_248_addr = 6'h24;
  assign pht_1_1_MPORT_248_mask = 1'h1;
  assign pht_1_1_MPORT_248_en = reset;
  assign pht_1_1_MPORT_250_data = 1'h0;
  assign pht_1_1_MPORT_250_addr = 6'h25;
  assign pht_1_1_MPORT_250_mask = 1'h1;
  assign pht_1_1_MPORT_250_en = reset;
  assign pht_1_1_MPORT_252_data = 1'h0;
  assign pht_1_1_MPORT_252_addr = 6'h26;
  assign pht_1_1_MPORT_252_mask = 1'h1;
  assign pht_1_1_MPORT_252_en = reset;
  assign pht_1_1_MPORT_254_data = 1'h0;
  assign pht_1_1_MPORT_254_addr = 6'h27;
  assign pht_1_1_MPORT_254_mask = 1'h1;
  assign pht_1_1_MPORT_254_en = reset;
  assign pht_1_1_MPORT_256_data = 1'h0;
  assign pht_1_1_MPORT_256_addr = 6'h28;
  assign pht_1_1_MPORT_256_mask = 1'h1;
  assign pht_1_1_MPORT_256_en = reset;
  assign pht_1_1_MPORT_258_data = 1'h0;
  assign pht_1_1_MPORT_258_addr = 6'h29;
  assign pht_1_1_MPORT_258_mask = 1'h1;
  assign pht_1_1_MPORT_258_en = reset;
  assign pht_1_1_MPORT_260_data = 1'h0;
  assign pht_1_1_MPORT_260_addr = 6'h2a;
  assign pht_1_1_MPORT_260_mask = 1'h1;
  assign pht_1_1_MPORT_260_en = reset;
  assign pht_1_1_MPORT_262_data = 1'h0;
  assign pht_1_1_MPORT_262_addr = 6'h2b;
  assign pht_1_1_MPORT_262_mask = 1'h1;
  assign pht_1_1_MPORT_262_en = reset;
  assign pht_1_1_MPORT_264_data = 1'h0;
  assign pht_1_1_MPORT_264_addr = 6'h2c;
  assign pht_1_1_MPORT_264_mask = 1'h1;
  assign pht_1_1_MPORT_264_en = reset;
  assign pht_1_1_MPORT_266_data = 1'h0;
  assign pht_1_1_MPORT_266_addr = 6'h2d;
  assign pht_1_1_MPORT_266_mask = 1'h1;
  assign pht_1_1_MPORT_266_en = reset;
  assign pht_1_1_MPORT_268_data = 1'h0;
  assign pht_1_1_MPORT_268_addr = 6'h2e;
  assign pht_1_1_MPORT_268_mask = 1'h1;
  assign pht_1_1_MPORT_268_en = reset;
  assign pht_1_1_MPORT_270_data = 1'h0;
  assign pht_1_1_MPORT_270_addr = 6'h2f;
  assign pht_1_1_MPORT_270_mask = 1'h1;
  assign pht_1_1_MPORT_270_en = reset;
  assign pht_1_1_MPORT_272_data = 1'h0;
  assign pht_1_1_MPORT_272_addr = 6'h30;
  assign pht_1_1_MPORT_272_mask = 1'h1;
  assign pht_1_1_MPORT_272_en = reset;
  assign pht_1_1_MPORT_274_data = 1'h0;
  assign pht_1_1_MPORT_274_addr = 6'h31;
  assign pht_1_1_MPORT_274_mask = 1'h1;
  assign pht_1_1_MPORT_274_en = reset;
  assign pht_1_1_MPORT_276_data = 1'h0;
  assign pht_1_1_MPORT_276_addr = 6'h32;
  assign pht_1_1_MPORT_276_mask = 1'h1;
  assign pht_1_1_MPORT_276_en = reset;
  assign pht_1_1_MPORT_278_data = 1'h0;
  assign pht_1_1_MPORT_278_addr = 6'h33;
  assign pht_1_1_MPORT_278_mask = 1'h1;
  assign pht_1_1_MPORT_278_en = reset;
  assign pht_1_1_MPORT_280_data = 1'h0;
  assign pht_1_1_MPORT_280_addr = 6'h34;
  assign pht_1_1_MPORT_280_mask = 1'h1;
  assign pht_1_1_MPORT_280_en = reset;
  assign pht_1_1_MPORT_282_data = 1'h0;
  assign pht_1_1_MPORT_282_addr = 6'h35;
  assign pht_1_1_MPORT_282_mask = 1'h1;
  assign pht_1_1_MPORT_282_en = reset;
  assign pht_1_1_MPORT_284_data = 1'h0;
  assign pht_1_1_MPORT_284_addr = 6'h36;
  assign pht_1_1_MPORT_284_mask = 1'h1;
  assign pht_1_1_MPORT_284_en = reset;
  assign pht_1_1_MPORT_286_data = 1'h0;
  assign pht_1_1_MPORT_286_addr = 6'h37;
  assign pht_1_1_MPORT_286_mask = 1'h1;
  assign pht_1_1_MPORT_286_en = reset;
  assign pht_1_1_MPORT_288_data = 1'h0;
  assign pht_1_1_MPORT_288_addr = 6'h38;
  assign pht_1_1_MPORT_288_mask = 1'h1;
  assign pht_1_1_MPORT_288_en = reset;
  assign pht_1_1_MPORT_290_data = 1'h0;
  assign pht_1_1_MPORT_290_addr = 6'h39;
  assign pht_1_1_MPORT_290_mask = 1'h1;
  assign pht_1_1_MPORT_290_en = reset;
  assign pht_1_1_MPORT_292_data = 1'h0;
  assign pht_1_1_MPORT_292_addr = 6'h3a;
  assign pht_1_1_MPORT_292_mask = 1'h1;
  assign pht_1_1_MPORT_292_en = reset;
  assign pht_1_1_MPORT_294_data = 1'h0;
  assign pht_1_1_MPORT_294_addr = 6'h3b;
  assign pht_1_1_MPORT_294_mask = 1'h1;
  assign pht_1_1_MPORT_294_en = reset;
  assign pht_1_1_MPORT_296_data = 1'h0;
  assign pht_1_1_MPORT_296_addr = 6'h3c;
  assign pht_1_1_MPORT_296_mask = 1'h1;
  assign pht_1_1_MPORT_296_en = reset;
  assign pht_1_1_MPORT_298_data = 1'h0;
  assign pht_1_1_MPORT_298_addr = 6'h3d;
  assign pht_1_1_MPORT_298_mask = 1'h1;
  assign pht_1_1_MPORT_298_en = reset;
  assign pht_1_1_MPORT_300_data = 1'h0;
  assign pht_1_1_MPORT_300_addr = 6'h3e;
  assign pht_1_1_MPORT_300_mask = 1'h1;
  assign pht_1_1_MPORT_300_en = reset;
  assign pht_1_1_MPORT_302_data = 1'h0;
  assign pht_1_1_MPORT_302_addr = 6'h3f;
  assign pht_1_1_MPORT_302_mask = 1'h1;
  assign pht_1_1_MPORT_302_en = reset;
//   assign pht_1_2_MPORT_2_en = pht_1_2_MPORT_2_en_pipe_0;
  assign pht_1_2_MPORT_2_addr = pht_1_2_MPORT_2_addr_pipe_0;
  assign pht_1_2_MPORT_2_data = pht_1_2[pht_1_2_MPORT_2_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_2_MPORT_10_en = pht_1_2_MPORT_10_en_pipe_0;
  assign pht_1_2_MPORT_10_addr = pht_1_2_MPORT_10_addr_pipe_0;
  assign pht_1_2_MPORT_10_data = pht_1_2[pht_1_2_MPORT_10_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_2_MPORT_20_en = pht_1_2_MPORT_20_en_pipe_0;
  assign pht_1_2_MPORT_20_addr = pht_1_2_MPORT_20_addr_pipe_0;
  assign pht_1_2_MPORT_20_data = pht_1_2[pht_1_2_MPORT_20_addr]; // @[PatternHistoryTable.scala 21:28]
  assign pht_1_2_MPORT_36_data = pht_wdata_w[1];
  assign pht_1_2_MPORT_36_addr = REG_37;
  assign pht_1_2_MPORT_36_mask = 1'h1;
  assign pht_1_2_MPORT_36_en = REG_29 & REG_36;
  assign pht_1_2_MPORT_304_data = 1'h0;
  assign pht_1_2_MPORT_304_addr = 6'h0;
  assign pht_1_2_MPORT_304_mask = 1'h1;
  assign pht_1_2_MPORT_304_en = reset;
  assign pht_1_2_MPORT_306_data = 1'h0;
  assign pht_1_2_MPORT_306_addr = 6'h1;
  assign pht_1_2_MPORT_306_mask = 1'h1;
  assign pht_1_2_MPORT_306_en = reset;
  assign pht_1_2_MPORT_308_data = 1'h0;
  assign pht_1_2_MPORT_308_addr = 6'h2;
  assign pht_1_2_MPORT_308_mask = 1'h1;
  assign pht_1_2_MPORT_308_en = reset;
  assign pht_1_2_MPORT_310_data = 1'h0;
  assign pht_1_2_MPORT_310_addr = 6'h3;
  assign pht_1_2_MPORT_310_mask = 1'h1;
  assign pht_1_2_MPORT_310_en = reset;
  assign pht_1_2_MPORT_312_data = 1'h0;
  assign pht_1_2_MPORT_312_addr = 6'h4;
  assign pht_1_2_MPORT_312_mask = 1'h1;
  assign pht_1_2_MPORT_312_en = reset;
  assign pht_1_2_MPORT_314_data = 1'h0;
  assign pht_1_2_MPORT_314_addr = 6'h5;
  assign pht_1_2_MPORT_314_mask = 1'h1;
  assign pht_1_2_MPORT_314_en = reset;
  assign pht_1_2_MPORT_316_data = 1'h0;
  assign pht_1_2_MPORT_316_addr = 6'h6;
  assign pht_1_2_MPORT_316_mask = 1'h1;
  assign pht_1_2_MPORT_316_en = reset;
  assign pht_1_2_MPORT_318_data = 1'h0;
  assign pht_1_2_MPORT_318_addr = 6'h7;
  assign pht_1_2_MPORT_318_mask = 1'h1;
  assign pht_1_2_MPORT_318_en = reset;
  assign pht_1_2_MPORT_320_data = 1'h0;
  assign pht_1_2_MPORT_320_addr = 6'h8;
  assign pht_1_2_MPORT_320_mask = 1'h1;
  assign pht_1_2_MPORT_320_en = reset;
  assign pht_1_2_MPORT_322_data = 1'h0;
  assign pht_1_2_MPORT_322_addr = 6'h9;
  assign pht_1_2_MPORT_322_mask = 1'h1;
  assign pht_1_2_MPORT_322_en = reset;
  assign pht_1_2_MPORT_324_data = 1'h0;
  assign pht_1_2_MPORT_324_addr = 6'ha;
  assign pht_1_2_MPORT_324_mask = 1'h1;
  assign pht_1_2_MPORT_324_en = reset;
  assign pht_1_2_MPORT_326_data = 1'h0;
  assign pht_1_2_MPORT_326_addr = 6'hb;
  assign pht_1_2_MPORT_326_mask = 1'h1;
  assign pht_1_2_MPORT_326_en = reset;
  assign pht_1_2_MPORT_328_data = 1'h0;
  assign pht_1_2_MPORT_328_addr = 6'hc;
  assign pht_1_2_MPORT_328_mask = 1'h1;
  assign pht_1_2_MPORT_328_en = reset;
  assign pht_1_2_MPORT_330_data = 1'h0;
  assign pht_1_2_MPORT_330_addr = 6'hd;
  assign pht_1_2_MPORT_330_mask = 1'h1;
  assign pht_1_2_MPORT_330_en = reset;
  assign pht_1_2_MPORT_332_data = 1'h0;
  assign pht_1_2_MPORT_332_addr = 6'he;
  assign pht_1_2_MPORT_332_mask = 1'h1;
  assign pht_1_2_MPORT_332_en = reset;
  assign pht_1_2_MPORT_334_data = 1'h0;
  assign pht_1_2_MPORT_334_addr = 6'hf;
  assign pht_1_2_MPORT_334_mask = 1'h1;
  assign pht_1_2_MPORT_334_en = reset;
  assign pht_1_2_MPORT_336_data = 1'h0;
  assign pht_1_2_MPORT_336_addr = 6'h10;
  assign pht_1_2_MPORT_336_mask = 1'h1;
  assign pht_1_2_MPORT_336_en = reset;
  assign pht_1_2_MPORT_338_data = 1'h0;
  assign pht_1_2_MPORT_338_addr = 6'h11;
  assign pht_1_2_MPORT_338_mask = 1'h1;
  assign pht_1_2_MPORT_338_en = reset;
  assign pht_1_2_MPORT_340_data = 1'h0;
  assign pht_1_2_MPORT_340_addr = 6'h12;
  assign pht_1_2_MPORT_340_mask = 1'h1;
  assign pht_1_2_MPORT_340_en = reset;
  assign pht_1_2_MPORT_342_data = 1'h0;
  assign pht_1_2_MPORT_342_addr = 6'h13;
  assign pht_1_2_MPORT_342_mask = 1'h1;
  assign pht_1_2_MPORT_342_en = reset;
  assign pht_1_2_MPORT_344_data = 1'h0;
  assign pht_1_2_MPORT_344_addr = 6'h14;
  assign pht_1_2_MPORT_344_mask = 1'h1;
  assign pht_1_2_MPORT_344_en = reset;
  assign pht_1_2_MPORT_346_data = 1'h0;
  assign pht_1_2_MPORT_346_addr = 6'h15;
  assign pht_1_2_MPORT_346_mask = 1'h1;
  assign pht_1_2_MPORT_346_en = reset;
  assign pht_1_2_MPORT_348_data = 1'h0;
  assign pht_1_2_MPORT_348_addr = 6'h16;
  assign pht_1_2_MPORT_348_mask = 1'h1;
  assign pht_1_2_MPORT_348_en = reset;
  assign pht_1_2_MPORT_350_data = 1'h0;
  assign pht_1_2_MPORT_350_addr = 6'h17;
  assign pht_1_2_MPORT_350_mask = 1'h1;
  assign pht_1_2_MPORT_350_en = reset;
  assign pht_1_2_MPORT_352_data = 1'h0;
  assign pht_1_2_MPORT_352_addr = 6'h18;
  assign pht_1_2_MPORT_352_mask = 1'h1;
  assign pht_1_2_MPORT_352_en = reset;
  assign pht_1_2_MPORT_354_data = 1'h0;
  assign pht_1_2_MPORT_354_addr = 6'h19;
  assign pht_1_2_MPORT_354_mask = 1'h1;
  assign pht_1_2_MPORT_354_en = reset;
  assign pht_1_2_MPORT_356_data = 1'h0;
  assign pht_1_2_MPORT_356_addr = 6'h1a;
  assign pht_1_2_MPORT_356_mask = 1'h1;
  assign pht_1_2_MPORT_356_en = reset;
  assign pht_1_2_MPORT_358_data = 1'h0;
  assign pht_1_2_MPORT_358_addr = 6'h1b;
  assign pht_1_2_MPORT_358_mask = 1'h1;
  assign pht_1_2_MPORT_358_en = reset;
  assign pht_1_2_MPORT_360_data = 1'h0;
  assign pht_1_2_MPORT_360_addr = 6'h1c;
  assign pht_1_2_MPORT_360_mask = 1'h1;
  assign pht_1_2_MPORT_360_en = reset;
  assign pht_1_2_MPORT_362_data = 1'h0;
  assign pht_1_2_MPORT_362_addr = 6'h1d;
  assign pht_1_2_MPORT_362_mask = 1'h1;
  assign pht_1_2_MPORT_362_en = reset;
  assign pht_1_2_MPORT_364_data = 1'h0;
  assign pht_1_2_MPORT_364_addr = 6'h1e;
  assign pht_1_2_MPORT_364_mask = 1'h1;
  assign pht_1_2_MPORT_364_en = reset;
  assign pht_1_2_MPORT_366_data = 1'h0;
  assign pht_1_2_MPORT_366_addr = 6'h1f;
  assign pht_1_2_MPORT_366_mask = 1'h1;
  assign pht_1_2_MPORT_366_en = reset;
  assign pht_1_2_MPORT_368_data = 1'h0;
  assign pht_1_2_MPORT_368_addr = 6'h20;
  assign pht_1_2_MPORT_368_mask = 1'h1;
  assign pht_1_2_MPORT_368_en = reset;
  assign pht_1_2_MPORT_370_data = 1'h0;
  assign pht_1_2_MPORT_370_addr = 6'h21;
  assign pht_1_2_MPORT_370_mask = 1'h1;
  assign pht_1_2_MPORT_370_en = reset;
  assign pht_1_2_MPORT_372_data = 1'h0;
  assign pht_1_2_MPORT_372_addr = 6'h22;
  assign pht_1_2_MPORT_372_mask = 1'h1;
  assign pht_1_2_MPORT_372_en = reset;
  assign pht_1_2_MPORT_374_data = 1'h0;
  assign pht_1_2_MPORT_374_addr = 6'h23;
  assign pht_1_2_MPORT_374_mask = 1'h1;
  assign pht_1_2_MPORT_374_en = reset;
  assign pht_1_2_MPORT_376_data = 1'h0;
  assign pht_1_2_MPORT_376_addr = 6'h24;
  assign pht_1_2_MPORT_376_mask = 1'h1;
  assign pht_1_2_MPORT_376_en = reset;
  assign pht_1_2_MPORT_378_data = 1'h0;
  assign pht_1_2_MPORT_378_addr = 6'h25;
  assign pht_1_2_MPORT_378_mask = 1'h1;
  assign pht_1_2_MPORT_378_en = reset;
  assign pht_1_2_MPORT_380_data = 1'h0;
  assign pht_1_2_MPORT_380_addr = 6'h26;
  assign pht_1_2_MPORT_380_mask = 1'h1;
  assign pht_1_2_MPORT_380_en = reset;
  assign pht_1_2_MPORT_382_data = 1'h0;
  assign pht_1_2_MPORT_382_addr = 6'h27;
  assign pht_1_2_MPORT_382_mask = 1'h1;
  assign pht_1_2_MPORT_382_en = reset;
  assign pht_1_2_MPORT_384_data = 1'h0;
  assign pht_1_2_MPORT_384_addr = 6'h28;
  assign pht_1_2_MPORT_384_mask = 1'h1;
  assign pht_1_2_MPORT_384_en = reset;
  assign pht_1_2_MPORT_386_data = 1'h0;
  assign pht_1_2_MPORT_386_addr = 6'h29;
  assign pht_1_2_MPORT_386_mask = 1'h1;
  assign pht_1_2_MPORT_386_en = reset;
  assign pht_1_2_MPORT_388_data = 1'h0;
  assign pht_1_2_MPORT_388_addr = 6'h2a;
  assign pht_1_2_MPORT_388_mask = 1'h1;
  assign pht_1_2_MPORT_388_en = reset;
  assign pht_1_2_MPORT_390_data = 1'h0;
  assign pht_1_2_MPORT_390_addr = 6'h2b;
  assign pht_1_2_MPORT_390_mask = 1'h1;
  assign pht_1_2_MPORT_390_en = reset;
  assign pht_1_2_MPORT_392_data = 1'h0;
  assign pht_1_2_MPORT_392_addr = 6'h2c;
  assign pht_1_2_MPORT_392_mask = 1'h1;
  assign pht_1_2_MPORT_392_en = reset;
  assign pht_1_2_MPORT_394_data = 1'h0;
  assign pht_1_2_MPORT_394_addr = 6'h2d;
  assign pht_1_2_MPORT_394_mask = 1'h1;
  assign pht_1_2_MPORT_394_en = reset;
  assign pht_1_2_MPORT_396_data = 1'h0;
  assign pht_1_2_MPORT_396_addr = 6'h2e;
  assign pht_1_2_MPORT_396_mask = 1'h1;
  assign pht_1_2_MPORT_396_en = reset;
  assign pht_1_2_MPORT_398_data = 1'h0;
  assign pht_1_2_MPORT_398_addr = 6'h2f;
  assign pht_1_2_MPORT_398_mask = 1'h1;
  assign pht_1_2_MPORT_398_en = reset;
  assign pht_1_2_MPORT_400_data = 1'h0;
  assign pht_1_2_MPORT_400_addr = 6'h30;
  assign pht_1_2_MPORT_400_mask = 1'h1;
  assign pht_1_2_MPORT_400_en = reset;
  assign pht_1_2_MPORT_402_data = 1'h0;
  assign pht_1_2_MPORT_402_addr = 6'h31;
  assign pht_1_2_MPORT_402_mask = 1'h1;
  assign pht_1_2_MPORT_402_en = reset;
  assign pht_1_2_MPORT_404_data = 1'h0;
  assign pht_1_2_MPORT_404_addr = 6'h32;
  assign pht_1_2_MPORT_404_mask = 1'h1;
  assign pht_1_2_MPORT_404_en = reset;
  assign pht_1_2_MPORT_406_data = 1'h0;
  assign pht_1_2_MPORT_406_addr = 6'h33;
  assign pht_1_2_MPORT_406_mask = 1'h1;
  assign pht_1_2_MPORT_406_en = reset;
  assign pht_1_2_MPORT_408_data = 1'h0;
  assign pht_1_2_MPORT_408_addr = 6'h34;
  assign pht_1_2_MPORT_408_mask = 1'h1;
  assign pht_1_2_MPORT_408_en = reset;
  assign pht_1_2_MPORT_410_data = 1'h0;
  assign pht_1_2_MPORT_410_addr = 6'h35;
  assign pht_1_2_MPORT_410_mask = 1'h1;
  assign pht_1_2_MPORT_410_en = reset;
  assign pht_1_2_MPORT_412_data = 1'h0;
  assign pht_1_2_MPORT_412_addr = 6'h36;
  assign pht_1_2_MPORT_412_mask = 1'h1;
  assign pht_1_2_MPORT_412_en = reset;
  assign pht_1_2_MPORT_414_data = 1'h0;
  assign pht_1_2_MPORT_414_addr = 6'h37;
  assign pht_1_2_MPORT_414_mask = 1'h1;
  assign pht_1_2_MPORT_414_en = reset;
  assign pht_1_2_MPORT_416_data = 1'h0;
  assign pht_1_2_MPORT_416_addr = 6'h38;
  assign pht_1_2_MPORT_416_mask = 1'h1;
  assign pht_1_2_MPORT_416_en = reset;
  assign pht_1_2_MPORT_418_data = 1'h0;
  assign pht_1_2_MPORT_418_addr = 6'h39;
  assign pht_1_2_MPORT_418_mask = 1'h1;
  assign pht_1_2_MPORT_418_en = reset;
  assign pht_1_2_MPORT_420_data = 1'h0;
  assign pht_1_2_MPORT_420_addr = 6'h3a;
  assign pht_1_2_MPORT_420_mask = 1'h1;
  assign pht_1_2_MPORT_420_en = reset;
  assign pht_1_2_MPORT_422_data = 1'h0;
  assign pht_1_2_MPORT_422_addr = 6'h3b;
  assign pht_1_2_MPORT_422_mask = 1'h1;
  assign pht_1_2_MPORT_422_en = reset;
  assign pht_1_2_MPORT_424_data = 1'h0;
  assign pht_1_2_MPORT_424_addr = 6'h3c;
  assign pht_1_2_MPORT_424_mask = 1'h1;
  assign pht_1_2_MPORT_424_en = reset;
  assign pht_1_2_MPORT_426_data = 1'h0;
  assign pht_1_2_MPORT_426_addr = 6'h3d;
  assign pht_1_2_MPORT_426_mask = 1'h1;
  assign pht_1_2_MPORT_426_en = reset;
  assign pht_1_2_MPORT_428_data = 1'h0;
  assign pht_1_2_MPORT_428_addr = 6'h3e;
  assign pht_1_2_MPORT_428_mask = 1'h1;
  assign pht_1_2_MPORT_428_en = reset;
  assign pht_1_2_MPORT_430_data = 1'h0;
  assign pht_1_2_MPORT_430_addr = 6'h3f;
  assign pht_1_2_MPORT_430_mask = 1'h1;
  assign pht_1_2_MPORT_430_en = reset;
//   assign pht_1_3_MPORT_3_en = pht_1_3_MPORT_3_en_pipe_0;
  assign pht_1_3_MPORT_3_addr = pht_1_3_MPORT_3_addr_pipe_0;
  assign pht_1_3_MPORT_3_data = pht_1_3[pht_1_3_MPORT_3_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_3_MPORT_11_en = pht_1_3_MPORT_11_en_pipe_0;
  assign pht_1_3_MPORT_11_addr = pht_1_3_MPORT_11_addr_pipe_0;
  assign pht_1_3_MPORT_11_data = pht_1_3[pht_1_3_MPORT_11_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_3_MPORT_22_en = pht_1_3_MPORT_22_en_pipe_0;
  assign pht_1_3_MPORT_22_addr = pht_1_3_MPORT_22_addr_pipe_0;
  assign pht_1_3_MPORT_22_data = pht_1_3[pht_1_3_MPORT_22_addr]; // @[PatternHistoryTable.scala 21:28]
  assign pht_1_3_MPORT_38_data = pht_wdata_w[1];
  assign pht_1_3_MPORT_38_addr = REG_40;
  assign pht_1_3_MPORT_38_mask = 1'h1;
  assign pht_1_3_MPORT_38_en = REG_29 & REG_39;
  assign pht_1_3_MPORT_432_data = 1'h0;
  assign pht_1_3_MPORT_432_addr = 6'h0;
  assign pht_1_3_MPORT_432_mask = 1'h1;
  assign pht_1_3_MPORT_432_en = reset;
  assign pht_1_3_MPORT_434_data = 1'h0;
  assign pht_1_3_MPORT_434_addr = 6'h1;
  assign pht_1_3_MPORT_434_mask = 1'h1;
  assign pht_1_3_MPORT_434_en = reset;
  assign pht_1_3_MPORT_436_data = 1'h0;
  assign pht_1_3_MPORT_436_addr = 6'h2;
  assign pht_1_3_MPORT_436_mask = 1'h1;
  assign pht_1_3_MPORT_436_en = reset;
  assign pht_1_3_MPORT_438_data = 1'h0;
  assign pht_1_3_MPORT_438_addr = 6'h3;
  assign pht_1_3_MPORT_438_mask = 1'h1;
  assign pht_1_3_MPORT_438_en = reset;
  assign pht_1_3_MPORT_440_data = 1'h0;
  assign pht_1_3_MPORT_440_addr = 6'h4;
  assign pht_1_3_MPORT_440_mask = 1'h1;
  assign pht_1_3_MPORT_440_en = reset;
  assign pht_1_3_MPORT_442_data = 1'h0;
  assign pht_1_3_MPORT_442_addr = 6'h5;
  assign pht_1_3_MPORT_442_mask = 1'h1;
  assign pht_1_3_MPORT_442_en = reset;
  assign pht_1_3_MPORT_444_data = 1'h0;
  assign pht_1_3_MPORT_444_addr = 6'h6;
  assign pht_1_3_MPORT_444_mask = 1'h1;
  assign pht_1_3_MPORT_444_en = reset;
  assign pht_1_3_MPORT_446_data = 1'h0;
  assign pht_1_3_MPORT_446_addr = 6'h7;
  assign pht_1_3_MPORT_446_mask = 1'h1;
  assign pht_1_3_MPORT_446_en = reset;
  assign pht_1_3_MPORT_448_data = 1'h0;
  assign pht_1_3_MPORT_448_addr = 6'h8;
  assign pht_1_3_MPORT_448_mask = 1'h1;
  assign pht_1_3_MPORT_448_en = reset;
  assign pht_1_3_MPORT_450_data = 1'h0;
  assign pht_1_3_MPORT_450_addr = 6'h9;
  assign pht_1_3_MPORT_450_mask = 1'h1;
  assign pht_1_3_MPORT_450_en = reset;
  assign pht_1_3_MPORT_452_data = 1'h0;
  assign pht_1_3_MPORT_452_addr = 6'ha;
  assign pht_1_3_MPORT_452_mask = 1'h1;
  assign pht_1_3_MPORT_452_en = reset;
  assign pht_1_3_MPORT_454_data = 1'h0;
  assign pht_1_3_MPORT_454_addr = 6'hb;
  assign pht_1_3_MPORT_454_mask = 1'h1;
  assign pht_1_3_MPORT_454_en = reset;
  assign pht_1_3_MPORT_456_data = 1'h0;
  assign pht_1_3_MPORT_456_addr = 6'hc;
  assign pht_1_3_MPORT_456_mask = 1'h1;
  assign pht_1_3_MPORT_456_en = reset;
  assign pht_1_3_MPORT_458_data = 1'h0;
  assign pht_1_3_MPORT_458_addr = 6'hd;
  assign pht_1_3_MPORT_458_mask = 1'h1;
  assign pht_1_3_MPORT_458_en = reset;
  assign pht_1_3_MPORT_460_data = 1'h0;
  assign pht_1_3_MPORT_460_addr = 6'he;
  assign pht_1_3_MPORT_460_mask = 1'h1;
  assign pht_1_3_MPORT_460_en = reset;
  assign pht_1_3_MPORT_462_data = 1'h0;
  assign pht_1_3_MPORT_462_addr = 6'hf;
  assign pht_1_3_MPORT_462_mask = 1'h1;
  assign pht_1_3_MPORT_462_en = reset;
  assign pht_1_3_MPORT_464_data = 1'h0;
  assign pht_1_3_MPORT_464_addr = 6'h10;
  assign pht_1_3_MPORT_464_mask = 1'h1;
  assign pht_1_3_MPORT_464_en = reset;
  assign pht_1_3_MPORT_466_data = 1'h0;
  assign pht_1_3_MPORT_466_addr = 6'h11;
  assign pht_1_3_MPORT_466_mask = 1'h1;
  assign pht_1_3_MPORT_466_en = reset;
  assign pht_1_3_MPORT_468_data = 1'h0;
  assign pht_1_3_MPORT_468_addr = 6'h12;
  assign pht_1_3_MPORT_468_mask = 1'h1;
  assign pht_1_3_MPORT_468_en = reset;
  assign pht_1_3_MPORT_470_data = 1'h0;
  assign pht_1_3_MPORT_470_addr = 6'h13;
  assign pht_1_3_MPORT_470_mask = 1'h1;
  assign pht_1_3_MPORT_470_en = reset;
  assign pht_1_3_MPORT_472_data = 1'h0;
  assign pht_1_3_MPORT_472_addr = 6'h14;
  assign pht_1_3_MPORT_472_mask = 1'h1;
  assign pht_1_3_MPORT_472_en = reset;
  assign pht_1_3_MPORT_474_data = 1'h0;
  assign pht_1_3_MPORT_474_addr = 6'h15;
  assign pht_1_3_MPORT_474_mask = 1'h1;
  assign pht_1_3_MPORT_474_en = reset;
  assign pht_1_3_MPORT_476_data = 1'h0;
  assign pht_1_3_MPORT_476_addr = 6'h16;
  assign pht_1_3_MPORT_476_mask = 1'h1;
  assign pht_1_3_MPORT_476_en = reset;
  assign pht_1_3_MPORT_478_data = 1'h0;
  assign pht_1_3_MPORT_478_addr = 6'h17;
  assign pht_1_3_MPORT_478_mask = 1'h1;
  assign pht_1_3_MPORT_478_en = reset;
  assign pht_1_3_MPORT_480_data = 1'h0;
  assign pht_1_3_MPORT_480_addr = 6'h18;
  assign pht_1_3_MPORT_480_mask = 1'h1;
  assign pht_1_3_MPORT_480_en = reset;
  assign pht_1_3_MPORT_482_data = 1'h0;
  assign pht_1_3_MPORT_482_addr = 6'h19;
  assign pht_1_3_MPORT_482_mask = 1'h1;
  assign pht_1_3_MPORT_482_en = reset;
  assign pht_1_3_MPORT_484_data = 1'h0;
  assign pht_1_3_MPORT_484_addr = 6'h1a;
  assign pht_1_3_MPORT_484_mask = 1'h1;
  assign pht_1_3_MPORT_484_en = reset;
  assign pht_1_3_MPORT_486_data = 1'h0;
  assign pht_1_3_MPORT_486_addr = 6'h1b;
  assign pht_1_3_MPORT_486_mask = 1'h1;
  assign pht_1_3_MPORT_486_en = reset;
  assign pht_1_3_MPORT_488_data = 1'h0;
  assign pht_1_3_MPORT_488_addr = 6'h1c;
  assign pht_1_3_MPORT_488_mask = 1'h1;
  assign pht_1_3_MPORT_488_en = reset;
  assign pht_1_3_MPORT_490_data = 1'h0;
  assign pht_1_3_MPORT_490_addr = 6'h1d;
  assign pht_1_3_MPORT_490_mask = 1'h1;
  assign pht_1_3_MPORT_490_en = reset;
  assign pht_1_3_MPORT_492_data = 1'h0;
  assign pht_1_3_MPORT_492_addr = 6'h1e;
  assign pht_1_3_MPORT_492_mask = 1'h1;
  assign pht_1_3_MPORT_492_en = reset;
  assign pht_1_3_MPORT_494_data = 1'h0;
  assign pht_1_3_MPORT_494_addr = 6'h1f;
  assign pht_1_3_MPORT_494_mask = 1'h1;
  assign pht_1_3_MPORT_494_en = reset;
  assign pht_1_3_MPORT_496_data = 1'h0;
  assign pht_1_3_MPORT_496_addr = 6'h20;
  assign pht_1_3_MPORT_496_mask = 1'h1;
  assign pht_1_3_MPORT_496_en = reset;
  assign pht_1_3_MPORT_498_data = 1'h0;
  assign pht_1_3_MPORT_498_addr = 6'h21;
  assign pht_1_3_MPORT_498_mask = 1'h1;
  assign pht_1_3_MPORT_498_en = reset;
  assign pht_1_3_MPORT_500_data = 1'h0;
  assign pht_1_3_MPORT_500_addr = 6'h22;
  assign pht_1_3_MPORT_500_mask = 1'h1;
  assign pht_1_3_MPORT_500_en = reset;
  assign pht_1_3_MPORT_502_data = 1'h0;
  assign pht_1_3_MPORT_502_addr = 6'h23;
  assign pht_1_3_MPORT_502_mask = 1'h1;
  assign pht_1_3_MPORT_502_en = reset;
  assign pht_1_3_MPORT_504_data = 1'h0;
  assign pht_1_3_MPORT_504_addr = 6'h24;
  assign pht_1_3_MPORT_504_mask = 1'h1;
  assign pht_1_3_MPORT_504_en = reset;
  assign pht_1_3_MPORT_506_data = 1'h0;
  assign pht_1_3_MPORT_506_addr = 6'h25;
  assign pht_1_3_MPORT_506_mask = 1'h1;
  assign pht_1_3_MPORT_506_en = reset;
  assign pht_1_3_MPORT_508_data = 1'h0;
  assign pht_1_3_MPORT_508_addr = 6'h26;
  assign pht_1_3_MPORT_508_mask = 1'h1;
  assign pht_1_3_MPORT_508_en = reset;
  assign pht_1_3_MPORT_510_data = 1'h0;
  assign pht_1_3_MPORT_510_addr = 6'h27;
  assign pht_1_3_MPORT_510_mask = 1'h1;
  assign pht_1_3_MPORT_510_en = reset;
  assign pht_1_3_MPORT_512_data = 1'h0;
  assign pht_1_3_MPORT_512_addr = 6'h28;
  assign pht_1_3_MPORT_512_mask = 1'h1;
  assign pht_1_3_MPORT_512_en = reset;
  assign pht_1_3_MPORT_514_data = 1'h0;
  assign pht_1_3_MPORT_514_addr = 6'h29;
  assign pht_1_3_MPORT_514_mask = 1'h1;
  assign pht_1_3_MPORT_514_en = reset;
  assign pht_1_3_MPORT_516_data = 1'h0;
  assign pht_1_3_MPORT_516_addr = 6'h2a;
  assign pht_1_3_MPORT_516_mask = 1'h1;
  assign pht_1_3_MPORT_516_en = reset;
  assign pht_1_3_MPORT_518_data = 1'h0;
  assign pht_1_3_MPORT_518_addr = 6'h2b;
  assign pht_1_3_MPORT_518_mask = 1'h1;
  assign pht_1_3_MPORT_518_en = reset;
  assign pht_1_3_MPORT_520_data = 1'h0;
  assign pht_1_3_MPORT_520_addr = 6'h2c;
  assign pht_1_3_MPORT_520_mask = 1'h1;
  assign pht_1_3_MPORT_520_en = reset;
  assign pht_1_3_MPORT_522_data = 1'h0;
  assign pht_1_3_MPORT_522_addr = 6'h2d;
  assign pht_1_3_MPORT_522_mask = 1'h1;
  assign pht_1_3_MPORT_522_en = reset;
  assign pht_1_3_MPORT_524_data = 1'h0;
  assign pht_1_3_MPORT_524_addr = 6'h2e;
  assign pht_1_3_MPORT_524_mask = 1'h1;
  assign pht_1_3_MPORT_524_en = reset;
  assign pht_1_3_MPORT_526_data = 1'h0;
  assign pht_1_3_MPORT_526_addr = 6'h2f;
  assign pht_1_3_MPORT_526_mask = 1'h1;
  assign pht_1_3_MPORT_526_en = reset;
  assign pht_1_3_MPORT_528_data = 1'h0;
  assign pht_1_3_MPORT_528_addr = 6'h30;
  assign pht_1_3_MPORT_528_mask = 1'h1;
  assign pht_1_3_MPORT_528_en = reset;
  assign pht_1_3_MPORT_530_data = 1'h0;
  assign pht_1_3_MPORT_530_addr = 6'h31;
  assign pht_1_3_MPORT_530_mask = 1'h1;
  assign pht_1_3_MPORT_530_en = reset;
  assign pht_1_3_MPORT_532_data = 1'h0;
  assign pht_1_3_MPORT_532_addr = 6'h32;
  assign pht_1_3_MPORT_532_mask = 1'h1;
  assign pht_1_3_MPORT_532_en = reset;
  assign pht_1_3_MPORT_534_data = 1'h0;
  assign pht_1_3_MPORT_534_addr = 6'h33;
  assign pht_1_3_MPORT_534_mask = 1'h1;
  assign pht_1_3_MPORT_534_en = reset;
  assign pht_1_3_MPORT_536_data = 1'h0;
  assign pht_1_3_MPORT_536_addr = 6'h34;
  assign pht_1_3_MPORT_536_mask = 1'h1;
  assign pht_1_3_MPORT_536_en = reset;
  assign pht_1_3_MPORT_538_data = 1'h0;
  assign pht_1_3_MPORT_538_addr = 6'h35;
  assign pht_1_3_MPORT_538_mask = 1'h1;
  assign pht_1_3_MPORT_538_en = reset;
  assign pht_1_3_MPORT_540_data = 1'h0;
  assign pht_1_3_MPORT_540_addr = 6'h36;
  assign pht_1_3_MPORT_540_mask = 1'h1;
  assign pht_1_3_MPORT_540_en = reset;
  assign pht_1_3_MPORT_542_data = 1'h0;
  assign pht_1_3_MPORT_542_addr = 6'h37;
  assign pht_1_3_MPORT_542_mask = 1'h1;
  assign pht_1_3_MPORT_542_en = reset;
  assign pht_1_3_MPORT_544_data = 1'h0;
  assign pht_1_3_MPORT_544_addr = 6'h38;
  assign pht_1_3_MPORT_544_mask = 1'h1;
  assign pht_1_3_MPORT_544_en = reset;
  assign pht_1_3_MPORT_546_data = 1'h0;
  assign pht_1_3_MPORT_546_addr = 6'h39;
  assign pht_1_3_MPORT_546_mask = 1'h1;
  assign pht_1_3_MPORT_546_en = reset;
  assign pht_1_3_MPORT_548_data = 1'h0;
  assign pht_1_3_MPORT_548_addr = 6'h3a;
  assign pht_1_3_MPORT_548_mask = 1'h1;
  assign pht_1_3_MPORT_548_en = reset;
  assign pht_1_3_MPORT_550_data = 1'h0;
  assign pht_1_3_MPORT_550_addr = 6'h3b;
  assign pht_1_3_MPORT_550_mask = 1'h1;
  assign pht_1_3_MPORT_550_en = reset;
  assign pht_1_3_MPORT_552_data = 1'h0;
  assign pht_1_3_MPORT_552_addr = 6'h3c;
  assign pht_1_3_MPORT_552_mask = 1'h1;
  assign pht_1_3_MPORT_552_en = reset;
  assign pht_1_3_MPORT_554_data = 1'h0;
  assign pht_1_3_MPORT_554_addr = 6'h3d;
  assign pht_1_3_MPORT_554_mask = 1'h1;
  assign pht_1_3_MPORT_554_en = reset;
  assign pht_1_3_MPORT_556_data = 1'h0;
  assign pht_1_3_MPORT_556_addr = 6'h3e;
  assign pht_1_3_MPORT_556_mask = 1'h1;
  assign pht_1_3_MPORT_556_en = reset;
  assign pht_1_3_MPORT_558_data = 1'h0;
  assign pht_1_3_MPORT_558_addr = 6'h3f;
  assign pht_1_3_MPORT_558_mask = 1'h1;
  assign pht_1_3_MPORT_558_en = reset;
//   assign pht_1_4_MPORT_4_en = pht_1_4_MPORT_4_en_pipe_0;
  assign pht_1_4_MPORT_4_addr = pht_1_4_MPORT_4_addr_pipe_0;
  assign pht_1_4_MPORT_4_data = pht_1_4[pht_1_4_MPORT_4_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_4_MPORT_12_en = pht_1_4_MPORT_12_en_pipe_0;
  assign pht_1_4_MPORT_12_addr = pht_1_4_MPORT_12_addr_pipe_0;
  assign pht_1_4_MPORT_12_data = pht_1_4[pht_1_4_MPORT_12_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_4_MPORT_24_en = pht_1_4_MPORT_24_en_pipe_0;
  assign pht_1_4_MPORT_24_addr = pht_1_4_MPORT_24_addr_pipe_0;
  assign pht_1_4_MPORT_24_data = pht_1_4[pht_1_4_MPORT_24_addr]; // @[PatternHistoryTable.scala 21:28]
  assign pht_1_4_MPORT_40_data = pht_wdata_w[1];
  assign pht_1_4_MPORT_40_addr = REG_43;
  assign pht_1_4_MPORT_40_mask = 1'h1;
  assign pht_1_4_MPORT_40_en = REG_29 & REG_42;
  assign pht_1_4_MPORT_560_data = 1'h0;
  assign pht_1_4_MPORT_560_addr = 6'h0;
  assign pht_1_4_MPORT_560_mask = 1'h1;
  assign pht_1_4_MPORT_560_en = reset;
  assign pht_1_4_MPORT_562_data = 1'h0;
  assign pht_1_4_MPORT_562_addr = 6'h1;
  assign pht_1_4_MPORT_562_mask = 1'h1;
  assign pht_1_4_MPORT_562_en = reset;
  assign pht_1_4_MPORT_564_data = 1'h0;
  assign pht_1_4_MPORT_564_addr = 6'h2;
  assign pht_1_4_MPORT_564_mask = 1'h1;
  assign pht_1_4_MPORT_564_en = reset;
  assign pht_1_4_MPORT_566_data = 1'h0;
  assign pht_1_4_MPORT_566_addr = 6'h3;
  assign pht_1_4_MPORT_566_mask = 1'h1;
  assign pht_1_4_MPORT_566_en = reset;
  assign pht_1_4_MPORT_568_data = 1'h0;
  assign pht_1_4_MPORT_568_addr = 6'h4;
  assign pht_1_4_MPORT_568_mask = 1'h1;
  assign pht_1_4_MPORT_568_en = reset;
  assign pht_1_4_MPORT_570_data = 1'h0;
  assign pht_1_4_MPORT_570_addr = 6'h5;
  assign pht_1_4_MPORT_570_mask = 1'h1;
  assign pht_1_4_MPORT_570_en = reset;
  assign pht_1_4_MPORT_572_data = 1'h0;
  assign pht_1_4_MPORT_572_addr = 6'h6;
  assign pht_1_4_MPORT_572_mask = 1'h1;
  assign pht_1_4_MPORT_572_en = reset;
  assign pht_1_4_MPORT_574_data = 1'h0;
  assign pht_1_4_MPORT_574_addr = 6'h7;
  assign pht_1_4_MPORT_574_mask = 1'h1;
  assign pht_1_4_MPORT_574_en = reset;
  assign pht_1_4_MPORT_576_data = 1'h0;
  assign pht_1_4_MPORT_576_addr = 6'h8;
  assign pht_1_4_MPORT_576_mask = 1'h1;
  assign pht_1_4_MPORT_576_en = reset;
  assign pht_1_4_MPORT_578_data = 1'h0;
  assign pht_1_4_MPORT_578_addr = 6'h9;
  assign pht_1_4_MPORT_578_mask = 1'h1;
  assign pht_1_4_MPORT_578_en = reset;
  assign pht_1_4_MPORT_580_data = 1'h0;
  assign pht_1_4_MPORT_580_addr = 6'ha;
  assign pht_1_4_MPORT_580_mask = 1'h1;
  assign pht_1_4_MPORT_580_en = reset;
  assign pht_1_4_MPORT_582_data = 1'h0;
  assign pht_1_4_MPORT_582_addr = 6'hb;
  assign pht_1_4_MPORT_582_mask = 1'h1;
  assign pht_1_4_MPORT_582_en = reset;
  assign pht_1_4_MPORT_584_data = 1'h0;
  assign pht_1_4_MPORT_584_addr = 6'hc;
  assign pht_1_4_MPORT_584_mask = 1'h1;
  assign pht_1_4_MPORT_584_en = reset;
  assign pht_1_4_MPORT_586_data = 1'h0;
  assign pht_1_4_MPORT_586_addr = 6'hd;
  assign pht_1_4_MPORT_586_mask = 1'h1;
  assign pht_1_4_MPORT_586_en = reset;
  assign pht_1_4_MPORT_588_data = 1'h0;
  assign pht_1_4_MPORT_588_addr = 6'he;
  assign pht_1_4_MPORT_588_mask = 1'h1;
  assign pht_1_4_MPORT_588_en = reset;
  assign pht_1_4_MPORT_590_data = 1'h0;
  assign pht_1_4_MPORT_590_addr = 6'hf;
  assign pht_1_4_MPORT_590_mask = 1'h1;
  assign pht_1_4_MPORT_590_en = reset;
  assign pht_1_4_MPORT_592_data = 1'h0;
  assign pht_1_4_MPORT_592_addr = 6'h10;
  assign pht_1_4_MPORT_592_mask = 1'h1;
  assign pht_1_4_MPORT_592_en = reset;
  assign pht_1_4_MPORT_594_data = 1'h0;
  assign pht_1_4_MPORT_594_addr = 6'h11;
  assign pht_1_4_MPORT_594_mask = 1'h1;
  assign pht_1_4_MPORT_594_en = reset;
  assign pht_1_4_MPORT_596_data = 1'h0;
  assign pht_1_4_MPORT_596_addr = 6'h12;
  assign pht_1_4_MPORT_596_mask = 1'h1;
  assign pht_1_4_MPORT_596_en = reset;
  assign pht_1_4_MPORT_598_data = 1'h0;
  assign pht_1_4_MPORT_598_addr = 6'h13;
  assign pht_1_4_MPORT_598_mask = 1'h1;
  assign pht_1_4_MPORT_598_en = reset;
  assign pht_1_4_MPORT_600_data = 1'h0;
  assign pht_1_4_MPORT_600_addr = 6'h14;
  assign pht_1_4_MPORT_600_mask = 1'h1;
  assign pht_1_4_MPORT_600_en = reset;
  assign pht_1_4_MPORT_602_data = 1'h0;
  assign pht_1_4_MPORT_602_addr = 6'h15;
  assign pht_1_4_MPORT_602_mask = 1'h1;
  assign pht_1_4_MPORT_602_en = reset;
  assign pht_1_4_MPORT_604_data = 1'h0;
  assign pht_1_4_MPORT_604_addr = 6'h16;
  assign pht_1_4_MPORT_604_mask = 1'h1;
  assign pht_1_4_MPORT_604_en = reset;
  assign pht_1_4_MPORT_606_data = 1'h0;
  assign pht_1_4_MPORT_606_addr = 6'h17;
  assign pht_1_4_MPORT_606_mask = 1'h1;
  assign pht_1_4_MPORT_606_en = reset;
  assign pht_1_4_MPORT_608_data = 1'h0;
  assign pht_1_4_MPORT_608_addr = 6'h18;
  assign pht_1_4_MPORT_608_mask = 1'h1;
  assign pht_1_4_MPORT_608_en = reset;
  assign pht_1_4_MPORT_610_data = 1'h0;
  assign pht_1_4_MPORT_610_addr = 6'h19;
  assign pht_1_4_MPORT_610_mask = 1'h1;
  assign pht_1_4_MPORT_610_en = reset;
  assign pht_1_4_MPORT_612_data = 1'h0;
  assign pht_1_4_MPORT_612_addr = 6'h1a;
  assign pht_1_4_MPORT_612_mask = 1'h1;
  assign pht_1_4_MPORT_612_en = reset;
  assign pht_1_4_MPORT_614_data = 1'h0;
  assign pht_1_4_MPORT_614_addr = 6'h1b;
  assign pht_1_4_MPORT_614_mask = 1'h1;
  assign pht_1_4_MPORT_614_en = reset;
  assign pht_1_4_MPORT_616_data = 1'h0;
  assign pht_1_4_MPORT_616_addr = 6'h1c;
  assign pht_1_4_MPORT_616_mask = 1'h1;
  assign pht_1_4_MPORT_616_en = reset;
  assign pht_1_4_MPORT_618_data = 1'h0;
  assign pht_1_4_MPORT_618_addr = 6'h1d;
  assign pht_1_4_MPORT_618_mask = 1'h1;
  assign pht_1_4_MPORT_618_en = reset;
  assign pht_1_4_MPORT_620_data = 1'h0;
  assign pht_1_4_MPORT_620_addr = 6'h1e;
  assign pht_1_4_MPORT_620_mask = 1'h1;
  assign pht_1_4_MPORT_620_en = reset;
  assign pht_1_4_MPORT_622_data = 1'h0;
  assign pht_1_4_MPORT_622_addr = 6'h1f;
  assign pht_1_4_MPORT_622_mask = 1'h1;
  assign pht_1_4_MPORT_622_en = reset;
  assign pht_1_4_MPORT_624_data = 1'h0;
  assign pht_1_4_MPORT_624_addr = 6'h20;
  assign pht_1_4_MPORT_624_mask = 1'h1;
  assign pht_1_4_MPORT_624_en = reset;
  assign pht_1_4_MPORT_626_data = 1'h0;
  assign pht_1_4_MPORT_626_addr = 6'h21;
  assign pht_1_4_MPORT_626_mask = 1'h1;
  assign pht_1_4_MPORT_626_en = reset;
  assign pht_1_4_MPORT_628_data = 1'h0;
  assign pht_1_4_MPORT_628_addr = 6'h22;
  assign pht_1_4_MPORT_628_mask = 1'h1;
  assign pht_1_4_MPORT_628_en = reset;
  assign pht_1_4_MPORT_630_data = 1'h0;
  assign pht_1_4_MPORT_630_addr = 6'h23;
  assign pht_1_4_MPORT_630_mask = 1'h1;
  assign pht_1_4_MPORT_630_en = reset;
  assign pht_1_4_MPORT_632_data = 1'h0;
  assign pht_1_4_MPORT_632_addr = 6'h24;
  assign pht_1_4_MPORT_632_mask = 1'h1;
  assign pht_1_4_MPORT_632_en = reset;
  assign pht_1_4_MPORT_634_data = 1'h0;
  assign pht_1_4_MPORT_634_addr = 6'h25;
  assign pht_1_4_MPORT_634_mask = 1'h1;
  assign pht_1_4_MPORT_634_en = reset;
  assign pht_1_4_MPORT_636_data = 1'h0;
  assign pht_1_4_MPORT_636_addr = 6'h26;
  assign pht_1_4_MPORT_636_mask = 1'h1;
  assign pht_1_4_MPORT_636_en = reset;
  assign pht_1_4_MPORT_638_data = 1'h0;
  assign pht_1_4_MPORT_638_addr = 6'h27;
  assign pht_1_4_MPORT_638_mask = 1'h1;
  assign pht_1_4_MPORT_638_en = reset;
  assign pht_1_4_MPORT_640_data = 1'h0;
  assign pht_1_4_MPORT_640_addr = 6'h28;
  assign pht_1_4_MPORT_640_mask = 1'h1;
  assign pht_1_4_MPORT_640_en = reset;
  assign pht_1_4_MPORT_642_data = 1'h0;
  assign pht_1_4_MPORT_642_addr = 6'h29;
  assign pht_1_4_MPORT_642_mask = 1'h1;
  assign pht_1_4_MPORT_642_en = reset;
  assign pht_1_4_MPORT_644_data = 1'h0;
  assign pht_1_4_MPORT_644_addr = 6'h2a;
  assign pht_1_4_MPORT_644_mask = 1'h1;
  assign pht_1_4_MPORT_644_en = reset;
  assign pht_1_4_MPORT_646_data = 1'h0;
  assign pht_1_4_MPORT_646_addr = 6'h2b;
  assign pht_1_4_MPORT_646_mask = 1'h1;
  assign pht_1_4_MPORT_646_en = reset;
  assign pht_1_4_MPORT_648_data = 1'h0;
  assign pht_1_4_MPORT_648_addr = 6'h2c;
  assign pht_1_4_MPORT_648_mask = 1'h1;
  assign pht_1_4_MPORT_648_en = reset;
  assign pht_1_4_MPORT_650_data = 1'h0;
  assign pht_1_4_MPORT_650_addr = 6'h2d;
  assign pht_1_4_MPORT_650_mask = 1'h1;
  assign pht_1_4_MPORT_650_en = reset;
  assign pht_1_4_MPORT_652_data = 1'h0;
  assign pht_1_4_MPORT_652_addr = 6'h2e;
  assign pht_1_4_MPORT_652_mask = 1'h1;
  assign pht_1_4_MPORT_652_en = reset;
  assign pht_1_4_MPORT_654_data = 1'h0;
  assign pht_1_4_MPORT_654_addr = 6'h2f;
  assign pht_1_4_MPORT_654_mask = 1'h1;
  assign pht_1_4_MPORT_654_en = reset;
  assign pht_1_4_MPORT_656_data = 1'h0;
  assign pht_1_4_MPORT_656_addr = 6'h30;
  assign pht_1_4_MPORT_656_mask = 1'h1;
  assign pht_1_4_MPORT_656_en = reset;
  assign pht_1_4_MPORT_658_data = 1'h0;
  assign pht_1_4_MPORT_658_addr = 6'h31;
  assign pht_1_4_MPORT_658_mask = 1'h1;
  assign pht_1_4_MPORT_658_en = reset;
  assign pht_1_4_MPORT_660_data = 1'h0;
  assign pht_1_4_MPORT_660_addr = 6'h32;
  assign pht_1_4_MPORT_660_mask = 1'h1;
  assign pht_1_4_MPORT_660_en = reset;
  assign pht_1_4_MPORT_662_data = 1'h0;
  assign pht_1_4_MPORT_662_addr = 6'h33;
  assign pht_1_4_MPORT_662_mask = 1'h1;
  assign pht_1_4_MPORT_662_en = reset;
  assign pht_1_4_MPORT_664_data = 1'h0;
  assign pht_1_4_MPORT_664_addr = 6'h34;
  assign pht_1_4_MPORT_664_mask = 1'h1;
  assign pht_1_4_MPORT_664_en = reset;
  assign pht_1_4_MPORT_666_data = 1'h0;
  assign pht_1_4_MPORT_666_addr = 6'h35;
  assign pht_1_4_MPORT_666_mask = 1'h1;
  assign pht_1_4_MPORT_666_en = reset;
  assign pht_1_4_MPORT_668_data = 1'h0;
  assign pht_1_4_MPORT_668_addr = 6'h36;
  assign pht_1_4_MPORT_668_mask = 1'h1;
  assign pht_1_4_MPORT_668_en = reset;
  assign pht_1_4_MPORT_670_data = 1'h0;
  assign pht_1_4_MPORT_670_addr = 6'h37;
  assign pht_1_4_MPORT_670_mask = 1'h1;
  assign pht_1_4_MPORT_670_en = reset;
  assign pht_1_4_MPORT_672_data = 1'h0;
  assign pht_1_4_MPORT_672_addr = 6'h38;
  assign pht_1_4_MPORT_672_mask = 1'h1;
  assign pht_1_4_MPORT_672_en = reset;
  assign pht_1_4_MPORT_674_data = 1'h0;
  assign pht_1_4_MPORT_674_addr = 6'h39;
  assign pht_1_4_MPORT_674_mask = 1'h1;
  assign pht_1_4_MPORT_674_en = reset;
  assign pht_1_4_MPORT_676_data = 1'h0;
  assign pht_1_4_MPORT_676_addr = 6'h3a;
  assign pht_1_4_MPORT_676_mask = 1'h1;
  assign pht_1_4_MPORT_676_en = reset;
  assign pht_1_4_MPORT_678_data = 1'h0;
  assign pht_1_4_MPORT_678_addr = 6'h3b;
  assign pht_1_4_MPORT_678_mask = 1'h1;
  assign pht_1_4_MPORT_678_en = reset;
  assign pht_1_4_MPORT_680_data = 1'h0;
  assign pht_1_4_MPORT_680_addr = 6'h3c;
  assign pht_1_4_MPORT_680_mask = 1'h1;
  assign pht_1_4_MPORT_680_en = reset;
  assign pht_1_4_MPORT_682_data = 1'h0;
  assign pht_1_4_MPORT_682_addr = 6'h3d;
  assign pht_1_4_MPORT_682_mask = 1'h1;
  assign pht_1_4_MPORT_682_en = reset;
  assign pht_1_4_MPORT_684_data = 1'h0;
  assign pht_1_4_MPORT_684_addr = 6'h3e;
  assign pht_1_4_MPORT_684_mask = 1'h1;
  assign pht_1_4_MPORT_684_en = reset;
  assign pht_1_4_MPORT_686_data = 1'h0;
  assign pht_1_4_MPORT_686_addr = 6'h3f;
  assign pht_1_4_MPORT_686_mask = 1'h1;
  assign pht_1_4_MPORT_686_en = reset;
//   assign pht_1_5_MPORT_5_en = pht_1_5_MPORT_5_en_pipe_0;
  assign pht_1_5_MPORT_5_addr = pht_1_5_MPORT_5_addr_pipe_0;
  assign pht_1_5_MPORT_5_data = pht_1_5[pht_1_5_MPORT_5_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_5_MPORT_13_en = pht_1_5_MPORT_13_en_pipe_0;
  assign pht_1_5_MPORT_13_addr = pht_1_5_MPORT_13_addr_pipe_0;
  assign pht_1_5_MPORT_13_data = pht_1_5[pht_1_5_MPORT_13_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_5_MPORT_26_en = pht_1_5_MPORT_26_en_pipe_0;
  assign pht_1_5_MPORT_26_addr = pht_1_5_MPORT_26_addr_pipe_0;
  assign pht_1_5_MPORT_26_data = pht_1_5[pht_1_5_MPORT_26_addr]; // @[PatternHistoryTable.scala 21:28]
  assign pht_1_5_MPORT_42_data = pht_wdata_w[1];
  assign pht_1_5_MPORT_42_addr = REG_46;
  assign pht_1_5_MPORT_42_mask = 1'h1;
  assign pht_1_5_MPORT_42_en = REG_29 & REG_45;
  assign pht_1_5_MPORT_688_data = 1'h0;
  assign pht_1_5_MPORT_688_addr = 6'h0;
  assign pht_1_5_MPORT_688_mask = 1'h1;
  assign pht_1_5_MPORT_688_en = reset;
  assign pht_1_5_MPORT_690_data = 1'h0;
  assign pht_1_5_MPORT_690_addr = 6'h1;
  assign pht_1_5_MPORT_690_mask = 1'h1;
  assign pht_1_5_MPORT_690_en = reset;
  assign pht_1_5_MPORT_692_data = 1'h0;
  assign pht_1_5_MPORT_692_addr = 6'h2;
  assign pht_1_5_MPORT_692_mask = 1'h1;
  assign pht_1_5_MPORT_692_en = reset;
  assign pht_1_5_MPORT_694_data = 1'h0;
  assign pht_1_5_MPORT_694_addr = 6'h3;
  assign pht_1_5_MPORT_694_mask = 1'h1;
  assign pht_1_5_MPORT_694_en = reset;
  assign pht_1_5_MPORT_696_data = 1'h0;
  assign pht_1_5_MPORT_696_addr = 6'h4;
  assign pht_1_5_MPORT_696_mask = 1'h1;
  assign pht_1_5_MPORT_696_en = reset;
  assign pht_1_5_MPORT_698_data = 1'h0;
  assign pht_1_5_MPORT_698_addr = 6'h5;
  assign pht_1_5_MPORT_698_mask = 1'h1;
  assign pht_1_5_MPORT_698_en = reset;
  assign pht_1_5_MPORT_700_data = 1'h0;
  assign pht_1_5_MPORT_700_addr = 6'h6;
  assign pht_1_5_MPORT_700_mask = 1'h1;
  assign pht_1_5_MPORT_700_en = reset;
  assign pht_1_5_MPORT_702_data = 1'h0;
  assign pht_1_5_MPORT_702_addr = 6'h7;
  assign pht_1_5_MPORT_702_mask = 1'h1;
  assign pht_1_5_MPORT_702_en = reset;
  assign pht_1_5_MPORT_704_data = 1'h0;
  assign pht_1_5_MPORT_704_addr = 6'h8;
  assign pht_1_5_MPORT_704_mask = 1'h1;
  assign pht_1_5_MPORT_704_en = reset;
  assign pht_1_5_MPORT_706_data = 1'h0;
  assign pht_1_5_MPORT_706_addr = 6'h9;
  assign pht_1_5_MPORT_706_mask = 1'h1;
  assign pht_1_5_MPORT_706_en = reset;
  assign pht_1_5_MPORT_708_data = 1'h0;
  assign pht_1_5_MPORT_708_addr = 6'ha;
  assign pht_1_5_MPORT_708_mask = 1'h1;
  assign pht_1_5_MPORT_708_en = reset;
  assign pht_1_5_MPORT_710_data = 1'h0;
  assign pht_1_5_MPORT_710_addr = 6'hb;
  assign pht_1_5_MPORT_710_mask = 1'h1;
  assign pht_1_5_MPORT_710_en = reset;
  assign pht_1_5_MPORT_712_data = 1'h0;
  assign pht_1_5_MPORT_712_addr = 6'hc;
  assign pht_1_5_MPORT_712_mask = 1'h1;
  assign pht_1_5_MPORT_712_en = reset;
  assign pht_1_5_MPORT_714_data = 1'h0;
  assign pht_1_5_MPORT_714_addr = 6'hd;
  assign pht_1_5_MPORT_714_mask = 1'h1;
  assign pht_1_5_MPORT_714_en = reset;
  assign pht_1_5_MPORT_716_data = 1'h0;
  assign pht_1_5_MPORT_716_addr = 6'he;
  assign pht_1_5_MPORT_716_mask = 1'h1;
  assign pht_1_5_MPORT_716_en = reset;
  assign pht_1_5_MPORT_718_data = 1'h0;
  assign pht_1_5_MPORT_718_addr = 6'hf;
  assign pht_1_5_MPORT_718_mask = 1'h1;
  assign pht_1_5_MPORT_718_en = reset;
  assign pht_1_5_MPORT_720_data = 1'h0;
  assign pht_1_5_MPORT_720_addr = 6'h10;
  assign pht_1_5_MPORT_720_mask = 1'h1;
  assign pht_1_5_MPORT_720_en = reset;
  assign pht_1_5_MPORT_722_data = 1'h0;
  assign pht_1_5_MPORT_722_addr = 6'h11;
  assign pht_1_5_MPORT_722_mask = 1'h1;
  assign pht_1_5_MPORT_722_en = reset;
  assign pht_1_5_MPORT_724_data = 1'h0;
  assign pht_1_5_MPORT_724_addr = 6'h12;
  assign pht_1_5_MPORT_724_mask = 1'h1;
  assign pht_1_5_MPORT_724_en = reset;
  assign pht_1_5_MPORT_726_data = 1'h0;
  assign pht_1_5_MPORT_726_addr = 6'h13;
  assign pht_1_5_MPORT_726_mask = 1'h1;
  assign pht_1_5_MPORT_726_en = reset;
  assign pht_1_5_MPORT_728_data = 1'h0;
  assign pht_1_5_MPORT_728_addr = 6'h14;
  assign pht_1_5_MPORT_728_mask = 1'h1;
  assign pht_1_5_MPORT_728_en = reset;
  assign pht_1_5_MPORT_730_data = 1'h0;
  assign pht_1_5_MPORT_730_addr = 6'h15;
  assign pht_1_5_MPORT_730_mask = 1'h1;
  assign pht_1_5_MPORT_730_en = reset;
  assign pht_1_5_MPORT_732_data = 1'h0;
  assign pht_1_5_MPORT_732_addr = 6'h16;
  assign pht_1_5_MPORT_732_mask = 1'h1;
  assign pht_1_5_MPORT_732_en = reset;
  assign pht_1_5_MPORT_734_data = 1'h0;
  assign pht_1_5_MPORT_734_addr = 6'h17;
  assign pht_1_5_MPORT_734_mask = 1'h1;
  assign pht_1_5_MPORT_734_en = reset;
  assign pht_1_5_MPORT_736_data = 1'h0;
  assign pht_1_5_MPORT_736_addr = 6'h18;
  assign pht_1_5_MPORT_736_mask = 1'h1;
  assign pht_1_5_MPORT_736_en = reset;
  assign pht_1_5_MPORT_738_data = 1'h0;
  assign pht_1_5_MPORT_738_addr = 6'h19;
  assign pht_1_5_MPORT_738_mask = 1'h1;
  assign pht_1_5_MPORT_738_en = reset;
  assign pht_1_5_MPORT_740_data = 1'h0;
  assign pht_1_5_MPORT_740_addr = 6'h1a;
  assign pht_1_5_MPORT_740_mask = 1'h1;
  assign pht_1_5_MPORT_740_en = reset;
  assign pht_1_5_MPORT_742_data = 1'h0;
  assign pht_1_5_MPORT_742_addr = 6'h1b;
  assign pht_1_5_MPORT_742_mask = 1'h1;
  assign pht_1_5_MPORT_742_en = reset;
  assign pht_1_5_MPORT_744_data = 1'h0;
  assign pht_1_5_MPORT_744_addr = 6'h1c;
  assign pht_1_5_MPORT_744_mask = 1'h1;
  assign pht_1_5_MPORT_744_en = reset;
  assign pht_1_5_MPORT_746_data = 1'h0;
  assign pht_1_5_MPORT_746_addr = 6'h1d;
  assign pht_1_5_MPORT_746_mask = 1'h1;
  assign pht_1_5_MPORT_746_en = reset;
  assign pht_1_5_MPORT_748_data = 1'h0;
  assign pht_1_5_MPORT_748_addr = 6'h1e;
  assign pht_1_5_MPORT_748_mask = 1'h1;
  assign pht_1_5_MPORT_748_en = reset;
  assign pht_1_5_MPORT_750_data = 1'h0;
  assign pht_1_5_MPORT_750_addr = 6'h1f;
  assign pht_1_5_MPORT_750_mask = 1'h1;
  assign pht_1_5_MPORT_750_en = reset;
  assign pht_1_5_MPORT_752_data = 1'h0;
  assign pht_1_5_MPORT_752_addr = 6'h20;
  assign pht_1_5_MPORT_752_mask = 1'h1;
  assign pht_1_5_MPORT_752_en = reset;
  assign pht_1_5_MPORT_754_data = 1'h0;
  assign pht_1_5_MPORT_754_addr = 6'h21;
  assign pht_1_5_MPORT_754_mask = 1'h1;
  assign pht_1_5_MPORT_754_en = reset;
  assign pht_1_5_MPORT_756_data = 1'h0;
  assign pht_1_5_MPORT_756_addr = 6'h22;
  assign pht_1_5_MPORT_756_mask = 1'h1;
  assign pht_1_5_MPORT_756_en = reset;
  assign pht_1_5_MPORT_758_data = 1'h0;
  assign pht_1_5_MPORT_758_addr = 6'h23;
  assign pht_1_5_MPORT_758_mask = 1'h1;
  assign pht_1_5_MPORT_758_en = reset;
  assign pht_1_5_MPORT_760_data = 1'h0;
  assign pht_1_5_MPORT_760_addr = 6'h24;
  assign pht_1_5_MPORT_760_mask = 1'h1;
  assign pht_1_5_MPORT_760_en = reset;
  assign pht_1_5_MPORT_762_data = 1'h0;
  assign pht_1_5_MPORT_762_addr = 6'h25;
  assign pht_1_5_MPORT_762_mask = 1'h1;
  assign pht_1_5_MPORT_762_en = reset;
  assign pht_1_5_MPORT_764_data = 1'h0;
  assign pht_1_5_MPORT_764_addr = 6'h26;
  assign pht_1_5_MPORT_764_mask = 1'h1;
  assign pht_1_5_MPORT_764_en = reset;
  assign pht_1_5_MPORT_766_data = 1'h0;
  assign pht_1_5_MPORT_766_addr = 6'h27;
  assign pht_1_5_MPORT_766_mask = 1'h1;
  assign pht_1_5_MPORT_766_en = reset;
  assign pht_1_5_MPORT_768_data = 1'h0;
  assign pht_1_5_MPORT_768_addr = 6'h28;
  assign pht_1_5_MPORT_768_mask = 1'h1;
  assign pht_1_5_MPORT_768_en = reset;
  assign pht_1_5_MPORT_770_data = 1'h0;
  assign pht_1_5_MPORT_770_addr = 6'h29;
  assign pht_1_5_MPORT_770_mask = 1'h1;
  assign pht_1_5_MPORT_770_en = reset;
  assign pht_1_5_MPORT_772_data = 1'h0;
  assign pht_1_5_MPORT_772_addr = 6'h2a;
  assign pht_1_5_MPORT_772_mask = 1'h1;
  assign pht_1_5_MPORT_772_en = reset;
  assign pht_1_5_MPORT_774_data = 1'h0;
  assign pht_1_5_MPORT_774_addr = 6'h2b;
  assign pht_1_5_MPORT_774_mask = 1'h1;
  assign pht_1_5_MPORT_774_en = reset;
  assign pht_1_5_MPORT_776_data = 1'h0;
  assign pht_1_5_MPORT_776_addr = 6'h2c;
  assign pht_1_5_MPORT_776_mask = 1'h1;
  assign pht_1_5_MPORT_776_en = reset;
  assign pht_1_5_MPORT_778_data = 1'h0;
  assign pht_1_5_MPORT_778_addr = 6'h2d;
  assign pht_1_5_MPORT_778_mask = 1'h1;
  assign pht_1_5_MPORT_778_en = reset;
  assign pht_1_5_MPORT_780_data = 1'h0;
  assign pht_1_5_MPORT_780_addr = 6'h2e;
  assign pht_1_5_MPORT_780_mask = 1'h1;
  assign pht_1_5_MPORT_780_en = reset;
  assign pht_1_5_MPORT_782_data = 1'h0;
  assign pht_1_5_MPORT_782_addr = 6'h2f;
  assign pht_1_5_MPORT_782_mask = 1'h1;
  assign pht_1_5_MPORT_782_en = reset;
  assign pht_1_5_MPORT_784_data = 1'h0;
  assign pht_1_5_MPORT_784_addr = 6'h30;
  assign pht_1_5_MPORT_784_mask = 1'h1;
  assign pht_1_5_MPORT_784_en = reset;
  assign pht_1_5_MPORT_786_data = 1'h0;
  assign pht_1_5_MPORT_786_addr = 6'h31;
  assign pht_1_5_MPORT_786_mask = 1'h1;
  assign pht_1_5_MPORT_786_en = reset;
  assign pht_1_5_MPORT_788_data = 1'h0;
  assign pht_1_5_MPORT_788_addr = 6'h32;
  assign pht_1_5_MPORT_788_mask = 1'h1;
  assign pht_1_5_MPORT_788_en = reset;
  assign pht_1_5_MPORT_790_data = 1'h0;
  assign pht_1_5_MPORT_790_addr = 6'h33;
  assign pht_1_5_MPORT_790_mask = 1'h1;
  assign pht_1_5_MPORT_790_en = reset;
  assign pht_1_5_MPORT_792_data = 1'h0;
  assign pht_1_5_MPORT_792_addr = 6'h34;
  assign pht_1_5_MPORT_792_mask = 1'h1;
  assign pht_1_5_MPORT_792_en = reset;
  assign pht_1_5_MPORT_794_data = 1'h0;
  assign pht_1_5_MPORT_794_addr = 6'h35;
  assign pht_1_5_MPORT_794_mask = 1'h1;
  assign pht_1_5_MPORT_794_en = reset;
  assign pht_1_5_MPORT_796_data = 1'h0;
  assign pht_1_5_MPORT_796_addr = 6'h36;
  assign pht_1_5_MPORT_796_mask = 1'h1;
  assign pht_1_5_MPORT_796_en = reset;
  assign pht_1_5_MPORT_798_data = 1'h0;
  assign pht_1_5_MPORT_798_addr = 6'h37;
  assign pht_1_5_MPORT_798_mask = 1'h1;
  assign pht_1_5_MPORT_798_en = reset;
  assign pht_1_5_MPORT_800_data = 1'h0;
  assign pht_1_5_MPORT_800_addr = 6'h38;
  assign pht_1_5_MPORT_800_mask = 1'h1;
  assign pht_1_5_MPORT_800_en = reset;
  assign pht_1_5_MPORT_802_data = 1'h0;
  assign pht_1_5_MPORT_802_addr = 6'h39;
  assign pht_1_5_MPORT_802_mask = 1'h1;
  assign pht_1_5_MPORT_802_en = reset;
  assign pht_1_5_MPORT_804_data = 1'h0;
  assign pht_1_5_MPORT_804_addr = 6'h3a;
  assign pht_1_5_MPORT_804_mask = 1'h1;
  assign pht_1_5_MPORT_804_en = reset;
  assign pht_1_5_MPORT_806_data = 1'h0;
  assign pht_1_5_MPORT_806_addr = 6'h3b;
  assign pht_1_5_MPORT_806_mask = 1'h1;
  assign pht_1_5_MPORT_806_en = reset;
  assign pht_1_5_MPORT_808_data = 1'h0;
  assign pht_1_5_MPORT_808_addr = 6'h3c;
  assign pht_1_5_MPORT_808_mask = 1'h1;
  assign pht_1_5_MPORT_808_en = reset;
  assign pht_1_5_MPORT_810_data = 1'h0;
  assign pht_1_5_MPORT_810_addr = 6'h3d;
  assign pht_1_5_MPORT_810_mask = 1'h1;
  assign pht_1_5_MPORT_810_en = reset;
  assign pht_1_5_MPORT_812_data = 1'h0;
  assign pht_1_5_MPORT_812_addr = 6'h3e;
  assign pht_1_5_MPORT_812_mask = 1'h1;
  assign pht_1_5_MPORT_812_en = reset;
  assign pht_1_5_MPORT_814_data = 1'h0;
  assign pht_1_5_MPORT_814_addr = 6'h3f;
  assign pht_1_5_MPORT_814_mask = 1'h1;
  assign pht_1_5_MPORT_814_en = reset;
//   assign pht_1_6_MPORT_6_en = pht_1_6_MPORT_6_en_pipe_0;
  assign pht_1_6_MPORT_6_addr = pht_1_6_MPORT_6_addr_pipe_0;
  assign pht_1_6_MPORT_6_data = pht_1_6[pht_1_6_MPORT_6_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_6_MPORT_14_en = pht_1_6_MPORT_14_en_pipe_0;
  assign pht_1_6_MPORT_14_addr = pht_1_6_MPORT_14_addr_pipe_0;
  assign pht_1_6_MPORT_14_data = pht_1_6[pht_1_6_MPORT_14_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_6_MPORT_28_en = pht_1_6_MPORT_28_en_pipe_0;
  assign pht_1_6_MPORT_28_addr = pht_1_6_MPORT_28_addr_pipe_0;
  assign pht_1_6_MPORT_28_data = pht_1_6[pht_1_6_MPORT_28_addr]; // @[PatternHistoryTable.scala 21:28]
  assign pht_1_6_MPORT_44_data = pht_wdata_w[1];
  assign pht_1_6_MPORT_44_addr = REG_49;
  assign pht_1_6_MPORT_44_mask = 1'h1;
  assign pht_1_6_MPORT_44_en = REG_29 & REG_48;
  assign pht_1_6_MPORT_816_data = 1'h0;
  assign pht_1_6_MPORT_816_addr = 6'h0;
  assign pht_1_6_MPORT_816_mask = 1'h1;
  assign pht_1_6_MPORT_816_en = reset;
  assign pht_1_6_MPORT_818_data = 1'h0;
  assign pht_1_6_MPORT_818_addr = 6'h1;
  assign pht_1_6_MPORT_818_mask = 1'h1;
  assign pht_1_6_MPORT_818_en = reset;
  assign pht_1_6_MPORT_820_data = 1'h0;
  assign pht_1_6_MPORT_820_addr = 6'h2;
  assign pht_1_6_MPORT_820_mask = 1'h1;
  assign pht_1_6_MPORT_820_en = reset;
  assign pht_1_6_MPORT_822_data = 1'h0;
  assign pht_1_6_MPORT_822_addr = 6'h3;
  assign pht_1_6_MPORT_822_mask = 1'h1;
  assign pht_1_6_MPORT_822_en = reset;
  assign pht_1_6_MPORT_824_data = 1'h0;
  assign pht_1_6_MPORT_824_addr = 6'h4;
  assign pht_1_6_MPORT_824_mask = 1'h1;
  assign pht_1_6_MPORT_824_en = reset;
  assign pht_1_6_MPORT_826_data = 1'h0;
  assign pht_1_6_MPORT_826_addr = 6'h5;
  assign pht_1_6_MPORT_826_mask = 1'h1;
  assign pht_1_6_MPORT_826_en = reset;
  assign pht_1_6_MPORT_828_data = 1'h0;
  assign pht_1_6_MPORT_828_addr = 6'h6;
  assign pht_1_6_MPORT_828_mask = 1'h1;
  assign pht_1_6_MPORT_828_en = reset;
  assign pht_1_6_MPORT_830_data = 1'h0;
  assign pht_1_6_MPORT_830_addr = 6'h7;
  assign pht_1_6_MPORT_830_mask = 1'h1;
  assign pht_1_6_MPORT_830_en = reset;
  assign pht_1_6_MPORT_832_data = 1'h0;
  assign pht_1_6_MPORT_832_addr = 6'h8;
  assign pht_1_6_MPORT_832_mask = 1'h1;
  assign pht_1_6_MPORT_832_en = reset;
  assign pht_1_6_MPORT_834_data = 1'h0;
  assign pht_1_6_MPORT_834_addr = 6'h9;
  assign pht_1_6_MPORT_834_mask = 1'h1;
  assign pht_1_6_MPORT_834_en = reset;
  assign pht_1_6_MPORT_836_data = 1'h0;
  assign pht_1_6_MPORT_836_addr = 6'ha;
  assign pht_1_6_MPORT_836_mask = 1'h1;
  assign pht_1_6_MPORT_836_en = reset;
  assign pht_1_6_MPORT_838_data = 1'h0;
  assign pht_1_6_MPORT_838_addr = 6'hb;
  assign pht_1_6_MPORT_838_mask = 1'h1;
  assign pht_1_6_MPORT_838_en = reset;
  assign pht_1_6_MPORT_840_data = 1'h0;
  assign pht_1_6_MPORT_840_addr = 6'hc;
  assign pht_1_6_MPORT_840_mask = 1'h1;
  assign pht_1_6_MPORT_840_en = reset;
  assign pht_1_6_MPORT_842_data = 1'h0;
  assign pht_1_6_MPORT_842_addr = 6'hd;
  assign pht_1_6_MPORT_842_mask = 1'h1;
  assign pht_1_6_MPORT_842_en = reset;
  assign pht_1_6_MPORT_844_data = 1'h0;
  assign pht_1_6_MPORT_844_addr = 6'he;
  assign pht_1_6_MPORT_844_mask = 1'h1;
  assign pht_1_6_MPORT_844_en = reset;
  assign pht_1_6_MPORT_846_data = 1'h0;
  assign pht_1_6_MPORT_846_addr = 6'hf;
  assign pht_1_6_MPORT_846_mask = 1'h1;
  assign pht_1_6_MPORT_846_en = reset;
  assign pht_1_6_MPORT_848_data = 1'h0;
  assign pht_1_6_MPORT_848_addr = 6'h10;
  assign pht_1_6_MPORT_848_mask = 1'h1;
  assign pht_1_6_MPORT_848_en = reset;
  assign pht_1_6_MPORT_850_data = 1'h0;
  assign pht_1_6_MPORT_850_addr = 6'h11;
  assign pht_1_6_MPORT_850_mask = 1'h1;
  assign pht_1_6_MPORT_850_en = reset;
  assign pht_1_6_MPORT_852_data = 1'h0;
  assign pht_1_6_MPORT_852_addr = 6'h12;
  assign pht_1_6_MPORT_852_mask = 1'h1;
  assign pht_1_6_MPORT_852_en = reset;
  assign pht_1_6_MPORT_854_data = 1'h0;
  assign pht_1_6_MPORT_854_addr = 6'h13;
  assign pht_1_6_MPORT_854_mask = 1'h1;
  assign pht_1_6_MPORT_854_en = reset;
  assign pht_1_6_MPORT_856_data = 1'h0;
  assign pht_1_6_MPORT_856_addr = 6'h14;
  assign pht_1_6_MPORT_856_mask = 1'h1;
  assign pht_1_6_MPORT_856_en = reset;
  assign pht_1_6_MPORT_858_data = 1'h0;
  assign pht_1_6_MPORT_858_addr = 6'h15;
  assign pht_1_6_MPORT_858_mask = 1'h1;
  assign pht_1_6_MPORT_858_en = reset;
  assign pht_1_6_MPORT_860_data = 1'h0;
  assign pht_1_6_MPORT_860_addr = 6'h16;
  assign pht_1_6_MPORT_860_mask = 1'h1;
  assign pht_1_6_MPORT_860_en = reset;
  assign pht_1_6_MPORT_862_data = 1'h0;
  assign pht_1_6_MPORT_862_addr = 6'h17;
  assign pht_1_6_MPORT_862_mask = 1'h1;
  assign pht_1_6_MPORT_862_en = reset;
  assign pht_1_6_MPORT_864_data = 1'h0;
  assign pht_1_6_MPORT_864_addr = 6'h18;
  assign pht_1_6_MPORT_864_mask = 1'h1;
  assign pht_1_6_MPORT_864_en = reset;
  assign pht_1_6_MPORT_866_data = 1'h0;
  assign pht_1_6_MPORT_866_addr = 6'h19;
  assign pht_1_6_MPORT_866_mask = 1'h1;
  assign pht_1_6_MPORT_866_en = reset;
  assign pht_1_6_MPORT_868_data = 1'h0;
  assign pht_1_6_MPORT_868_addr = 6'h1a;
  assign pht_1_6_MPORT_868_mask = 1'h1;
  assign pht_1_6_MPORT_868_en = reset;
  assign pht_1_6_MPORT_870_data = 1'h0;
  assign pht_1_6_MPORT_870_addr = 6'h1b;
  assign pht_1_6_MPORT_870_mask = 1'h1;
  assign pht_1_6_MPORT_870_en = reset;
  assign pht_1_6_MPORT_872_data = 1'h0;
  assign pht_1_6_MPORT_872_addr = 6'h1c;
  assign pht_1_6_MPORT_872_mask = 1'h1;
  assign pht_1_6_MPORT_872_en = reset;
  assign pht_1_6_MPORT_874_data = 1'h0;
  assign pht_1_6_MPORT_874_addr = 6'h1d;
  assign pht_1_6_MPORT_874_mask = 1'h1;
  assign pht_1_6_MPORT_874_en = reset;
  assign pht_1_6_MPORT_876_data = 1'h0;
  assign pht_1_6_MPORT_876_addr = 6'h1e;
  assign pht_1_6_MPORT_876_mask = 1'h1;
  assign pht_1_6_MPORT_876_en = reset;
  assign pht_1_6_MPORT_878_data = 1'h0;
  assign pht_1_6_MPORT_878_addr = 6'h1f;
  assign pht_1_6_MPORT_878_mask = 1'h1;
  assign pht_1_6_MPORT_878_en = reset;
  assign pht_1_6_MPORT_880_data = 1'h0;
  assign pht_1_6_MPORT_880_addr = 6'h20;
  assign pht_1_6_MPORT_880_mask = 1'h1;
  assign pht_1_6_MPORT_880_en = reset;
  assign pht_1_6_MPORT_882_data = 1'h0;
  assign pht_1_6_MPORT_882_addr = 6'h21;
  assign pht_1_6_MPORT_882_mask = 1'h1;
  assign pht_1_6_MPORT_882_en = reset;
  assign pht_1_6_MPORT_884_data = 1'h0;
  assign pht_1_6_MPORT_884_addr = 6'h22;
  assign pht_1_6_MPORT_884_mask = 1'h1;
  assign pht_1_6_MPORT_884_en = reset;
  assign pht_1_6_MPORT_886_data = 1'h0;
  assign pht_1_6_MPORT_886_addr = 6'h23;
  assign pht_1_6_MPORT_886_mask = 1'h1;
  assign pht_1_6_MPORT_886_en = reset;
  assign pht_1_6_MPORT_888_data = 1'h0;
  assign pht_1_6_MPORT_888_addr = 6'h24;
  assign pht_1_6_MPORT_888_mask = 1'h1;
  assign pht_1_6_MPORT_888_en = reset;
  assign pht_1_6_MPORT_890_data = 1'h0;
  assign pht_1_6_MPORT_890_addr = 6'h25;
  assign pht_1_6_MPORT_890_mask = 1'h1;
  assign pht_1_6_MPORT_890_en = reset;
  assign pht_1_6_MPORT_892_data = 1'h0;
  assign pht_1_6_MPORT_892_addr = 6'h26;
  assign pht_1_6_MPORT_892_mask = 1'h1;
  assign pht_1_6_MPORT_892_en = reset;
  assign pht_1_6_MPORT_894_data = 1'h0;
  assign pht_1_6_MPORT_894_addr = 6'h27;
  assign pht_1_6_MPORT_894_mask = 1'h1;
  assign pht_1_6_MPORT_894_en = reset;
  assign pht_1_6_MPORT_896_data = 1'h0;
  assign pht_1_6_MPORT_896_addr = 6'h28;
  assign pht_1_6_MPORT_896_mask = 1'h1;
  assign pht_1_6_MPORT_896_en = reset;
  assign pht_1_6_MPORT_898_data = 1'h0;
  assign pht_1_6_MPORT_898_addr = 6'h29;
  assign pht_1_6_MPORT_898_mask = 1'h1;
  assign pht_1_6_MPORT_898_en = reset;
  assign pht_1_6_MPORT_900_data = 1'h0;
  assign pht_1_6_MPORT_900_addr = 6'h2a;
  assign pht_1_6_MPORT_900_mask = 1'h1;
  assign pht_1_6_MPORT_900_en = reset;
  assign pht_1_6_MPORT_902_data = 1'h0;
  assign pht_1_6_MPORT_902_addr = 6'h2b;
  assign pht_1_6_MPORT_902_mask = 1'h1;
  assign pht_1_6_MPORT_902_en = reset;
  assign pht_1_6_MPORT_904_data = 1'h0;
  assign pht_1_6_MPORT_904_addr = 6'h2c;
  assign pht_1_6_MPORT_904_mask = 1'h1;
  assign pht_1_6_MPORT_904_en = reset;
  assign pht_1_6_MPORT_906_data = 1'h0;
  assign pht_1_6_MPORT_906_addr = 6'h2d;
  assign pht_1_6_MPORT_906_mask = 1'h1;
  assign pht_1_6_MPORT_906_en = reset;
  assign pht_1_6_MPORT_908_data = 1'h0;
  assign pht_1_6_MPORT_908_addr = 6'h2e;
  assign pht_1_6_MPORT_908_mask = 1'h1;
  assign pht_1_6_MPORT_908_en = reset;
  assign pht_1_6_MPORT_910_data = 1'h0;
  assign pht_1_6_MPORT_910_addr = 6'h2f;
  assign pht_1_6_MPORT_910_mask = 1'h1;
  assign pht_1_6_MPORT_910_en = reset;
  assign pht_1_6_MPORT_912_data = 1'h0;
  assign pht_1_6_MPORT_912_addr = 6'h30;
  assign pht_1_6_MPORT_912_mask = 1'h1;
  assign pht_1_6_MPORT_912_en = reset;
  assign pht_1_6_MPORT_914_data = 1'h0;
  assign pht_1_6_MPORT_914_addr = 6'h31;
  assign pht_1_6_MPORT_914_mask = 1'h1;
  assign pht_1_6_MPORT_914_en = reset;
  assign pht_1_6_MPORT_916_data = 1'h0;
  assign pht_1_6_MPORT_916_addr = 6'h32;
  assign pht_1_6_MPORT_916_mask = 1'h1;
  assign pht_1_6_MPORT_916_en = reset;
  assign pht_1_6_MPORT_918_data = 1'h0;
  assign pht_1_6_MPORT_918_addr = 6'h33;
  assign pht_1_6_MPORT_918_mask = 1'h1;
  assign pht_1_6_MPORT_918_en = reset;
  assign pht_1_6_MPORT_920_data = 1'h0;
  assign pht_1_6_MPORT_920_addr = 6'h34;
  assign pht_1_6_MPORT_920_mask = 1'h1;
  assign pht_1_6_MPORT_920_en = reset;
  assign pht_1_6_MPORT_922_data = 1'h0;
  assign pht_1_6_MPORT_922_addr = 6'h35;
  assign pht_1_6_MPORT_922_mask = 1'h1;
  assign pht_1_6_MPORT_922_en = reset;
  assign pht_1_6_MPORT_924_data = 1'h0;
  assign pht_1_6_MPORT_924_addr = 6'h36;
  assign pht_1_6_MPORT_924_mask = 1'h1;
  assign pht_1_6_MPORT_924_en = reset;
  assign pht_1_6_MPORT_926_data = 1'h0;
  assign pht_1_6_MPORT_926_addr = 6'h37;
  assign pht_1_6_MPORT_926_mask = 1'h1;
  assign pht_1_6_MPORT_926_en = reset;
  assign pht_1_6_MPORT_928_data = 1'h0;
  assign pht_1_6_MPORT_928_addr = 6'h38;
  assign pht_1_6_MPORT_928_mask = 1'h1;
  assign pht_1_6_MPORT_928_en = reset;
  assign pht_1_6_MPORT_930_data = 1'h0;
  assign pht_1_6_MPORT_930_addr = 6'h39;
  assign pht_1_6_MPORT_930_mask = 1'h1;
  assign pht_1_6_MPORT_930_en = reset;
  assign pht_1_6_MPORT_932_data = 1'h0;
  assign pht_1_6_MPORT_932_addr = 6'h3a;
  assign pht_1_6_MPORT_932_mask = 1'h1;
  assign pht_1_6_MPORT_932_en = reset;
  assign pht_1_6_MPORT_934_data = 1'h0;
  assign pht_1_6_MPORT_934_addr = 6'h3b;
  assign pht_1_6_MPORT_934_mask = 1'h1;
  assign pht_1_6_MPORT_934_en = reset;
  assign pht_1_6_MPORT_936_data = 1'h0;
  assign pht_1_6_MPORT_936_addr = 6'h3c;
  assign pht_1_6_MPORT_936_mask = 1'h1;
  assign pht_1_6_MPORT_936_en = reset;
  assign pht_1_6_MPORT_938_data = 1'h0;
  assign pht_1_6_MPORT_938_addr = 6'h3d;
  assign pht_1_6_MPORT_938_mask = 1'h1;
  assign pht_1_6_MPORT_938_en = reset;
  assign pht_1_6_MPORT_940_data = 1'h0;
  assign pht_1_6_MPORT_940_addr = 6'h3e;
  assign pht_1_6_MPORT_940_mask = 1'h1;
  assign pht_1_6_MPORT_940_en = reset;
  assign pht_1_6_MPORT_942_data = 1'h0;
  assign pht_1_6_MPORT_942_addr = 6'h3f;
  assign pht_1_6_MPORT_942_mask = 1'h1;
  assign pht_1_6_MPORT_942_en = reset;
//   assign pht_1_7_MPORT_7_en = pht_1_7_MPORT_7_en_pipe_0;
  assign pht_1_7_MPORT_7_addr = pht_1_7_MPORT_7_addr_pipe_0;
  assign pht_1_7_MPORT_7_data = pht_1_7[pht_1_7_MPORT_7_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_7_MPORT_15_en = pht_1_7_MPORT_15_en_pipe_0;
  assign pht_1_7_MPORT_15_addr = pht_1_7_MPORT_15_addr_pipe_0;
  assign pht_1_7_MPORT_15_data = pht_1_7[pht_1_7_MPORT_15_addr]; // @[PatternHistoryTable.scala 21:28]
//   assign pht_1_7_MPORT_30_en = pht_1_7_MPORT_30_en_pipe_0;
  assign pht_1_7_MPORT_30_addr = pht_1_7_MPORT_30_addr_pipe_0;
  assign pht_1_7_MPORT_30_data = pht_1_7[pht_1_7_MPORT_30_addr]; // @[PatternHistoryTable.scala 21:28]
  assign pht_1_7_MPORT_46_data = pht_wdata_w[1];
  assign pht_1_7_MPORT_46_addr = REG_52;
  assign pht_1_7_MPORT_46_mask = 1'h1;
  assign pht_1_7_MPORT_46_en = REG_29 & REG_51;
  assign pht_1_7_MPORT_944_data = 1'h0;
  assign pht_1_7_MPORT_944_addr = 6'h0;
  assign pht_1_7_MPORT_944_mask = 1'h1;
  assign pht_1_7_MPORT_944_en = reset;
  assign pht_1_7_MPORT_946_data = 1'h0;
  assign pht_1_7_MPORT_946_addr = 6'h1;
  assign pht_1_7_MPORT_946_mask = 1'h1;
  assign pht_1_7_MPORT_946_en = reset;
  assign pht_1_7_MPORT_948_data = 1'h0;
  assign pht_1_7_MPORT_948_addr = 6'h2;
  assign pht_1_7_MPORT_948_mask = 1'h1;
  assign pht_1_7_MPORT_948_en = reset;
  assign pht_1_7_MPORT_950_data = 1'h0;
  assign pht_1_7_MPORT_950_addr = 6'h3;
  assign pht_1_7_MPORT_950_mask = 1'h1;
  assign pht_1_7_MPORT_950_en = reset;
  assign pht_1_7_MPORT_952_data = 1'h0;
  assign pht_1_7_MPORT_952_addr = 6'h4;
  assign pht_1_7_MPORT_952_mask = 1'h1;
  assign pht_1_7_MPORT_952_en = reset;
  assign pht_1_7_MPORT_954_data = 1'h0;
  assign pht_1_7_MPORT_954_addr = 6'h5;
  assign pht_1_7_MPORT_954_mask = 1'h1;
  assign pht_1_7_MPORT_954_en = reset;
  assign pht_1_7_MPORT_956_data = 1'h0;
  assign pht_1_7_MPORT_956_addr = 6'h6;
  assign pht_1_7_MPORT_956_mask = 1'h1;
  assign pht_1_7_MPORT_956_en = reset;
  assign pht_1_7_MPORT_958_data = 1'h0;
  assign pht_1_7_MPORT_958_addr = 6'h7;
  assign pht_1_7_MPORT_958_mask = 1'h1;
  assign pht_1_7_MPORT_958_en = reset;
  assign pht_1_7_MPORT_960_data = 1'h0;
  assign pht_1_7_MPORT_960_addr = 6'h8;
  assign pht_1_7_MPORT_960_mask = 1'h1;
  assign pht_1_7_MPORT_960_en = reset;
  assign pht_1_7_MPORT_962_data = 1'h0;
  assign pht_1_7_MPORT_962_addr = 6'h9;
  assign pht_1_7_MPORT_962_mask = 1'h1;
  assign pht_1_7_MPORT_962_en = reset;
  assign pht_1_7_MPORT_964_data = 1'h0;
  assign pht_1_7_MPORT_964_addr = 6'ha;
  assign pht_1_7_MPORT_964_mask = 1'h1;
  assign pht_1_7_MPORT_964_en = reset;
  assign pht_1_7_MPORT_966_data = 1'h0;
  assign pht_1_7_MPORT_966_addr = 6'hb;
  assign pht_1_7_MPORT_966_mask = 1'h1;
  assign pht_1_7_MPORT_966_en = reset;
  assign pht_1_7_MPORT_968_data = 1'h0;
  assign pht_1_7_MPORT_968_addr = 6'hc;
  assign pht_1_7_MPORT_968_mask = 1'h1;
  assign pht_1_7_MPORT_968_en = reset;
  assign pht_1_7_MPORT_970_data = 1'h0;
  assign pht_1_7_MPORT_970_addr = 6'hd;
  assign pht_1_7_MPORT_970_mask = 1'h1;
  assign pht_1_7_MPORT_970_en = reset;
  assign pht_1_7_MPORT_972_data = 1'h0;
  assign pht_1_7_MPORT_972_addr = 6'he;
  assign pht_1_7_MPORT_972_mask = 1'h1;
  assign pht_1_7_MPORT_972_en = reset;
  assign pht_1_7_MPORT_974_data = 1'h0;
  assign pht_1_7_MPORT_974_addr = 6'hf;
  assign pht_1_7_MPORT_974_mask = 1'h1;
  assign pht_1_7_MPORT_974_en = reset;
  assign pht_1_7_MPORT_976_data = 1'h0;
  assign pht_1_7_MPORT_976_addr = 6'h10;
  assign pht_1_7_MPORT_976_mask = 1'h1;
  assign pht_1_7_MPORT_976_en = reset;
  assign pht_1_7_MPORT_978_data = 1'h0;
  assign pht_1_7_MPORT_978_addr = 6'h11;
  assign pht_1_7_MPORT_978_mask = 1'h1;
  assign pht_1_7_MPORT_978_en = reset;
  assign pht_1_7_MPORT_980_data = 1'h0;
  assign pht_1_7_MPORT_980_addr = 6'h12;
  assign pht_1_7_MPORT_980_mask = 1'h1;
  assign pht_1_7_MPORT_980_en = reset;
  assign pht_1_7_MPORT_982_data = 1'h0;
  assign pht_1_7_MPORT_982_addr = 6'h13;
  assign pht_1_7_MPORT_982_mask = 1'h1;
  assign pht_1_7_MPORT_982_en = reset;
  assign pht_1_7_MPORT_984_data = 1'h0;
  assign pht_1_7_MPORT_984_addr = 6'h14;
  assign pht_1_7_MPORT_984_mask = 1'h1;
  assign pht_1_7_MPORT_984_en = reset;
  assign pht_1_7_MPORT_986_data = 1'h0;
  assign pht_1_7_MPORT_986_addr = 6'h15;
  assign pht_1_7_MPORT_986_mask = 1'h1;
  assign pht_1_7_MPORT_986_en = reset;
  assign pht_1_7_MPORT_988_data = 1'h0;
  assign pht_1_7_MPORT_988_addr = 6'h16;
  assign pht_1_7_MPORT_988_mask = 1'h1;
  assign pht_1_7_MPORT_988_en = reset;
  assign pht_1_7_MPORT_990_data = 1'h0;
  assign pht_1_7_MPORT_990_addr = 6'h17;
  assign pht_1_7_MPORT_990_mask = 1'h1;
  assign pht_1_7_MPORT_990_en = reset;
  assign pht_1_7_MPORT_992_data = 1'h0;
  assign pht_1_7_MPORT_992_addr = 6'h18;
  assign pht_1_7_MPORT_992_mask = 1'h1;
  assign pht_1_7_MPORT_992_en = reset;
  assign pht_1_7_MPORT_994_data = 1'h0;
  assign pht_1_7_MPORT_994_addr = 6'h19;
  assign pht_1_7_MPORT_994_mask = 1'h1;
  assign pht_1_7_MPORT_994_en = reset;
  assign pht_1_7_MPORT_996_data = 1'h0;
  assign pht_1_7_MPORT_996_addr = 6'h1a;
  assign pht_1_7_MPORT_996_mask = 1'h1;
  assign pht_1_7_MPORT_996_en = reset;
  assign pht_1_7_MPORT_998_data = 1'h0;
  assign pht_1_7_MPORT_998_addr = 6'h1b;
  assign pht_1_7_MPORT_998_mask = 1'h1;
  assign pht_1_7_MPORT_998_en = reset;
  assign pht_1_7_MPORT_1000_data = 1'h0;
  assign pht_1_7_MPORT_1000_addr = 6'h1c;
  assign pht_1_7_MPORT_1000_mask = 1'h1;
  assign pht_1_7_MPORT_1000_en = reset;
  assign pht_1_7_MPORT_1002_data = 1'h0;
  assign pht_1_7_MPORT_1002_addr = 6'h1d;
  assign pht_1_7_MPORT_1002_mask = 1'h1;
  assign pht_1_7_MPORT_1002_en = reset;
  assign pht_1_7_MPORT_1004_data = 1'h0;
  assign pht_1_7_MPORT_1004_addr = 6'h1e;
  assign pht_1_7_MPORT_1004_mask = 1'h1;
  assign pht_1_7_MPORT_1004_en = reset;
  assign pht_1_7_MPORT_1006_data = 1'h0;
  assign pht_1_7_MPORT_1006_addr = 6'h1f;
  assign pht_1_7_MPORT_1006_mask = 1'h1;
  assign pht_1_7_MPORT_1006_en = reset;
  assign pht_1_7_MPORT_1008_data = 1'h0;
  assign pht_1_7_MPORT_1008_addr = 6'h20;
  assign pht_1_7_MPORT_1008_mask = 1'h1;
  assign pht_1_7_MPORT_1008_en = reset;
  assign pht_1_7_MPORT_1010_data = 1'h0;
  assign pht_1_7_MPORT_1010_addr = 6'h21;
  assign pht_1_7_MPORT_1010_mask = 1'h1;
  assign pht_1_7_MPORT_1010_en = reset;
  assign pht_1_7_MPORT_1012_data = 1'h0;
  assign pht_1_7_MPORT_1012_addr = 6'h22;
  assign pht_1_7_MPORT_1012_mask = 1'h1;
  assign pht_1_7_MPORT_1012_en = reset;
  assign pht_1_7_MPORT_1014_data = 1'h0;
  assign pht_1_7_MPORT_1014_addr = 6'h23;
  assign pht_1_7_MPORT_1014_mask = 1'h1;
  assign pht_1_7_MPORT_1014_en = reset;
  assign pht_1_7_MPORT_1016_data = 1'h0;
  assign pht_1_7_MPORT_1016_addr = 6'h24;
  assign pht_1_7_MPORT_1016_mask = 1'h1;
  assign pht_1_7_MPORT_1016_en = reset;
  assign pht_1_7_MPORT_1018_data = 1'h0;
  assign pht_1_7_MPORT_1018_addr = 6'h25;
  assign pht_1_7_MPORT_1018_mask = 1'h1;
  assign pht_1_7_MPORT_1018_en = reset;
  assign pht_1_7_MPORT_1020_data = 1'h0;
  assign pht_1_7_MPORT_1020_addr = 6'h26;
  assign pht_1_7_MPORT_1020_mask = 1'h1;
  assign pht_1_7_MPORT_1020_en = reset;
  assign pht_1_7_MPORT_1022_data = 1'h0;
  assign pht_1_7_MPORT_1022_addr = 6'h27;
  assign pht_1_7_MPORT_1022_mask = 1'h1;
  assign pht_1_7_MPORT_1022_en = reset;
  assign pht_1_7_MPORT_1024_data = 1'h0;
  assign pht_1_7_MPORT_1024_addr = 6'h28;
  assign pht_1_7_MPORT_1024_mask = 1'h1;
  assign pht_1_7_MPORT_1024_en = reset;
  assign pht_1_7_MPORT_1026_data = 1'h0;
  assign pht_1_7_MPORT_1026_addr = 6'h29;
  assign pht_1_7_MPORT_1026_mask = 1'h1;
  assign pht_1_7_MPORT_1026_en = reset;
  assign pht_1_7_MPORT_1028_data = 1'h0;
  assign pht_1_7_MPORT_1028_addr = 6'h2a;
  assign pht_1_7_MPORT_1028_mask = 1'h1;
  assign pht_1_7_MPORT_1028_en = reset;
  assign pht_1_7_MPORT_1030_data = 1'h0;
  assign pht_1_7_MPORT_1030_addr = 6'h2b;
  assign pht_1_7_MPORT_1030_mask = 1'h1;
  assign pht_1_7_MPORT_1030_en = reset;
  assign pht_1_7_MPORT_1032_data = 1'h0;
  assign pht_1_7_MPORT_1032_addr = 6'h2c;
  assign pht_1_7_MPORT_1032_mask = 1'h1;
  assign pht_1_7_MPORT_1032_en = reset;
  assign pht_1_7_MPORT_1034_data = 1'h0;
  assign pht_1_7_MPORT_1034_addr = 6'h2d;
  assign pht_1_7_MPORT_1034_mask = 1'h1;
  assign pht_1_7_MPORT_1034_en = reset;
  assign pht_1_7_MPORT_1036_data = 1'h0;
  assign pht_1_7_MPORT_1036_addr = 6'h2e;
  assign pht_1_7_MPORT_1036_mask = 1'h1;
  assign pht_1_7_MPORT_1036_en = reset;
  assign pht_1_7_MPORT_1038_data = 1'h0;
  assign pht_1_7_MPORT_1038_addr = 6'h2f;
  assign pht_1_7_MPORT_1038_mask = 1'h1;
  assign pht_1_7_MPORT_1038_en = reset;
  assign pht_1_7_MPORT_1040_data = 1'h0;
  assign pht_1_7_MPORT_1040_addr = 6'h30;
  assign pht_1_7_MPORT_1040_mask = 1'h1;
  assign pht_1_7_MPORT_1040_en = reset;
  assign pht_1_7_MPORT_1042_data = 1'h0;
  assign pht_1_7_MPORT_1042_addr = 6'h31;
  assign pht_1_7_MPORT_1042_mask = 1'h1;
  assign pht_1_7_MPORT_1042_en = reset;
  assign pht_1_7_MPORT_1044_data = 1'h0;
  assign pht_1_7_MPORT_1044_addr = 6'h32;
  assign pht_1_7_MPORT_1044_mask = 1'h1;
  assign pht_1_7_MPORT_1044_en = reset;
  assign pht_1_7_MPORT_1046_data = 1'h0;
  assign pht_1_7_MPORT_1046_addr = 6'h33;
  assign pht_1_7_MPORT_1046_mask = 1'h1;
  assign pht_1_7_MPORT_1046_en = reset;
  assign pht_1_7_MPORT_1048_data = 1'h0;
  assign pht_1_7_MPORT_1048_addr = 6'h34;
  assign pht_1_7_MPORT_1048_mask = 1'h1;
  assign pht_1_7_MPORT_1048_en = reset;
  assign pht_1_7_MPORT_1050_data = 1'h0;
  assign pht_1_7_MPORT_1050_addr = 6'h35;
  assign pht_1_7_MPORT_1050_mask = 1'h1;
  assign pht_1_7_MPORT_1050_en = reset;
  assign pht_1_7_MPORT_1052_data = 1'h0;
  assign pht_1_7_MPORT_1052_addr = 6'h36;
  assign pht_1_7_MPORT_1052_mask = 1'h1;
  assign pht_1_7_MPORT_1052_en = reset;
  assign pht_1_7_MPORT_1054_data = 1'h0;
  assign pht_1_7_MPORT_1054_addr = 6'h37;
  assign pht_1_7_MPORT_1054_mask = 1'h1;
  assign pht_1_7_MPORT_1054_en = reset;
  assign pht_1_7_MPORT_1056_data = 1'h0;
  assign pht_1_7_MPORT_1056_addr = 6'h38;
  assign pht_1_7_MPORT_1056_mask = 1'h1;
  assign pht_1_7_MPORT_1056_en = reset;
  assign pht_1_7_MPORT_1058_data = 1'h0;
  assign pht_1_7_MPORT_1058_addr = 6'h39;
  assign pht_1_7_MPORT_1058_mask = 1'h1;
  assign pht_1_7_MPORT_1058_en = reset;
  assign pht_1_7_MPORT_1060_data = 1'h0;
  assign pht_1_7_MPORT_1060_addr = 6'h3a;
  assign pht_1_7_MPORT_1060_mask = 1'h1;
  assign pht_1_7_MPORT_1060_en = reset;
  assign pht_1_7_MPORT_1062_data = 1'h0;
  assign pht_1_7_MPORT_1062_addr = 6'h3b;
  assign pht_1_7_MPORT_1062_mask = 1'h1;
  assign pht_1_7_MPORT_1062_en = reset;
  assign pht_1_7_MPORT_1064_data = 1'h0;
  assign pht_1_7_MPORT_1064_addr = 6'h3c;
  assign pht_1_7_MPORT_1064_mask = 1'h1;
  assign pht_1_7_MPORT_1064_en = reset;
  assign pht_1_7_MPORT_1066_data = 1'h0;
  assign pht_1_7_MPORT_1066_addr = 6'h3d;
  assign pht_1_7_MPORT_1066_mask = 1'h1;
  assign pht_1_7_MPORT_1066_en = reset;
  assign pht_1_7_MPORT_1068_data = 1'h0;
  assign pht_1_7_MPORT_1068_addr = 6'h3e;
  assign pht_1_7_MPORT_1068_mask = 1'h1;
  assign pht_1_7_MPORT_1068_en = reset;
  assign pht_1_7_MPORT_1070_data = 1'h0;
  assign pht_1_7_MPORT_1070_addr = 6'h3f;
  assign pht_1_7_MPORT_1070_mask = 1'h1;
  assign pht_1_7_MPORT_1070_en = reset;
//   assign pht_0_0_MPORT_17_en = pht_0_0_MPORT_17_en_pipe_0;
  assign pht_0_0_MPORT_17_addr = pht_0_0_MPORT_17_addr_pipe_0;
  assign pht_0_0_MPORT_17_data = pht_0_0[pht_0_0_MPORT_17_addr]; // @[PatternHistoryTable.scala 26:28]
  assign pht_0_0_MPORT_33_data = pht_wdata_w[0];
  assign pht_0_0_MPORT_33_addr = REG_32;
  assign pht_0_0_MPORT_33_mask = 1'h1;
  assign pht_0_0_MPORT_33_en = REG_29 & REG_30;
  assign pht_0_0_MPORT_49_data = 1'h0;
  assign pht_0_0_MPORT_49_addr = 6'h0;
  assign pht_0_0_MPORT_49_mask = 1'h1;
  assign pht_0_0_MPORT_49_en = reset;
  assign pht_0_0_MPORT_51_data = 1'h0;
  assign pht_0_0_MPORT_51_addr = 6'h1;
  assign pht_0_0_MPORT_51_mask = 1'h1;
  assign pht_0_0_MPORT_51_en = reset;
  assign pht_0_0_MPORT_53_data = 1'h0;
  assign pht_0_0_MPORT_53_addr = 6'h2;
  assign pht_0_0_MPORT_53_mask = 1'h1;
  assign pht_0_0_MPORT_53_en = reset;
  assign pht_0_0_MPORT_55_data = 1'h0;
  assign pht_0_0_MPORT_55_addr = 6'h3;
  assign pht_0_0_MPORT_55_mask = 1'h1;
  assign pht_0_0_MPORT_55_en = reset;
  assign pht_0_0_MPORT_57_data = 1'h0;
  assign pht_0_0_MPORT_57_addr = 6'h4;
  assign pht_0_0_MPORT_57_mask = 1'h1;
  assign pht_0_0_MPORT_57_en = reset;
  assign pht_0_0_MPORT_59_data = 1'h0;
  assign pht_0_0_MPORT_59_addr = 6'h5;
  assign pht_0_0_MPORT_59_mask = 1'h1;
  assign pht_0_0_MPORT_59_en = reset;
  assign pht_0_0_MPORT_61_data = 1'h0;
  assign pht_0_0_MPORT_61_addr = 6'h6;
  assign pht_0_0_MPORT_61_mask = 1'h1;
  assign pht_0_0_MPORT_61_en = reset;
  assign pht_0_0_MPORT_63_data = 1'h0;
  assign pht_0_0_MPORT_63_addr = 6'h7;
  assign pht_0_0_MPORT_63_mask = 1'h1;
  assign pht_0_0_MPORT_63_en = reset;
  assign pht_0_0_MPORT_65_data = 1'h0;
  assign pht_0_0_MPORT_65_addr = 6'h8;
  assign pht_0_0_MPORT_65_mask = 1'h1;
  assign pht_0_0_MPORT_65_en = reset;
  assign pht_0_0_MPORT_67_data = 1'h0;
  assign pht_0_0_MPORT_67_addr = 6'h9;
  assign pht_0_0_MPORT_67_mask = 1'h1;
  assign pht_0_0_MPORT_67_en = reset;
  assign pht_0_0_MPORT_69_data = 1'h0;
  assign pht_0_0_MPORT_69_addr = 6'ha;
  assign pht_0_0_MPORT_69_mask = 1'h1;
  assign pht_0_0_MPORT_69_en = reset;
  assign pht_0_0_MPORT_71_data = 1'h0;
  assign pht_0_0_MPORT_71_addr = 6'hb;
  assign pht_0_0_MPORT_71_mask = 1'h1;
  assign pht_0_0_MPORT_71_en = reset;
  assign pht_0_0_MPORT_73_data = 1'h0;
  assign pht_0_0_MPORT_73_addr = 6'hc;
  assign pht_0_0_MPORT_73_mask = 1'h1;
  assign pht_0_0_MPORT_73_en = reset;
  assign pht_0_0_MPORT_75_data = 1'h0;
  assign pht_0_0_MPORT_75_addr = 6'hd;
  assign pht_0_0_MPORT_75_mask = 1'h1;
  assign pht_0_0_MPORT_75_en = reset;
  assign pht_0_0_MPORT_77_data = 1'h0;
  assign pht_0_0_MPORT_77_addr = 6'he;
  assign pht_0_0_MPORT_77_mask = 1'h1;
  assign pht_0_0_MPORT_77_en = reset;
  assign pht_0_0_MPORT_79_data = 1'h0;
  assign pht_0_0_MPORT_79_addr = 6'hf;
  assign pht_0_0_MPORT_79_mask = 1'h1;
  assign pht_0_0_MPORT_79_en = reset;
  assign pht_0_0_MPORT_81_data = 1'h0;
  assign pht_0_0_MPORT_81_addr = 6'h10;
  assign pht_0_0_MPORT_81_mask = 1'h1;
  assign pht_0_0_MPORT_81_en = reset;
  assign pht_0_0_MPORT_83_data = 1'h0;
  assign pht_0_0_MPORT_83_addr = 6'h11;
  assign pht_0_0_MPORT_83_mask = 1'h1;
  assign pht_0_0_MPORT_83_en = reset;
  assign pht_0_0_MPORT_85_data = 1'h0;
  assign pht_0_0_MPORT_85_addr = 6'h12;
  assign pht_0_0_MPORT_85_mask = 1'h1;
  assign pht_0_0_MPORT_85_en = reset;
  assign pht_0_0_MPORT_87_data = 1'h0;
  assign pht_0_0_MPORT_87_addr = 6'h13;
  assign pht_0_0_MPORT_87_mask = 1'h1;
  assign pht_0_0_MPORT_87_en = reset;
  assign pht_0_0_MPORT_89_data = 1'h0;
  assign pht_0_0_MPORT_89_addr = 6'h14;
  assign pht_0_0_MPORT_89_mask = 1'h1;
  assign pht_0_0_MPORT_89_en = reset;
  assign pht_0_0_MPORT_91_data = 1'h0;
  assign pht_0_0_MPORT_91_addr = 6'h15;
  assign pht_0_0_MPORT_91_mask = 1'h1;
  assign pht_0_0_MPORT_91_en = reset;
  assign pht_0_0_MPORT_93_data = 1'h0;
  assign pht_0_0_MPORT_93_addr = 6'h16;
  assign pht_0_0_MPORT_93_mask = 1'h1;
  assign pht_0_0_MPORT_93_en = reset;
  assign pht_0_0_MPORT_95_data = 1'h0;
  assign pht_0_0_MPORT_95_addr = 6'h17;
  assign pht_0_0_MPORT_95_mask = 1'h1;
  assign pht_0_0_MPORT_95_en = reset;
  assign pht_0_0_MPORT_97_data = 1'h0;
  assign pht_0_0_MPORT_97_addr = 6'h18;
  assign pht_0_0_MPORT_97_mask = 1'h1;
  assign pht_0_0_MPORT_97_en = reset;
  assign pht_0_0_MPORT_99_data = 1'h0;
  assign pht_0_0_MPORT_99_addr = 6'h19;
  assign pht_0_0_MPORT_99_mask = 1'h1;
  assign pht_0_0_MPORT_99_en = reset;
  assign pht_0_0_MPORT_101_data = 1'h0;
  assign pht_0_0_MPORT_101_addr = 6'h1a;
  assign pht_0_0_MPORT_101_mask = 1'h1;
  assign pht_0_0_MPORT_101_en = reset;
  assign pht_0_0_MPORT_103_data = 1'h0;
  assign pht_0_0_MPORT_103_addr = 6'h1b;
  assign pht_0_0_MPORT_103_mask = 1'h1;
  assign pht_0_0_MPORT_103_en = reset;
  assign pht_0_0_MPORT_105_data = 1'h0;
  assign pht_0_0_MPORT_105_addr = 6'h1c;
  assign pht_0_0_MPORT_105_mask = 1'h1;
  assign pht_0_0_MPORT_105_en = reset;
  assign pht_0_0_MPORT_107_data = 1'h0;
  assign pht_0_0_MPORT_107_addr = 6'h1d;
  assign pht_0_0_MPORT_107_mask = 1'h1;
  assign pht_0_0_MPORT_107_en = reset;
  assign pht_0_0_MPORT_109_data = 1'h0;
  assign pht_0_0_MPORT_109_addr = 6'h1e;
  assign pht_0_0_MPORT_109_mask = 1'h1;
  assign pht_0_0_MPORT_109_en = reset;
  assign pht_0_0_MPORT_111_data = 1'h0;
  assign pht_0_0_MPORT_111_addr = 6'h1f;
  assign pht_0_0_MPORT_111_mask = 1'h1;
  assign pht_0_0_MPORT_111_en = reset;
  assign pht_0_0_MPORT_113_data = 1'h0;
  assign pht_0_0_MPORT_113_addr = 6'h20;
  assign pht_0_0_MPORT_113_mask = 1'h1;
  assign pht_0_0_MPORT_113_en = reset;
  assign pht_0_0_MPORT_115_data = 1'h0;
  assign pht_0_0_MPORT_115_addr = 6'h21;
  assign pht_0_0_MPORT_115_mask = 1'h1;
  assign pht_0_0_MPORT_115_en = reset;
  assign pht_0_0_MPORT_117_data = 1'h0;
  assign pht_0_0_MPORT_117_addr = 6'h22;
  assign pht_0_0_MPORT_117_mask = 1'h1;
  assign pht_0_0_MPORT_117_en = reset;
  assign pht_0_0_MPORT_119_data = 1'h0;
  assign pht_0_0_MPORT_119_addr = 6'h23;
  assign pht_0_0_MPORT_119_mask = 1'h1;
  assign pht_0_0_MPORT_119_en = reset;
  assign pht_0_0_MPORT_121_data = 1'h0;
  assign pht_0_0_MPORT_121_addr = 6'h24;
  assign pht_0_0_MPORT_121_mask = 1'h1;
  assign pht_0_0_MPORT_121_en = reset;
  assign pht_0_0_MPORT_123_data = 1'h0;
  assign pht_0_0_MPORT_123_addr = 6'h25;
  assign pht_0_0_MPORT_123_mask = 1'h1;
  assign pht_0_0_MPORT_123_en = reset;
  assign pht_0_0_MPORT_125_data = 1'h0;
  assign pht_0_0_MPORT_125_addr = 6'h26;
  assign pht_0_0_MPORT_125_mask = 1'h1;
  assign pht_0_0_MPORT_125_en = reset;
  assign pht_0_0_MPORT_127_data = 1'h0;
  assign pht_0_0_MPORT_127_addr = 6'h27;
  assign pht_0_0_MPORT_127_mask = 1'h1;
  assign pht_0_0_MPORT_127_en = reset;
  assign pht_0_0_MPORT_129_data = 1'h0;
  assign pht_0_0_MPORT_129_addr = 6'h28;
  assign pht_0_0_MPORT_129_mask = 1'h1;
  assign pht_0_0_MPORT_129_en = reset;
  assign pht_0_0_MPORT_131_data = 1'h0;
  assign pht_0_0_MPORT_131_addr = 6'h29;
  assign pht_0_0_MPORT_131_mask = 1'h1;
  assign pht_0_0_MPORT_131_en = reset;
  assign pht_0_0_MPORT_133_data = 1'h0;
  assign pht_0_0_MPORT_133_addr = 6'h2a;
  assign pht_0_0_MPORT_133_mask = 1'h1;
  assign pht_0_0_MPORT_133_en = reset;
  assign pht_0_0_MPORT_135_data = 1'h0;
  assign pht_0_0_MPORT_135_addr = 6'h2b;
  assign pht_0_0_MPORT_135_mask = 1'h1;
  assign pht_0_0_MPORT_135_en = reset;
  assign pht_0_0_MPORT_137_data = 1'h0;
  assign pht_0_0_MPORT_137_addr = 6'h2c;
  assign pht_0_0_MPORT_137_mask = 1'h1;
  assign pht_0_0_MPORT_137_en = reset;
  assign pht_0_0_MPORT_139_data = 1'h0;
  assign pht_0_0_MPORT_139_addr = 6'h2d;
  assign pht_0_0_MPORT_139_mask = 1'h1;
  assign pht_0_0_MPORT_139_en = reset;
  assign pht_0_0_MPORT_141_data = 1'h0;
  assign pht_0_0_MPORT_141_addr = 6'h2e;
  assign pht_0_0_MPORT_141_mask = 1'h1;
  assign pht_0_0_MPORT_141_en = reset;
  assign pht_0_0_MPORT_143_data = 1'h0;
  assign pht_0_0_MPORT_143_addr = 6'h2f;
  assign pht_0_0_MPORT_143_mask = 1'h1;
  assign pht_0_0_MPORT_143_en = reset;
  assign pht_0_0_MPORT_145_data = 1'h0;
  assign pht_0_0_MPORT_145_addr = 6'h30;
  assign pht_0_0_MPORT_145_mask = 1'h1;
  assign pht_0_0_MPORT_145_en = reset;
  assign pht_0_0_MPORT_147_data = 1'h0;
  assign pht_0_0_MPORT_147_addr = 6'h31;
  assign pht_0_0_MPORT_147_mask = 1'h1;
  assign pht_0_0_MPORT_147_en = reset;
  assign pht_0_0_MPORT_149_data = 1'h0;
  assign pht_0_0_MPORT_149_addr = 6'h32;
  assign pht_0_0_MPORT_149_mask = 1'h1;
  assign pht_0_0_MPORT_149_en = reset;
  assign pht_0_0_MPORT_151_data = 1'h0;
  assign pht_0_0_MPORT_151_addr = 6'h33;
  assign pht_0_0_MPORT_151_mask = 1'h1;
  assign pht_0_0_MPORT_151_en = reset;
  assign pht_0_0_MPORT_153_data = 1'h0;
  assign pht_0_0_MPORT_153_addr = 6'h34;
  assign pht_0_0_MPORT_153_mask = 1'h1;
  assign pht_0_0_MPORT_153_en = reset;
  assign pht_0_0_MPORT_155_data = 1'h0;
  assign pht_0_0_MPORT_155_addr = 6'h35;
  assign pht_0_0_MPORT_155_mask = 1'h1;
  assign pht_0_0_MPORT_155_en = reset;
  assign pht_0_0_MPORT_157_data = 1'h0;
  assign pht_0_0_MPORT_157_addr = 6'h36;
  assign pht_0_0_MPORT_157_mask = 1'h1;
  assign pht_0_0_MPORT_157_en = reset;
  assign pht_0_0_MPORT_159_data = 1'h0;
  assign pht_0_0_MPORT_159_addr = 6'h37;
  assign pht_0_0_MPORT_159_mask = 1'h1;
  assign pht_0_0_MPORT_159_en = reset;
  assign pht_0_0_MPORT_161_data = 1'h0;
  assign pht_0_0_MPORT_161_addr = 6'h38;
  assign pht_0_0_MPORT_161_mask = 1'h1;
  assign pht_0_0_MPORT_161_en = reset;
  assign pht_0_0_MPORT_163_data = 1'h0;
  assign pht_0_0_MPORT_163_addr = 6'h39;
  assign pht_0_0_MPORT_163_mask = 1'h1;
  assign pht_0_0_MPORT_163_en = reset;
  assign pht_0_0_MPORT_165_data = 1'h0;
  assign pht_0_0_MPORT_165_addr = 6'h3a;
  assign pht_0_0_MPORT_165_mask = 1'h1;
  assign pht_0_0_MPORT_165_en = reset;
  assign pht_0_0_MPORT_167_data = 1'h0;
  assign pht_0_0_MPORT_167_addr = 6'h3b;
  assign pht_0_0_MPORT_167_mask = 1'h1;
  assign pht_0_0_MPORT_167_en = reset;
  assign pht_0_0_MPORT_169_data = 1'h0;
  assign pht_0_0_MPORT_169_addr = 6'h3c;
  assign pht_0_0_MPORT_169_mask = 1'h1;
  assign pht_0_0_MPORT_169_en = reset;
  assign pht_0_0_MPORT_171_data = 1'h0;
  assign pht_0_0_MPORT_171_addr = 6'h3d;
  assign pht_0_0_MPORT_171_mask = 1'h1;
  assign pht_0_0_MPORT_171_en = reset;
  assign pht_0_0_MPORT_173_data = 1'h0;
  assign pht_0_0_MPORT_173_addr = 6'h3e;
  assign pht_0_0_MPORT_173_mask = 1'h1;
  assign pht_0_0_MPORT_173_en = reset;
  assign pht_0_0_MPORT_175_data = 1'h0;
  assign pht_0_0_MPORT_175_addr = 6'h3f;
  assign pht_0_0_MPORT_175_mask = 1'h1;
  assign pht_0_0_MPORT_175_en = reset;
//   assign pht_0_1_MPORT_19_en = pht_0_1_MPORT_19_en_pipe_0;
  assign pht_0_1_MPORT_19_addr = pht_0_1_MPORT_19_addr_pipe_0;
  assign pht_0_1_MPORT_19_data = pht_0_1[pht_0_1_MPORT_19_addr]; // @[PatternHistoryTable.scala 26:28]
  assign pht_0_1_MPORT_35_data = pht_wdata_w[0];
  assign pht_0_1_MPORT_35_addr = REG_35;
  assign pht_0_1_MPORT_35_mask = 1'h1;
  assign pht_0_1_MPORT_35_en = REG_29 & REG_33;
  assign pht_0_1_MPORT_177_data = 1'h0;
  assign pht_0_1_MPORT_177_addr = 6'h0;
  assign pht_0_1_MPORT_177_mask = 1'h1;
  assign pht_0_1_MPORT_177_en = reset;
  assign pht_0_1_MPORT_179_data = 1'h0;
  assign pht_0_1_MPORT_179_addr = 6'h1;
  assign pht_0_1_MPORT_179_mask = 1'h1;
  assign pht_0_1_MPORT_179_en = reset;
  assign pht_0_1_MPORT_181_data = 1'h0;
  assign pht_0_1_MPORT_181_addr = 6'h2;
  assign pht_0_1_MPORT_181_mask = 1'h1;
  assign pht_0_1_MPORT_181_en = reset;
  assign pht_0_1_MPORT_183_data = 1'h0;
  assign pht_0_1_MPORT_183_addr = 6'h3;
  assign pht_0_1_MPORT_183_mask = 1'h1;
  assign pht_0_1_MPORT_183_en = reset;
  assign pht_0_1_MPORT_185_data = 1'h0;
  assign pht_0_1_MPORT_185_addr = 6'h4;
  assign pht_0_1_MPORT_185_mask = 1'h1;
  assign pht_0_1_MPORT_185_en = reset;
  assign pht_0_1_MPORT_187_data = 1'h0;
  assign pht_0_1_MPORT_187_addr = 6'h5;
  assign pht_0_1_MPORT_187_mask = 1'h1;
  assign pht_0_1_MPORT_187_en = reset;
  assign pht_0_1_MPORT_189_data = 1'h0;
  assign pht_0_1_MPORT_189_addr = 6'h6;
  assign pht_0_1_MPORT_189_mask = 1'h1;
  assign pht_0_1_MPORT_189_en = reset;
  assign pht_0_1_MPORT_191_data = 1'h0;
  assign pht_0_1_MPORT_191_addr = 6'h7;
  assign pht_0_1_MPORT_191_mask = 1'h1;
  assign pht_0_1_MPORT_191_en = reset;
  assign pht_0_1_MPORT_193_data = 1'h0;
  assign pht_0_1_MPORT_193_addr = 6'h8;
  assign pht_0_1_MPORT_193_mask = 1'h1;
  assign pht_0_1_MPORT_193_en = reset;
  assign pht_0_1_MPORT_195_data = 1'h0;
  assign pht_0_1_MPORT_195_addr = 6'h9;
  assign pht_0_1_MPORT_195_mask = 1'h1;
  assign pht_0_1_MPORT_195_en = reset;
  assign pht_0_1_MPORT_197_data = 1'h0;
  assign pht_0_1_MPORT_197_addr = 6'ha;
  assign pht_0_1_MPORT_197_mask = 1'h1;
  assign pht_0_1_MPORT_197_en = reset;
  assign pht_0_1_MPORT_199_data = 1'h0;
  assign pht_0_1_MPORT_199_addr = 6'hb;
  assign pht_0_1_MPORT_199_mask = 1'h1;
  assign pht_0_1_MPORT_199_en = reset;
  assign pht_0_1_MPORT_201_data = 1'h0;
  assign pht_0_1_MPORT_201_addr = 6'hc;
  assign pht_0_1_MPORT_201_mask = 1'h1;
  assign pht_0_1_MPORT_201_en = reset;
  assign pht_0_1_MPORT_203_data = 1'h0;
  assign pht_0_1_MPORT_203_addr = 6'hd;
  assign pht_0_1_MPORT_203_mask = 1'h1;
  assign pht_0_1_MPORT_203_en = reset;
  assign pht_0_1_MPORT_205_data = 1'h0;
  assign pht_0_1_MPORT_205_addr = 6'he;
  assign pht_0_1_MPORT_205_mask = 1'h1;
  assign pht_0_1_MPORT_205_en = reset;
  assign pht_0_1_MPORT_207_data = 1'h0;
  assign pht_0_1_MPORT_207_addr = 6'hf;
  assign pht_0_1_MPORT_207_mask = 1'h1;
  assign pht_0_1_MPORT_207_en = reset;
  assign pht_0_1_MPORT_209_data = 1'h0;
  assign pht_0_1_MPORT_209_addr = 6'h10;
  assign pht_0_1_MPORT_209_mask = 1'h1;
  assign pht_0_1_MPORT_209_en = reset;
  assign pht_0_1_MPORT_211_data = 1'h0;
  assign pht_0_1_MPORT_211_addr = 6'h11;
  assign pht_0_1_MPORT_211_mask = 1'h1;
  assign pht_0_1_MPORT_211_en = reset;
  assign pht_0_1_MPORT_213_data = 1'h0;
  assign pht_0_1_MPORT_213_addr = 6'h12;
  assign pht_0_1_MPORT_213_mask = 1'h1;
  assign pht_0_1_MPORT_213_en = reset;
  assign pht_0_1_MPORT_215_data = 1'h0;
  assign pht_0_1_MPORT_215_addr = 6'h13;
  assign pht_0_1_MPORT_215_mask = 1'h1;
  assign pht_0_1_MPORT_215_en = reset;
  assign pht_0_1_MPORT_217_data = 1'h0;
  assign pht_0_1_MPORT_217_addr = 6'h14;
  assign pht_0_1_MPORT_217_mask = 1'h1;
  assign pht_0_1_MPORT_217_en = reset;
  assign pht_0_1_MPORT_219_data = 1'h0;
  assign pht_0_1_MPORT_219_addr = 6'h15;
  assign pht_0_1_MPORT_219_mask = 1'h1;
  assign pht_0_1_MPORT_219_en = reset;
  assign pht_0_1_MPORT_221_data = 1'h0;
  assign pht_0_1_MPORT_221_addr = 6'h16;
  assign pht_0_1_MPORT_221_mask = 1'h1;
  assign pht_0_1_MPORT_221_en = reset;
  assign pht_0_1_MPORT_223_data = 1'h0;
  assign pht_0_1_MPORT_223_addr = 6'h17;
  assign pht_0_1_MPORT_223_mask = 1'h1;
  assign pht_0_1_MPORT_223_en = reset;
  assign pht_0_1_MPORT_225_data = 1'h0;
  assign pht_0_1_MPORT_225_addr = 6'h18;
  assign pht_0_1_MPORT_225_mask = 1'h1;
  assign pht_0_1_MPORT_225_en = reset;
  assign pht_0_1_MPORT_227_data = 1'h0;
  assign pht_0_1_MPORT_227_addr = 6'h19;
  assign pht_0_1_MPORT_227_mask = 1'h1;
  assign pht_0_1_MPORT_227_en = reset;
  assign pht_0_1_MPORT_229_data = 1'h0;
  assign pht_0_1_MPORT_229_addr = 6'h1a;
  assign pht_0_1_MPORT_229_mask = 1'h1;
  assign pht_0_1_MPORT_229_en = reset;
  assign pht_0_1_MPORT_231_data = 1'h0;
  assign pht_0_1_MPORT_231_addr = 6'h1b;
  assign pht_0_1_MPORT_231_mask = 1'h1;
  assign pht_0_1_MPORT_231_en = reset;
  assign pht_0_1_MPORT_233_data = 1'h0;
  assign pht_0_1_MPORT_233_addr = 6'h1c;
  assign pht_0_1_MPORT_233_mask = 1'h1;
  assign pht_0_1_MPORT_233_en = reset;
  assign pht_0_1_MPORT_235_data = 1'h0;
  assign pht_0_1_MPORT_235_addr = 6'h1d;
  assign pht_0_1_MPORT_235_mask = 1'h1;
  assign pht_0_1_MPORT_235_en = reset;
  assign pht_0_1_MPORT_237_data = 1'h0;
  assign pht_0_1_MPORT_237_addr = 6'h1e;
  assign pht_0_1_MPORT_237_mask = 1'h1;
  assign pht_0_1_MPORT_237_en = reset;
  assign pht_0_1_MPORT_239_data = 1'h0;
  assign pht_0_1_MPORT_239_addr = 6'h1f;
  assign pht_0_1_MPORT_239_mask = 1'h1;
  assign pht_0_1_MPORT_239_en = reset;
  assign pht_0_1_MPORT_241_data = 1'h0;
  assign pht_0_1_MPORT_241_addr = 6'h20;
  assign pht_0_1_MPORT_241_mask = 1'h1;
  assign pht_0_1_MPORT_241_en = reset;
  assign pht_0_1_MPORT_243_data = 1'h0;
  assign pht_0_1_MPORT_243_addr = 6'h21;
  assign pht_0_1_MPORT_243_mask = 1'h1;
  assign pht_0_1_MPORT_243_en = reset;
  assign pht_0_1_MPORT_245_data = 1'h0;
  assign pht_0_1_MPORT_245_addr = 6'h22;
  assign pht_0_1_MPORT_245_mask = 1'h1;
  assign pht_0_1_MPORT_245_en = reset;
  assign pht_0_1_MPORT_247_data = 1'h0;
  assign pht_0_1_MPORT_247_addr = 6'h23;
  assign pht_0_1_MPORT_247_mask = 1'h1;
  assign pht_0_1_MPORT_247_en = reset;
  assign pht_0_1_MPORT_249_data = 1'h0;
  assign pht_0_1_MPORT_249_addr = 6'h24;
  assign pht_0_1_MPORT_249_mask = 1'h1;
  assign pht_0_1_MPORT_249_en = reset;
  assign pht_0_1_MPORT_251_data = 1'h0;
  assign pht_0_1_MPORT_251_addr = 6'h25;
  assign pht_0_1_MPORT_251_mask = 1'h1;
  assign pht_0_1_MPORT_251_en = reset;
  assign pht_0_1_MPORT_253_data = 1'h0;
  assign pht_0_1_MPORT_253_addr = 6'h26;
  assign pht_0_1_MPORT_253_mask = 1'h1;
  assign pht_0_1_MPORT_253_en = reset;
  assign pht_0_1_MPORT_255_data = 1'h0;
  assign pht_0_1_MPORT_255_addr = 6'h27;
  assign pht_0_1_MPORT_255_mask = 1'h1;
  assign pht_0_1_MPORT_255_en = reset;
  assign pht_0_1_MPORT_257_data = 1'h0;
  assign pht_0_1_MPORT_257_addr = 6'h28;
  assign pht_0_1_MPORT_257_mask = 1'h1;
  assign pht_0_1_MPORT_257_en = reset;
  assign pht_0_1_MPORT_259_data = 1'h0;
  assign pht_0_1_MPORT_259_addr = 6'h29;
  assign pht_0_1_MPORT_259_mask = 1'h1;
  assign pht_0_1_MPORT_259_en = reset;
  assign pht_0_1_MPORT_261_data = 1'h0;
  assign pht_0_1_MPORT_261_addr = 6'h2a;
  assign pht_0_1_MPORT_261_mask = 1'h1;
  assign pht_0_1_MPORT_261_en = reset;
  assign pht_0_1_MPORT_263_data = 1'h0;
  assign pht_0_1_MPORT_263_addr = 6'h2b;
  assign pht_0_1_MPORT_263_mask = 1'h1;
  assign pht_0_1_MPORT_263_en = reset;
  assign pht_0_1_MPORT_265_data = 1'h0;
  assign pht_0_1_MPORT_265_addr = 6'h2c;
  assign pht_0_1_MPORT_265_mask = 1'h1;
  assign pht_0_1_MPORT_265_en = reset;
  assign pht_0_1_MPORT_267_data = 1'h0;
  assign pht_0_1_MPORT_267_addr = 6'h2d;
  assign pht_0_1_MPORT_267_mask = 1'h1;
  assign pht_0_1_MPORT_267_en = reset;
  assign pht_0_1_MPORT_269_data = 1'h0;
  assign pht_0_1_MPORT_269_addr = 6'h2e;
  assign pht_0_1_MPORT_269_mask = 1'h1;
  assign pht_0_1_MPORT_269_en = reset;
  assign pht_0_1_MPORT_271_data = 1'h0;
  assign pht_0_1_MPORT_271_addr = 6'h2f;
  assign pht_0_1_MPORT_271_mask = 1'h1;
  assign pht_0_1_MPORT_271_en = reset;
  assign pht_0_1_MPORT_273_data = 1'h0;
  assign pht_0_1_MPORT_273_addr = 6'h30;
  assign pht_0_1_MPORT_273_mask = 1'h1;
  assign pht_0_1_MPORT_273_en = reset;
  assign pht_0_1_MPORT_275_data = 1'h0;
  assign pht_0_1_MPORT_275_addr = 6'h31;
  assign pht_0_1_MPORT_275_mask = 1'h1;
  assign pht_0_1_MPORT_275_en = reset;
  assign pht_0_1_MPORT_277_data = 1'h0;
  assign pht_0_1_MPORT_277_addr = 6'h32;
  assign pht_0_1_MPORT_277_mask = 1'h1;
  assign pht_0_1_MPORT_277_en = reset;
  assign pht_0_1_MPORT_279_data = 1'h0;
  assign pht_0_1_MPORT_279_addr = 6'h33;
  assign pht_0_1_MPORT_279_mask = 1'h1;
  assign pht_0_1_MPORT_279_en = reset;
  assign pht_0_1_MPORT_281_data = 1'h0;
  assign pht_0_1_MPORT_281_addr = 6'h34;
  assign pht_0_1_MPORT_281_mask = 1'h1;
  assign pht_0_1_MPORT_281_en = reset;
  assign pht_0_1_MPORT_283_data = 1'h0;
  assign pht_0_1_MPORT_283_addr = 6'h35;
  assign pht_0_1_MPORT_283_mask = 1'h1;
  assign pht_0_1_MPORT_283_en = reset;
  assign pht_0_1_MPORT_285_data = 1'h0;
  assign pht_0_1_MPORT_285_addr = 6'h36;
  assign pht_0_1_MPORT_285_mask = 1'h1;
  assign pht_0_1_MPORT_285_en = reset;
  assign pht_0_1_MPORT_287_data = 1'h0;
  assign pht_0_1_MPORT_287_addr = 6'h37;
  assign pht_0_1_MPORT_287_mask = 1'h1;
  assign pht_0_1_MPORT_287_en = reset;
  assign pht_0_1_MPORT_289_data = 1'h0;
  assign pht_0_1_MPORT_289_addr = 6'h38;
  assign pht_0_1_MPORT_289_mask = 1'h1;
  assign pht_0_1_MPORT_289_en = reset;
  assign pht_0_1_MPORT_291_data = 1'h0;
  assign pht_0_1_MPORT_291_addr = 6'h39;
  assign pht_0_1_MPORT_291_mask = 1'h1;
  assign pht_0_1_MPORT_291_en = reset;
  assign pht_0_1_MPORT_293_data = 1'h0;
  assign pht_0_1_MPORT_293_addr = 6'h3a;
  assign pht_0_1_MPORT_293_mask = 1'h1;
  assign pht_0_1_MPORT_293_en = reset;
  assign pht_0_1_MPORT_295_data = 1'h0;
  assign pht_0_1_MPORT_295_addr = 6'h3b;
  assign pht_0_1_MPORT_295_mask = 1'h1;
  assign pht_0_1_MPORT_295_en = reset;
  assign pht_0_1_MPORT_297_data = 1'h0;
  assign pht_0_1_MPORT_297_addr = 6'h3c;
  assign pht_0_1_MPORT_297_mask = 1'h1;
  assign pht_0_1_MPORT_297_en = reset;
  assign pht_0_1_MPORT_299_data = 1'h0;
  assign pht_0_1_MPORT_299_addr = 6'h3d;
  assign pht_0_1_MPORT_299_mask = 1'h1;
  assign pht_0_1_MPORT_299_en = reset;
  assign pht_0_1_MPORT_301_data = 1'h0;
  assign pht_0_1_MPORT_301_addr = 6'h3e;
  assign pht_0_1_MPORT_301_mask = 1'h1;
  assign pht_0_1_MPORT_301_en = reset;
  assign pht_0_1_MPORT_303_data = 1'h0;
  assign pht_0_1_MPORT_303_addr = 6'h3f;
  assign pht_0_1_MPORT_303_mask = 1'h1;
  assign pht_0_1_MPORT_303_en = reset;
//   assign pht_0_2_MPORT_21_en = pht_0_2_MPORT_21_en_pipe_0;
  assign pht_0_2_MPORT_21_addr = pht_0_2_MPORT_21_addr_pipe_0;
  assign pht_0_2_MPORT_21_data = pht_0_2[pht_0_2_MPORT_21_addr]; // @[PatternHistoryTable.scala 26:28]
  assign pht_0_2_MPORT_37_data = pht_wdata_w[0];
  assign pht_0_2_MPORT_37_addr = REG_38;
  assign pht_0_2_MPORT_37_mask = 1'h1;
  assign pht_0_2_MPORT_37_en = REG_29 & REG_36;
  assign pht_0_2_MPORT_305_data = 1'h0;
  assign pht_0_2_MPORT_305_addr = 6'h0;
  assign pht_0_2_MPORT_305_mask = 1'h1;
  assign pht_0_2_MPORT_305_en = reset;
  assign pht_0_2_MPORT_307_data = 1'h0;
  assign pht_0_2_MPORT_307_addr = 6'h1;
  assign pht_0_2_MPORT_307_mask = 1'h1;
  assign pht_0_2_MPORT_307_en = reset;
  assign pht_0_2_MPORT_309_data = 1'h0;
  assign pht_0_2_MPORT_309_addr = 6'h2;
  assign pht_0_2_MPORT_309_mask = 1'h1;
  assign pht_0_2_MPORT_309_en = reset;
  assign pht_0_2_MPORT_311_data = 1'h0;
  assign pht_0_2_MPORT_311_addr = 6'h3;
  assign pht_0_2_MPORT_311_mask = 1'h1;
  assign pht_0_2_MPORT_311_en = reset;
  assign pht_0_2_MPORT_313_data = 1'h0;
  assign pht_0_2_MPORT_313_addr = 6'h4;
  assign pht_0_2_MPORT_313_mask = 1'h1;
  assign pht_0_2_MPORT_313_en = reset;
  assign pht_0_2_MPORT_315_data = 1'h0;
  assign pht_0_2_MPORT_315_addr = 6'h5;
  assign pht_0_2_MPORT_315_mask = 1'h1;
  assign pht_0_2_MPORT_315_en = reset;
  assign pht_0_2_MPORT_317_data = 1'h0;
  assign pht_0_2_MPORT_317_addr = 6'h6;
  assign pht_0_2_MPORT_317_mask = 1'h1;
  assign pht_0_2_MPORT_317_en = reset;
  assign pht_0_2_MPORT_319_data = 1'h0;
  assign pht_0_2_MPORT_319_addr = 6'h7;
  assign pht_0_2_MPORT_319_mask = 1'h1;
  assign pht_0_2_MPORT_319_en = reset;
  assign pht_0_2_MPORT_321_data = 1'h0;
  assign pht_0_2_MPORT_321_addr = 6'h8;
  assign pht_0_2_MPORT_321_mask = 1'h1;
  assign pht_0_2_MPORT_321_en = reset;
  assign pht_0_2_MPORT_323_data = 1'h0;
  assign pht_0_2_MPORT_323_addr = 6'h9;
  assign pht_0_2_MPORT_323_mask = 1'h1;
  assign pht_0_2_MPORT_323_en = reset;
  assign pht_0_2_MPORT_325_data = 1'h0;
  assign pht_0_2_MPORT_325_addr = 6'ha;
  assign pht_0_2_MPORT_325_mask = 1'h1;
  assign pht_0_2_MPORT_325_en = reset;
  assign pht_0_2_MPORT_327_data = 1'h0;
  assign pht_0_2_MPORT_327_addr = 6'hb;
  assign pht_0_2_MPORT_327_mask = 1'h1;
  assign pht_0_2_MPORT_327_en = reset;
  assign pht_0_2_MPORT_329_data = 1'h0;
  assign pht_0_2_MPORT_329_addr = 6'hc;
  assign pht_0_2_MPORT_329_mask = 1'h1;
  assign pht_0_2_MPORT_329_en = reset;
  assign pht_0_2_MPORT_331_data = 1'h0;
  assign pht_0_2_MPORT_331_addr = 6'hd;
  assign pht_0_2_MPORT_331_mask = 1'h1;
  assign pht_0_2_MPORT_331_en = reset;
  assign pht_0_2_MPORT_333_data = 1'h0;
  assign pht_0_2_MPORT_333_addr = 6'he;
  assign pht_0_2_MPORT_333_mask = 1'h1;
  assign pht_0_2_MPORT_333_en = reset;
  assign pht_0_2_MPORT_335_data = 1'h0;
  assign pht_0_2_MPORT_335_addr = 6'hf;
  assign pht_0_2_MPORT_335_mask = 1'h1;
  assign pht_0_2_MPORT_335_en = reset;
  assign pht_0_2_MPORT_337_data = 1'h0;
  assign pht_0_2_MPORT_337_addr = 6'h10;
  assign pht_0_2_MPORT_337_mask = 1'h1;
  assign pht_0_2_MPORT_337_en = reset;
  assign pht_0_2_MPORT_339_data = 1'h0;
  assign pht_0_2_MPORT_339_addr = 6'h11;
  assign pht_0_2_MPORT_339_mask = 1'h1;
  assign pht_0_2_MPORT_339_en = reset;
  assign pht_0_2_MPORT_341_data = 1'h0;
  assign pht_0_2_MPORT_341_addr = 6'h12;
  assign pht_0_2_MPORT_341_mask = 1'h1;
  assign pht_0_2_MPORT_341_en = reset;
  assign pht_0_2_MPORT_343_data = 1'h0;
  assign pht_0_2_MPORT_343_addr = 6'h13;
  assign pht_0_2_MPORT_343_mask = 1'h1;
  assign pht_0_2_MPORT_343_en = reset;
  assign pht_0_2_MPORT_345_data = 1'h0;
  assign pht_0_2_MPORT_345_addr = 6'h14;
  assign pht_0_2_MPORT_345_mask = 1'h1;
  assign pht_0_2_MPORT_345_en = reset;
  assign pht_0_2_MPORT_347_data = 1'h0;
  assign pht_0_2_MPORT_347_addr = 6'h15;
  assign pht_0_2_MPORT_347_mask = 1'h1;
  assign pht_0_2_MPORT_347_en = reset;
  assign pht_0_2_MPORT_349_data = 1'h0;
  assign pht_0_2_MPORT_349_addr = 6'h16;
  assign pht_0_2_MPORT_349_mask = 1'h1;
  assign pht_0_2_MPORT_349_en = reset;
  assign pht_0_2_MPORT_351_data = 1'h0;
  assign pht_0_2_MPORT_351_addr = 6'h17;
  assign pht_0_2_MPORT_351_mask = 1'h1;
  assign pht_0_2_MPORT_351_en = reset;
  assign pht_0_2_MPORT_353_data = 1'h0;
  assign pht_0_2_MPORT_353_addr = 6'h18;
  assign pht_0_2_MPORT_353_mask = 1'h1;
  assign pht_0_2_MPORT_353_en = reset;
  assign pht_0_2_MPORT_355_data = 1'h0;
  assign pht_0_2_MPORT_355_addr = 6'h19;
  assign pht_0_2_MPORT_355_mask = 1'h1;
  assign pht_0_2_MPORT_355_en = reset;
  assign pht_0_2_MPORT_357_data = 1'h0;
  assign pht_0_2_MPORT_357_addr = 6'h1a;
  assign pht_0_2_MPORT_357_mask = 1'h1;
  assign pht_0_2_MPORT_357_en = reset;
  assign pht_0_2_MPORT_359_data = 1'h0;
  assign pht_0_2_MPORT_359_addr = 6'h1b;
  assign pht_0_2_MPORT_359_mask = 1'h1;
  assign pht_0_2_MPORT_359_en = reset;
  assign pht_0_2_MPORT_361_data = 1'h0;
  assign pht_0_2_MPORT_361_addr = 6'h1c;
  assign pht_0_2_MPORT_361_mask = 1'h1;
  assign pht_0_2_MPORT_361_en = reset;
  assign pht_0_2_MPORT_363_data = 1'h0;
  assign pht_0_2_MPORT_363_addr = 6'h1d;
  assign pht_0_2_MPORT_363_mask = 1'h1;
  assign pht_0_2_MPORT_363_en = reset;
  assign pht_0_2_MPORT_365_data = 1'h0;
  assign pht_0_2_MPORT_365_addr = 6'h1e;
  assign pht_0_2_MPORT_365_mask = 1'h1;
  assign pht_0_2_MPORT_365_en = reset;
  assign pht_0_2_MPORT_367_data = 1'h0;
  assign pht_0_2_MPORT_367_addr = 6'h1f;
  assign pht_0_2_MPORT_367_mask = 1'h1;
  assign pht_0_2_MPORT_367_en = reset;
  assign pht_0_2_MPORT_369_data = 1'h0;
  assign pht_0_2_MPORT_369_addr = 6'h20;
  assign pht_0_2_MPORT_369_mask = 1'h1;
  assign pht_0_2_MPORT_369_en = reset;
  assign pht_0_2_MPORT_371_data = 1'h0;
  assign pht_0_2_MPORT_371_addr = 6'h21;
  assign pht_0_2_MPORT_371_mask = 1'h1;
  assign pht_0_2_MPORT_371_en = reset;
  assign pht_0_2_MPORT_373_data = 1'h0;
  assign pht_0_2_MPORT_373_addr = 6'h22;
  assign pht_0_2_MPORT_373_mask = 1'h1;
  assign pht_0_2_MPORT_373_en = reset;
  assign pht_0_2_MPORT_375_data = 1'h0;
  assign pht_0_2_MPORT_375_addr = 6'h23;
  assign pht_0_2_MPORT_375_mask = 1'h1;
  assign pht_0_2_MPORT_375_en = reset;
  assign pht_0_2_MPORT_377_data = 1'h0;
  assign pht_0_2_MPORT_377_addr = 6'h24;
  assign pht_0_2_MPORT_377_mask = 1'h1;
  assign pht_0_2_MPORT_377_en = reset;
  assign pht_0_2_MPORT_379_data = 1'h0;
  assign pht_0_2_MPORT_379_addr = 6'h25;
  assign pht_0_2_MPORT_379_mask = 1'h1;
  assign pht_0_2_MPORT_379_en = reset;
  assign pht_0_2_MPORT_381_data = 1'h0;
  assign pht_0_2_MPORT_381_addr = 6'h26;
  assign pht_0_2_MPORT_381_mask = 1'h1;
  assign pht_0_2_MPORT_381_en = reset;
  assign pht_0_2_MPORT_383_data = 1'h0;
  assign pht_0_2_MPORT_383_addr = 6'h27;
  assign pht_0_2_MPORT_383_mask = 1'h1;
  assign pht_0_2_MPORT_383_en = reset;
  assign pht_0_2_MPORT_385_data = 1'h0;
  assign pht_0_2_MPORT_385_addr = 6'h28;
  assign pht_0_2_MPORT_385_mask = 1'h1;
  assign pht_0_2_MPORT_385_en = reset;
  assign pht_0_2_MPORT_387_data = 1'h0;
  assign pht_0_2_MPORT_387_addr = 6'h29;
  assign pht_0_2_MPORT_387_mask = 1'h1;
  assign pht_0_2_MPORT_387_en = reset;
  assign pht_0_2_MPORT_389_data = 1'h0;
  assign pht_0_2_MPORT_389_addr = 6'h2a;
  assign pht_0_2_MPORT_389_mask = 1'h1;
  assign pht_0_2_MPORT_389_en = reset;
  assign pht_0_2_MPORT_391_data = 1'h0;
  assign pht_0_2_MPORT_391_addr = 6'h2b;
  assign pht_0_2_MPORT_391_mask = 1'h1;
  assign pht_0_2_MPORT_391_en = reset;
  assign pht_0_2_MPORT_393_data = 1'h0;
  assign pht_0_2_MPORT_393_addr = 6'h2c;
  assign pht_0_2_MPORT_393_mask = 1'h1;
  assign pht_0_2_MPORT_393_en = reset;
  assign pht_0_2_MPORT_395_data = 1'h0;
  assign pht_0_2_MPORT_395_addr = 6'h2d;
  assign pht_0_2_MPORT_395_mask = 1'h1;
  assign pht_0_2_MPORT_395_en = reset;
  assign pht_0_2_MPORT_397_data = 1'h0;
  assign pht_0_2_MPORT_397_addr = 6'h2e;
  assign pht_0_2_MPORT_397_mask = 1'h1;
  assign pht_0_2_MPORT_397_en = reset;
  assign pht_0_2_MPORT_399_data = 1'h0;
  assign pht_0_2_MPORT_399_addr = 6'h2f;
  assign pht_0_2_MPORT_399_mask = 1'h1;
  assign pht_0_2_MPORT_399_en = reset;
  assign pht_0_2_MPORT_401_data = 1'h0;
  assign pht_0_2_MPORT_401_addr = 6'h30;
  assign pht_0_2_MPORT_401_mask = 1'h1;
  assign pht_0_2_MPORT_401_en = reset;
  assign pht_0_2_MPORT_403_data = 1'h0;
  assign pht_0_2_MPORT_403_addr = 6'h31;
  assign pht_0_2_MPORT_403_mask = 1'h1;
  assign pht_0_2_MPORT_403_en = reset;
  assign pht_0_2_MPORT_405_data = 1'h0;
  assign pht_0_2_MPORT_405_addr = 6'h32;
  assign pht_0_2_MPORT_405_mask = 1'h1;
  assign pht_0_2_MPORT_405_en = reset;
  assign pht_0_2_MPORT_407_data = 1'h0;
  assign pht_0_2_MPORT_407_addr = 6'h33;
  assign pht_0_2_MPORT_407_mask = 1'h1;
  assign pht_0_2_MPORT_407_en = reset;
  assign pht_0_2_MPORT_409_data = 1'h0;
  assign pht_0_2_MPORT_409_addr = 6'h34;
  assign pht_0_2_MPORT_409_mask = 1'h1;
  assign pht_0_2_MPORT_409_en = reset;
  assign pht_0_2_MPORT_411_data = 1'h0;
  assign pht_0_2_MPORT_411_addr = 6'h35;
  assign pht_0_2_MPORT_411_mask = 1'h1;
  assign pht_0_2_MPORT_411_en = reset;
  assign pht_0_2_MPORT_413_data = 1'h0;
  assign pht_0_2_MPORT_413_addr = 6'h36;
  assign pht_0_2_MPORT_413_mask = 1'h1;
  assign pht_0_2_MPORT_413_en = reset;
  assign pht_0_2_MPORT_415_data = 1'h0;
  assign pht_0_2_MPORT_415_addr = 6'h37;
  assign pht_0_2_MPORT_415_mask = 1'h1;
  assign pht_0_2_MPORT_415_en = reset;
  assign pht_0_2_MPORT_417_data = 1'h0;
  assign pht_0_2_MPORT_417_addr = 6'h38;
  assign pht_0_2_MPORT_417_mask = 1'h1;
  assign pht_0_2_MPORT_417_en = reset;
  assign pht_0_2_MPORT_419_data = 1'h0;
  assign pht_0_2_MPORT_419_addr = 6'h39;
  assign pht_0_2_MPORT_419_mask = 1'h1;
  assign pht_0_2_MPORT_419_en = reset;
  assign pht_0_2_MPORT_421_data = 1'h0;
  assign pht_0_2_MPORT_421_addr = 6'h3a;
  assign pht_0_2_MPORT_421_mask = 1'h1;
  assign pht_0_2_MPORT_421_en = reset;
  assign pht_0_2_MPORT_423_data = 1'h0;
  assign pht_0_2_MPORT_423_addr = 6'h3b;
  assign pht_0_2_MPORT_423_mask = 1'h1;
  assign pht_0_2_MPORT_423_en = reset;
  assign pht_0_2_MPORT_425_data = 1'h0;
  assign pht_0_2_MPORT_425_addr = 6'h3c;
  assign pht_0_2_MPORT_425_mask = 1'h1;
  assign pht_0_2_MPORT_425_en = reset;
  assign pht_0_2_MPORT_427_data = 1'h0;
  assign pht_0_2_MPORT_427_addr = 6'h3d;
  assign pht_0_2_MPORT_427_mask = 1'h1;
  assign pht_0_2_MPORT_427_en = reset;
  assign pht_0_2_MPORT_429_data = 1'h0;
  assign pht_0_2_MPORT_429_addr = 6'h3e;
  assign pht_0_2_MPORT_429_mask = 1'h1;
  assign pht_0_2_MPORT_429_en = reset;
  assign pht_0_2_MPORT_431_data = 1'h0;
  assign pht_0_2_MPORT_431_addr = 6'h3f;
  assign pht_0_2_MPORT_431_mask = 1'h1;
  assign pht_0_2_MPORT_431_en = reset;
//   assign pht_0_3_MPORT_23_en = pht_0_3_MPORT_23_en_pipe_0;
  assign pht_0_3_MPORT_23_addr = pht_0_3_MPORT_23_addr_pipe_0;
  assign pht_0_3_MPORT_23_data = pht_0_3[pht_0_3_MPORT_23_addr]; // @[PatternHistoryTable.scala 26:28]
  assign pht_0_3_MPORT_39_data = pht_wdata_w[0];
  assign pht_0_3_MPORT_39_addr = REG_41;
  assign pht_0_3_MPORT_39_mask = 1'h1;
  assign pht_0_3_MPORT_39_en = REG_29 & REG_39;
  assign pht_0_3_MPORT_433_data = 1'h0;
  assign pht_0_3_MPORT_433_addr = 6'h0;
  assign pht_0_3_MPORT_433_mask = 1'h1;
  assign pht_0_3_MPORT_433_en = reset;
  assign pht_0_3_MPORT_435_data = 1'h0;
  assign pht_0_3_MPORT_435_addr = 6'h1;
  assign pht_0_3_MPORT_435_mask = 1'h1;
  assign pht_0_3_MPORT_435_en = reset;
  assign pht_0_3_MPORT_437_data = 1'h0;
  assign pht_0_3_MPORT_437_addr = 6'h2;
  assign pht_0_3_MPORT_437_mask = 1'h1;
  assign pht_0_3_MPORT_437_en = reset;
  assign pht_0_3_MPORT_439_data = 1'h0;
  assign pht_0_3_MPORT_439_addr = 6'h3;
  assign pht_0_3_MPORT_439_mask = 1'h1;
  assign pht_0_3_MPORT_439_en = reset;
  assign pht_0_3_MPORT_441_data = 1'h0;
  assign pht_0_3_MPORT_441_addr = 6'h4;
  assign pht_0_3_MPORT_441_mask = 1'h1;
  assign pht_0_3_MPORT_441_en = reset;
  assign pht_0_3_MPORT_443_data = 1'h0;
  assign pht_0_3_MPORT_443_addr = 6'h5;
  assign pht_0_3_MPORT_443_mask = 1'h1;
  assign pht_0_3_MPORT_443_en = reset;
  assign pht_0_3_MPORT_445_data = 1'h0;
  assign pht_0_3_MPORT_445_addr = 6'h6;
  assign pht_0_3_MPORT_445_mask = 1'h1;
  assign pht_0_3_MPORT_445_en = reset;
  assign pht_0_3_MPORT_447_data = 1'h0;
  assign pht_0_3_MPORT_447_addr = 6'h7;
  assign pht_0_3_MPORT_447_mask = 1'h1;
  assign pht_0_3_MPORT_447_en = reset;
  assign pht_0_3_MPORT_449_data = 1'h0;
  assign pht_0_3_MPORT_449_addr = 6'h8;
  assign pht_0_3_MPORT_449_mask = 1'h1;
  assign pht_0_3_MPORT_449_en = reset;
  assign pht_0_3_MPORT_451_data = 1'h0;
  assign pht_0_3_MPORT_451_addr = 6'h9;
  assign pht_0_3_MPORT_451_mask = 1'h1;
  assign pht_0_3_MPORT_451_en = reset;
  assign pht_0_3_MPORT_453_data = 1'h0;
  assign pht_0_3_MPORT_453_addr = 6'ha;
  assign pht_0_3_MPORT_453_mask = 1'h1;
  assign pht_0_3_MPORT_453_en = reset;
  assign pht_0_3_MPORT_455_data = 1'h0;
  assign pht_0_3_MPORT_455_addr = 6'hb;
  assign pht_0_3_MPORT_455_mask = 1'h1;
  assign pht_0_3_MPORT_455_en = reset;
  assign pht_0_3_MPORT_457_data = 1'h0;
  assign pht_0_3_MPORT_457_addr = 6'hc;
  assign pht_0_3_MPORT_457_mask = 1'h1;
  assign pht_0_3_MPORT_457_en = reset;
  assign pht_0_3_MPORT_459_data = 1'h0;
  assign pht_0_3_MPORT_459_addr = 6'hd;
  assign pht_0_3_MPORT_459_mask = 1'h1;
  assign pht_0_3_MPORT_459_en = reset;
  assign pht_0_3_MPORT_461_data = 1'h0;
  assign pht_0_3_MPORT_461_addr = 6'he;
  assign pht_0_3_MPORT_461_mask = 1'h1;
  assign pht_0_3_MPORT_461_en = reset;
  assign pht_0_3_MPORT_463_data = 1'h0;
  assign pht_0_3_MPORT_463_addr = 6'hf;
  assign pht_0_3_MPORT_463_mask = 1'h1;
  assign pht_0_3_MPORT_463_en = reset;
  assign pht_0_3_MPORT_465_data = 1'h0;
  assign pht_0_3_MPORT_465_addr = 6'h10;
  assign pht_0_3_MPORT_465_mask = 1'h1;
  assign pht_0_3_MPORT_465_en = reset;
  assign pht_0_3_MPORT_467_data = 1'h0;
  assign pht_0_3_MPORT_467_addr = 6'h11;
  assign pht_0_3_MPORT_467_mask = 1'h1;
  assign pht_0_3_MPORT_467_en = reset;
  assign pht_0_3_MPORT_469_data = 1'h0;
  assign pht_0_3_MPORT_469_addr = 6'h12;
  assign pht_0_3_MPORT_469_mask = 1'h1;
  assign pht_0_3_MPORT_469_en = reset;
  assign pht_0_3_MPORT_471_data = 1'h0;
  assign pht_0_3_MPORT_471_addr = 6'h13;
  assign pht_0_3_MPORT_471_mask = 1'h1;
  assign pht_0_3_MPORT_471_en = reset;
  assign pht_0_3_MPORT_473_data = 1'h0;
  assign pht_0_3_MPORT_473_addr = 6'h14;
  assign pht_0_3_MPORT_473_mask = 1'h1;
  assign pht_0_3_MPORT_473_en = reset;
  assign pht_0_3_MPORT_475_data = 1'h0;
  assign pht_0_3_MPORT_475_addr = 6'h15;
  assign pht_0_3_MPORT_475_mask = 1'h1;
  assign pht_0_3_MPORT_475_en = reset;
  assign pht_0_3_MPORT_477_data = 1'h0;
  assign pht_0_3_MPORT_477_addr = 6'h16;
  assign pht_0_3_MPORT_477_mask = 1'h1;
  assign pht_0_3_MPORT_477_en = reset;
  assign pht_0_3_MPORT_479_data = 1'h0;
  assign pht_0_3_MPORT_479_addr = 6'h17;
  assign pht_0_3_MPORT_479_mask = 1'h1;
  assign pht_0_3_MPORT_479_en = reset;
  assign pht_0_3_MPORT_481_data = 1'h0;
  assign pht_0_3_MPORT_481_addr = 6'h18;
  assign pht_0_3_MPORT_481_mask = 1'h1;
  assign pht_0_3_MPORT_481_en = reset;
  assign pht_0_3_MPORT_483_data = 1'h0;
  assign pht_0_3_MPORT_483_addr = 6'h19;
  assign pht_0_3_MPORT_483_mask = 1'h1;
  assign pht_0_3_MPORT_483_en = reset;
  assign pht_0_3_MPORT_485_data = 1'h0;
  assign pht_0_3_MPORT_485_addr = 6'h1a;
  assign pht_0_3_MPORT_485_mask = 1'h1;
  assign pht_0_3_MPORT_485_en = reset;
  assign pht_0_3_MPORT_487_data = 1'h0;
  assign pht_0_3_MPORT_487_addr = 6'h1b;
  assign pht_0_3_MPORT_487_mask = 1'h1;
  assign pht_0_3_MPORT_487_en = reset;
  assign pht_0_3_MPORT_489_data = 1'h0;
  assign pht_0_3_MPORT_489_addr = 6'h1c;
  assign pht_0_3_MPORT_489_mask = 1'h1;
  assign pht_0_3_MPORT_489_en = reset;
  assign pht_0_3_MPORT_491_data = 1'h0;
  assign pht_0_3_MPORT_491_addr = 6'h1d;
  assign pht_0_3_MPORT_491_mask = 1'h1;
  assign pht_0_3_MPORT_491_en = reset;
  assign pht_0_3_MPORT_493_data = 1'h0;
  assign pht_0_3_MPORT_493_addr = 6'h1e;
  assign pht_0_3_MPORT_493_mask = 1'h1;
  assign pht_0_3_MPORT_493_en = reset;
  assign pht_0_3_MPORT_495_data = 1'h0;
  assign pht_0_3_MPORT_495_addr = 6'h1f;
  assign pht_0_3_MPORT_495_mask = 1'h1;
  assign pht_0_3_MPORT_495_en = reset;
  assign pht_0_3_MPORT_497_data = 1'h0;
  assign pht_0_3_MPORT_497_addr = 6'h20;
  assign pht_0_3_MPORT_497_mask = 1'h1;
  assign pht_0_3_MPORT_497_en = reset;
  assign pht_0_3_MPORT_499_data = 1'h0;
  assign pht_0_3_MPORT_499_addr = 6'h21;
  assign pht_0_3_MPORT_499_mask = 1'h1;
  assign pht_0_3_MPORT_499_en = reset;
  assign pht_0_3_MPORT_501_data = 1'h0;
  assign pht_0_3_MPORT_501_addr = 6'h22;
  assign pht_0_3_MPORT_501_mask = 1'h1;
  assign pht_0_3_MPORT_501_en = reset;
  assign pht_0_3_MPORT_503_data = 1'h0;
  assign pht_0_3_MPORT_503_addr = 6'h23;
  assign pht_0_3_MPORT_503_mask = 1'h1;
  assign pht_0_3_MPORT_503_en = reset;
  assign pht_0_3_MPORT_505_data = 1'h0;
  assign pht_0_3_MPORT_505_addr = 6'h24;
  assign pht_0_3_MPORT_505_mask = 1'h1;
  assign pht_0_3_MPORT_505_en = reset;
  assign pht_0_3_MPORT_507_data = 1'h0;
  assign pht_0_3_MPORT_507_addr = 6'h25;
  assign pht_0_3_MPORT_507_mask = 1'h1;
  assign pht_0_3_MPORT_507_en = reset;
  assign pht_0_3_MPORT_509_data = 1'h0;
  assign pht_0_3_MPORT_509_addr = 6'h26;
  assign pht_0_3_MPORT_509_mask = 1'h1;
  assign pht_0_3_MPORT_509_en = reset;
  assign pht_0_3_MPORT_511_data = 1'h0;
  assign pht_0_3_MPORT_511_addr = 6'h27;
  assign pht_0_3_MPORT_511_mask = 1'h1;
  assign pht_0_3_MPORT_511_en = reset;
  assign pht_0_3_MPORT_513_data = 1'h0;
  assign pht_0_3_MPORT_513_addr = 6'h28;
  assign pht_0_3_MPORT_513_mask = 1'h1;
  assign pht_0_3_MPORT_513_en = reset;
  assign pht_0_3_MPORT_515_data = 1'h0;
  assign pht_0_3_MPORT_515_addr = 6'h29;
  assign pht_0_3_MPORT_515_mask = 1'h1;
  assign pht_0_3_MPORT_515_en = reset;
  assign pht_0_3_MPORT_517_data = 1'h0;
  assign pht_0_3_MPORT_517_addr = 6'h2a;
  assign pht_0_3_MPORT_517_mask = 1'h1;
  assign pht_0_3_MPORT_517_en = reset;
  assign pht_0_3_MPORT_519_data = 1'h0;
  assign pht_0_3_MPORT_519_addr = 6'h2b;
  assign pht_0_3_MPORT_519_mask = 1'h1;
  assign pht_0_3_MPORT_519_en = reset;
  assign pht_0_3_MPORT_521_data = 1'h0;
  assign pht_0_3_MPORT_521_addr = 6'h2c;
  assign pht_0_3_MPORT_521_mask = 1'h1;
  assign pht_0_3_MPORT_521_en = reset;
  assign pht_0_3_MPORT_523_data = 1'h0;
  assign pht_0_3_MPORT_523_addr = 6'h2d;
  assign pht_0_3_MPORT_523_mask = 1'h1;
  assign pht_0_3_MPORT_523_en = reset;
  assign pht_0_3_MPORT_525_data = 1'h0;
  assign pht_0_3_MPORT_525_addr = 6'h2e;
  assign pht_0_3_MPORT_525_mask = 1'h1;
  assign pht_0_3_MPORT_525_en = reset;
  assign pht_0_3_MPORT_527_data = 1'h0;
  assign pht_0_3_MPORT_527_addr = 6'h2f;
  assign pht_0_3_MPORT_527_mask = 1'h1;
  assign pht_0_3_MPORT_527_en = reset;
  assign pht_0_3_MPORT_529_data = 1'h0;
  assign pht_0_3_MPORT_529_addr = 6'h30;
  assign pht_0_3_MPORT_529_mask = 1'h1;
  assign pht_0_3_MPORT_529_en = reset;
  assign pht_0_3_MPORT_531_data = 1'h0;
  assign pht_0_3_MPORT_531_addr = 6'h31;
  assign pht_0_3_MPORT_531_mask = 1'h1;
  assign pht_0_3_MPORT_531_en = reset;
  assign pht_0_3_MPORT_533_data = 1'h0;
  assign pht_0_3_MPORT_533_addr = 6'h32;
  assign pht_0_3_MPORT_533_mask = 1'h1;
  assign pht_0_3_MPORT_533_en = reset;
  assign pht_0_3_MPORT_535_data = 1'h0;
  assign pht_0_3_MPORT_535_addr = 6'h33;
  assign pht_0_3_MPORT_535_mask = 1'h1;
  assign pht_0_3_MPORT_535_en = reset;
  assign pht_0_3_MPORT_537_data = 1'h0;
  assign pht_0_3_MPORT_537_addr = 6'h34;
  assign pht_0_3_MPORT_537_mask = 1'h1;
  assign pht_0_3_MPORT_537_en = reset;
  assign pht_0_3_MPORT_539_data = 1'h0;
  assign pht_0_3_MPORT_539_addr = 6'h35;
  assign pht_0_3_MPORT_539_mask = 1'h1;
  assign pht_0_3_MPORT_539_en = reset;
  assign pht_0_3_MPORT_541_data = 1'h0;
  assign pht_0_3_MPORT_541_addr = 6'h36;
  assign pht_0_3_MPORT_541_mask = 1'h1;
  assign pht_0_3_MPORT_541_en = reset;
  assign pht_0_3_MPORT_543_data = 1'h0;
  assign pht_0_3_MPORT_543_addr = 6'h37;
  assign pht_0_3_MPORT_543_mask = 1'h1;
  assign pht_0_3_MPORT_543_en = reset;
  assign pht_0_3_MPORT_545_data = 1'h0;
  assign pht_0_3_MPORT_545_addr = 6'h38;
  assign pht_0_3_MPORT_545_mask = 1'h1;
  assign pht_0_3_MPORT_545_en = reset;
  assign pht_0_3_MPORT_547_data = 1'h0;
  assign pht_0_3_MPORT_547_addr = 6'h39;
  assign pht_0_3_MPORT_547_mask = 1'h1;
  assign pht_0_3_MPORT_547_en = reset;
  assign pht_0_3_MPORT_549_data = 1'h0;
  assign pht_0_3_MPORT_549_addr = 6'h3a;
  assign pht_0_3_MPORT_549_mask = 1'h1;
  assign pht_0_3_MPORT_549_en = reset;
  assign pht_0_3_MPORT_551_data = 1'h0;
  assign pht_0_3_MPORT_551_addr = 6'h3b;
  assign pht_0_3_MPORT_551_mask = 1'h1;
  assign pht_0_3_MPORT_551_en = reset;
  assign pht_0_3_MPORT_553_data = 1'h0;
  assign pht_0_3_MPORT_553_addr = 6'h3c;
  assign pht_0_3_MPORT_553_mask = 1'h1;
  assign pht_0_3_MPORT_553_en = reset;
  assign pht_0_3_MPORT_555_data = 1'h0;
  assign pht_0_3_MPORT_555_addr = 6'h3d;
  assign pht_0_3_MPORT_555_mask = 1'h1;
  assign pht_0_3_MPORT_555_en = reset;
  assign pht_0_3_MPORT_557_data = 1'h0;
  assign pht_0_3_MPORT_557_addr = 6'h3e;
  assign pht_0_3_MPORT_557_mask = 1'h1;
  assign pht_0_3_MPORT_557_en = reset;
  assign pht_0_3_MPORT_559_data = 1'h0;
  assign pht_0_3_MPORT_559_addr = 6'h3f;
  assign pht_0_3_MPORT_559_mask = 1'h1;
  assign pht_0_3_MPORT_559_en = reset;
//   assign pht_0_4_MPORT_25_en = pht_0_4_MPORT_25_en_pipe_0;
  assign pht_0_4_MPORT_25_addr = pht_0_4_MPORT_25_addr_pipe_0;
  assign pht_0_4_MPORT_25_data = pht_0_4[pht_0_4_MPORT_25_addr]; // @[PatternHistoryTable.scala 26:28]
  assign pht_0_4_MPORT_41_data = pht_wdata_w[0];
  assign pht_0_4_MPORT_41_addr = REG_44;
  assign pht_0_4_MPORT_41_mask = 1'h1;
  assign pht_0_4_MPORT_41_en = REG_29 & REG_42;
  assign pht_0_4_MPORT_561_data = 1'h0;
  assign pht_0_4_MPORT_561_addr = 6'h0;
  assign pht_0_4_MPORT_561_mask = 1'h1;
  assign pht_0_4_MPORT_561_en = reset;
  assign pht_0_4_MPORT_563_data = 1'h0;
  assign pht_0_4_MPORT_563_addr = 6'h1;
  assign pht_0_4_MPORT_563_mask = 1'h1;
  assign pht_0_4_MPORT_563_en = reset;
  assign pht_0_4_MPORT_565_data = 1'h0;
  assign pht_0_4_MPORT_565_addr = 6'h2;
  assign pht_0_4_MPORT_565_mask = 1'h1;
  assign pht_0_4_MPORT_565_en = reset;
  assign pht_0_4_MPORT_567_data = 1'h0;
  assign pht_0_4_MPORT_567_addr = 6'h3;
  assign pht_0_4_MPORT_567_mask = 1'h1;
  assign pht_0_4_MPORT_567_en = reset;
  assign pht_0_4_MPORT_569_data = 1'h0;
  assign pht_0_4_MPORT_569_addr = 6'h4;
  assign pht_0_4_MPORT_569_mask = 1'h1;
  assign pht_0_4_MPORT_569_en = reset;
  assign pht_0_4_MPORT_571_data = 1'h0;
  assign pht_0_4_MPORT_571_addr = 6'h5;
  assign pht_0_4_MPORT_571_mask = 1'h1;
  assign pht_0_4_MPORT_571_en = reset;
  assign pht_0_4_MPORT_573_data = 1'h0;
  assign pht_0_4_MPORT_573_addr = 6'h6;
  assign pht_0_4_MPORT_573_mask = 1'h1;
  assign pht_0_4_MPORT_573_en = reset;
  assign pht_0_4_MPORT_575_data = 1'h0;
  assign pht_0_4_MPORT_575_addr = 6'h7;
  assign pht_0_4_MPORT_575_mask = 1'h1;
  assign pht_0_4_MPORT_575_en = reset;
  assign pht_0_4_MPORT_577_data = 1'h0;
  assign pht_0_4_MPORT_577_addr = 6'h8;
  assign pht_0_4_MPORT_577_mask = 1'h1;
  assign pht_0_4_MPORT_577_en = reset;
  assign pht_0_4_MPORT_579_data = 1'h0;
  assign pht_0_4_MPORT_579_addr = 6'h9;
  assign pht_0_4_MPORT_579_mask = 1'h1;
  assign pht_0_4_MPORT_579_en = reset;
  assign pht_0_4_MPORT_581_data = 1'h0;
  assign pht_0_4_MPORT_581_addr = 6'ha;
  assign pht_0_4_MPORT_581_mask = 1'h1;
  assign pht_0_4_MPORT_581_en = reset;
  assign pht_0_4_MPORT_583_data = 1'h0;
  assign pht_0_4_MPORT_583_addr = 6'hb;
  assign pht_0_4_MPORT_583_mask = 1'h1;
  assign pht_0_4_MPORT_583_en = reset;
  assign pht_0_4_MPORT_585_data = 1'h0;
  assign pht_0_4_MPORT_585_addr = 6'hc;
  assign pht_0_4_MPORT_585_mask = 1'h1;
  assign pht_0_4_MPORT_585_en = reset;
  assign pht_0_4_MPORT_587_data = 1'h0;
  assign pht_0_4_MPORT_587_addr = 6'hd;
  assign pht_0_4_MPORT_587_mask = 1'h1;
  assign pht_0_4_MPORT_587_en = reset;
  assign pht_0_4_MPORT_589_data = 1'h0;
  assign pht_0_4_MPORT_589_addr = 6'he;
  assign pht_0_4_MPORT_589_mask = 1'h1;
  assign pht_0_4_MPORT_589_en = reset;
  assign pht_0_4_MPORT_591_data = 1'h0;
  assign pht_0_4_MPORT_591_addr = 6'hf;
  assign pht_0_4_MPORT_591_mask = 1'h1;
  assign pht_0_4_MPORT_591_en = reset;
  assign pht_0_4_MPORT_593_data = 1'h0;
  assign pht_0_4_MPORT_593_addr = 6'h10;
  assign pht_0_4_MPORT_593_mask = 1'h1;
  assign pht_0_4_MPORT_593_en = reset;
  assign pht_0_4_MPORT_595_data = 1'h0;
  assign pht_0_4_MPORT_595_addr = 6'h11;
  assign pht_0_4_MPORT_595_mask = 1'h1;
  assign pht_0_4_MPORT_595_en = reset;
  assign pht_0_4_MPORT_597_data = 1'h0;
  assign pht_0_4_MPORT_597_addr = 6'h12;
  assign pht_0_4_MPORT_597_mask = 1'h1;
  assign pht_0_4_MPORT_597_en = reset;
  assign pht_0_4_MPORT_599_data = 1'h0;
  assign pht_0_4_MPORT_599_addr = 6'h13;
  assign pht_0_4_MPORT_599_mask = 1'h1;
  assign pht_0_4_MPORT_599_en = reset;
  assign pht_0_4_MPORT_601_data = 1'h0;
  assign pht_0_4_MPORT_601_addr = 6'h14;
  assign pht_0_4_MPORT_601_mask = 1'h1;
  assign pht_0_4_MPORT_601_en = reset;
  assign pht_0_4_MPORT_603_data = 1'h0;
  assign pht_0_4_MPORT_603_addr = 6'h15;
  assign pht_0_4_MPORT_603_mask = 1'h1;
  assign pht_0_4_MPORT_603_en = reset;
  assign pht_0_4_MPORT_605_data = 1'h0;
  assign pht_0_4_MPORT_605_addr = 6'h16;
  assign pht_0_4_MPORT_605_mask = 1'h1;
  assign pht_0_4_MPORT_605_en = reset;
  assign pht_0_4_MPORT_607_data = 1'h0;
  assign pht_0_4_MPORT_607_addr = 6'h17;
  assign pht_0_4_MPORT_607_mask = 1'h1;
  assign pht_0_4_MPORT_607_en = reset;
  assign pht_0_4_MPORT_609_data = 1'h0;
  assign pht_0_4_MPORT_609_addr = 6'h18;
  assign pht_0_4_MPORT_609_mask = 1'h1;
  assign pht_0_4_MPORT_609_en = reset;
  assign pht_0_4_MPORT_611_data = 1'h0;
  assign pht_0_4_MPORT_611_addr = 6'h19;
  assign pht_0_4_MPORT_611_mask = 1'h1;
  assign pht_0_4_MPORT_611_en = reset;
  assign pht_0_4_MPORT_613_data = 1'h0;
  assign pht_0_4_MPORT_613_addr = 6'h1a;
  assign pht_0_4_MPORT_613_mask = 1'h1;
  assign pht_0_4_MPORT_613_en = reset;
  assign pht_0_4_MPORT_615_data = 1'h0;
  assign pht_0_4_MPORT_615_addr = 6'h1b;
  assign pht_0_4_MPORT_615_mask = 1'h1;
  assign pht_0_4_MPORT_615_en = reset;
  assign pht_0_4_MPORT_617_data = 1'h0;
  assign pht_0_4_MPORT_617_addr = 6'h1c;
  assign pht_0_4_MPORT_617_mask = 1'h1;
  assign pht_0_4_MPORT_617_en = reset;
  assign pht_0_4_MPORT_619_data = 1'h0;
  assign pht_0_4_MPORT_619_addr = 6'h1d;
  assign pht_0_4_MPORT_619_mask = 1'h1;
  assign pht_0_4_MPORT_619_en = reset;
  assign pht_0_4_MPORT_621_data = 1'h0;
  assign pht_0_4_MPORT_621_addr = 6'h1e;
  assign pht_0_4_MPORT_621_mask = 1'h1;
  assign pht_0_4_MPORT_621_en = reset;
  assign pht_0_4_MPORT_623_data = 1'h0;
  assign pht_0_4_MPORT_623_addr = 6'h1f;
  assign pht_0_4_MPORT_623_mask = 1'h1;
  assign pht_0_4_MPORT_623_en = reset;
  assign pht_0_4_MPORT_625_data = 1'h0;
  assign pht_0_4_MPORT_625_addr = 6'h20;
  assign pht_0_4_MPORT_625_mask = 1'h1;
  assign pht_0_4_MPORT_625_en = reset;
  assign pht_0_4_MPORT_627_data = 1'h0;
  assign pht_0_4_MPORT_627_addr = 6'h21;
  assign pht_0_4_MPORT_627_mask = 1'h1;
  assign pht_0_4_MPORT_627_en = reset;
  assign pht_0_4_MPORT_629_data = 1'h0;
  assign pht_0_4_MPORT_629_addr = 6'h22;
  assign pht_0_4_MPORT_629_mask = 1'h1;
  assign pht_0_4_MPORT_629_en = reset;
  assign pht_0_4_MPORT_631_data = 1'h0;
  assign pht_0_4_MPORT_631_addr = 6'h23;
  assign pht_0_4_MPORT_631_mask = 1'h1;
  assign pht_0_4_MPORT_631_en = reset;
  assign pht_0_4_MPORT_633_data = 1'h0;
  assign pht_0_4_MPORT_633_addr = 6'h24;
  assign pht_0_4_MPORT_633_mask = 1'h1;
  assign pht_0_4_MPORT_633_en = reset;
  assign pht_0_4_MPORT_635_data = 1'h0;
  assign pht_0_4_MPORT_635_addr = 6'h25;
  assign pht_0_4_MPORT_635_mask = 1'h1;
  assign pht_0_4_MPORT_635_en = reset;
  assign pht_0_4_MPORT_637_data = 1'h0;
  assign pht_0_4_MPORT_637_addr = 6'h26;
  assign pht_0_4_MPORT_637_mask = 1'h1;
  assign pht_0_4_MPORT_637_en = reset;
  assign pht_0_4_MPORT_639_data = 1'h0;
  assign pht_0_4_MPORT_639_addr = 6'h27;
  assign pht_0_4_MPORT_639_mask = 1'h1;
  assign pht_0_4_MPORT_639_en = reset;
  assign pht_0_4_MPORT_641_data = 1'h0;
  assign pht_0_4_MPORT_641_addr = 6'h28;
  assign pht_0_4_MPORT_641_mask = 1'h1;
  assign pht_0_4_MPORT_641_en = reset;
  assign pht_0_4_MPORT_643_data = 1'h0;
  assign pht_0_4_MPORT_643_addr = 6'h29;
  assign pht_0_4_MPORT_643_mask = 1'h1;
  assign pht_0_4_MPORT_643_en = reset;
  assign pht_0_4_MPORT_645_data = 1'h0;
  assign pht_0_4_MPORT_645_addr = 6'h2a;
  assign pht_0_4_MPORT_645_mask = 1'h1;
  assign pht_0_4_MPORT_645_en = reset;
  assign pht_0_4_MPORT_647_data = 1'h0;
  assign pht_0_4_MPORT_647_addr = 6'h2b;
  assign pht_0_4_MPORT_647_mask = 1'h1;
  assign pht_0_4_MPORT_647_en = reset;
  assign pht_0_4_MPORT_649_data = 1'h0;
  assign pht_0_4_MPORT_649_addr = 6'h2c;
  assign pht_0_4_MPORT_649_mask = 1'h1;
  assign pht_0_4_MPORT_649_en = reset;
  assign pht_0_4_MPORT_651_data = 1'h0;
  assign pht_0_4_MPORT_651_addr = 6'h2d;
  assign pht_0_4_MPORT_651_mask = 1'h1;
  assign pht_0_4_MPORT_651_en = reset;
  assign pht_0_4_MPORT_653_data = 1'h0;
  assign pht_0_4_MPORT_653_addr = 6'h2e;
  assign pht_0_4_MPORT_653_mask = 1'h1;
  assign pht_0_4_MPORT_653_en = reset;
  assign pht_0_4_MPORT_655_data = 1'h0;
  assign pht_0_4_MPORT_655_addr = 6'h2f;
  assign pht_0_4_MPORT_655_mask = 1'h1;
  assign pht_0_4_MPORT_655_en = reset;
  assign pht_0_4_MPORT_657_data = 1'h0;
  assign pht_0_4_MPORT_657_addr = 6'h30;
  assign pht_0_4_MPORT_657_mask = 1'h1;
  assign pht_0_4_MPORT_657_en = reset;
  assign pht_0_4_MPORT_659_data = 1'h0;
  assign pht_0_4_MPORT_659_addr = 6'h31;
  assign pht_0_4_MPORT_659_mask = 1'h1;
  assign pht_0_4_MPORT_659_en = reset;
  assign pht_0_4_MPORT_661_data = 1'h0;
  assign pht_0_4_MPORT_661_addr = 6'h32;
  assign pht_0_4_MPORT_661_mask = 1'h1;
  assign pht_0_4_MPORT_661_en = reset;
  assign pht_0_4_MPORT_663_data = 1'h0;
  assign pht_0_4_MPORT_663_addr = 6'h33;
  assign pht_0_4_MPORT_663_mask = 1'h1;
  assign pht_0_4_MPORT_663_en = reset;
  assign pht_0_4_MPORT_665_data = 1'h0;
  assign pht_0_4_MPORT_665_addr = 6'h34;
  assign pht_0_4_MPORT_665_mask = 1'h1;
  assign pht_0_4_MPORT_665_en = reset;
  assign pht_0_4_MPORT_667_data = 1'h0;
  assign pht_0_4_MPORT_667_addr = 6'h35;
  assign pht_0_4_MPORT_667_mask = 1'h1;
  assign pht_0_4_MPORT_667_en = reset;
  assign pht_0_4_MPORT_669_data = 1'h0;
  assign pht_0_4_MPORT_669_addr = 6'h36;
  assign pht_0_4_MPORT_669_mask = 1'h1;
  assign pht_0_4_MPORT_669_en = reset;
  assign pht_0_4_MPORT_671_data = 1'h0;
  assign pht_0_4_MPORT_671_addr = 6'h37;
  assign pht_0_4_MPORT_671_mask = 1'h1;
  assign pht_0_4_MPORT_671_en = reset;
  assign pht_0_4_MPORT_673_data = 1'h0;
  assign pht_0_4_MPORT_673_addr = 6'h38;
  assign pht_0_4_MPORT_673_mask = 1'h1;
  assign pht_0_4_MPORT_673_en = reset;
  assign pht_0_4_MPORT_675_data = 1'h0;
  assign pht_0_4_MPORT_675_addr = 6'h39;
  assign pht_0_4_MPORT_675_mask = 1'h1;
  assign pht_0_4_MPORT_675_en = reset;
  assign pht_0_4_MPORT_677_data = 1'h0;
  assign pht_0_4_MPORT_677_addr = 6'h3a;
  assign pht_0_4_MPORT_677_mask = 1'h1;
  assign pht_0_4_MPORT_677_en = reset;
  assign pht_0_4_MPORT_679_data = 1'h0;
  assign pht_0_4_MPORT_679_addr = 6'h3b;
  assign pht_0_4_MPORT_679_mask = 1'h1;
  assign pht_0_4_MPORT_679_en = reset;
  assign pht_0_4_MPORT_681_data = 1'h0;
  assign pht_0_4_MPORT_681_addr = 6'h3c;
  assign pht_0_4_MPORT_681_mask = 1'h1;
  assign pht_0_4_MPORT_681_en = reset;
  assign pht_0_4_MPORT_683_data = 1'h0;
  assign pht_0_4_MPORT_683_addr = 6'h3d;
  assign pht_0_4_MPORT_683_mask = 1'h1;
  assign pht_0_4_MPORT_683_en = reset;
  assign pht_0_4_MPORT_685_data = 1'h0;
  assign pht_0_4_MPORT_685_addr = 6'h3e;
  assign pht_0_4_MPORT_685_mask = 1'h1;
  assign pht_0_4_MPORT_685_en = reset;
  assign pht_0_4_MPORT_687_data = 1'h0;
  assign pht_0_4_MPORT_687_addr = 6'h3f;
  assign pht_0_4_MPORT_687_mask = 1'h1;
  assign pht_0_4_MPORT_687_en = reset;
//   assign pht_0_5_MPORT_27_en = pht_0_5_MPORT_27_en_pipe_0;
  assign pht_0_5_MPORT_27_addr = pht_0_5_MPORT_27_addr_pipe_0;
  assign pht_0_5_MPORT_27_data = pht_0_5[pht_0_5_MPORT_27_addr]; // @[PatternHistoryTable.scala 26:28]
  assign pht_0_5_MPORT_43_data = pht_wdata_w[0];
  assign pht_0_5_MPORT_43_addr = REG_47;
  assign pht_0_5_MPORT_43_mask = 1'h1;
  assign pht_0_5_MPORT_43_en = REG_29 & REG_45;
  assign pht_0_5_MPORT_689_data = 1'h0;
  assign pht_0_5_MPORT_689_addr = 6'h0;
  assign pht_0_5_MPORT_689_mask = 1'h1;
  assign pht_0_5_MPORT_689_en = reset;
  assign pht_0_5_MPORT_691_data = 1'h0;
  assign pht_0_5_MPORT_691_addr = 6'h1;
  assign pht_0_5_MPORT_691_mask = 1'h1;
  assign pht_0_5_MPORT_691_en = reset;
  assign pht_0_5_MPORT_693_data = 1'h0;
  assign pht_0_5_MPORT_693_addr = 6'h2;
  assign pht_0_5_MPORT_693_mask = 1'h1;
  assign pht_0_5_MPORT_693_en = reset;
  assign pht_0_5_MPORT_695_data = 1'h0;
  assign pht_0_5_MPORT_695_addr = 6'h3;
  assign pht_0_5_MPORT_695_mask = 1'h1;
  assign pht_0_5_MPORT_695_en = reset;
  assign pht_0_5_MPORT_697_data = 1'h0;
  assign pht_0_5_MPORT_697_addr = 6'h4;
  assign pht_0_5_MPORT_697_mask = 1'h1;
  assign pht_0_5_MPORT_697_en = reset;
  assign pht_0_5_MPORT_699_data = 1'h0;
  assign pht_0_5_MPORT_699_addr = 6'h5;
  assign pht_0_5_MPORT_699_mask = 1'h1;
  assign pht_0_5_MPORT_699_en = reset;
  assign pht_0_5_MPORT_701_data = 1'h0;
  assign pht_0_5_MPORT_701_addr = 6'h6;
  assign pht_0_5_MPORT_701_mask = 1'h1;
  assign pht_0_5_MPORT_701_en = reset;
  assign pht_0_5_MPORT_703_data = 1'h0;
  assign pht_0_5_MPORT_703_addr = 6'h7;
  assign pht_0_5_MPORT_703_mask = 1'h1;
  assign pht_0_5_MPORT_703_en = reset;
  assign pht_0_5_MPORT_705_data = 1'h0;
  assign pht_0_5_MPORT_705_addr = 6'h8;
  assign pht_0_5_MPORT_705_mask = 1'h1;
  assign pht_0_5_MPORT_705_en = reset;
  assign pht_0_5_MPORT_707_data = 1'h0;
  assign pht_0_5_MPORT_707_addr = 6'h9;
  assign pht_0_5_MPORT_707_mask = 1'h1;
  assign pht_0_5_MPORT_707_en = reset;
  assign pht_0_5_MPORT_709_data = 1'h0;
  assign pht_0_5_MPORT_709_addr = 6'ha;
  assign pht_0_5_MPORT_709_mask = 1'h1;
  assign pht_0_5_MPORT_709_en = reset;
  assign pht_0_5_MPORT_711_data = 1'h0;
  assign pht_0_5_MPORT_711_addr = 6'hb;
  assign pht_0_5_MPORT_711_mask = 1'h1;
  assign pht_0_5_MPORT_711_en = reset;
  assign pht_0_5_MPORT_713_data = 1'h0;
  assign pht_0_5_MPORT_713_addr = 6'hc;
  assign pht_0_5_MPORT_713_mask = 1'h1;
  assign pht_0_5_MPORT_713_en = reset;
  assign pht_0_5_MPORT_715_data = 1'h0;
  assign pht_0_5_MPORT_715_addr = 6'hd;
  assign pht_0_5_MPORT_715_mask = 1'h1;
  assign pht_0_5_MPORT_715_en = reset;
  assign pht_0_5_MPORT_717_data = 1'h0;
  assign pht_0_5_MPORT_717_addr = 6'he;
  assign pht_0_5_MPORT_717_mask = 1'h1;
  assign pht_0_5_MPORT_717_en = reset;
  assign pht_0_5_MPORT_719_data = 1'h0;
  assign pht_0_5_MPORT_719_addr = 6'hf;
  assign pht_0_5_MPORT_719_mask = 1'h1;
  assign pht_0_5_MPORT_719_en = reset;
  assign pht_0_5_MPORT_721_data = 1'h0;
  assign pht_0_5_MPORT_721_addr = 6'h10;
  assign pht_0_5_MPORT_721_mask = 1'h1;
  assign pht_0_5_MPORT_721_en = reset;
  assign pht_0_5_MPORT_723_data = 1'h0;
  assign pht_0_5_MPORT_723_addr = 6'h11;
  assign pht_0_5_MPORT_723_mask = 1'h1;
  assign pht_0_5_MPORT_723_en = reset;
  assign pht_0_5_MPORT_725_data = 1'h0;
  assign pht_0_5_MPORT_725_addr = 6'h12;
  assign pht_0_5_MPORT_725_mask = 1'h1;
  assign pht_0_5_MPORT_725_en = reset;
  assign pht_0_5_MPORT_727_data = 1'h0;
  assign pht_0_5_MPORT_727_addr = 6'h13;
  assign pht_0_5_MPORT_727_mask = 1'h1;
  assign pht_0_5_MPORT_727_en = reset;
  assign pht_0_5_MPORT_729_data = 1'h0;
  assign pht_0_5_MPORT_729_addr = 6'h14;
  assign pht_0_5_MPORT_729_mask = 1'h1;
  assign pht_0_5_MPORT_729_en = reset;
  assign pht_0_5_MPORT_731_data = 1'h0;
  assign pht_0_5_MPORT_731_addr = 6'h15;
  assign pht_0_5_MPORT_731_mask = 1'h1;
  assign pht_0_5_MPORT_731_en = reset;
  assign pht_0_5_MPORT_733_data = 1'h0;
  assign pht_0_5_MPORT_733_addr = 6'h16;
  assign pht_0_5_MPORT_733_mask = 1'h1;
  assign pht_0_5_MPORT_733_en = reset;
  assign pht_0_5_MPORT_735_data = 1'h0;
  assign pht_0_5_MPORT_735_addr = 6'h17;
  assign pht_0_5_MPORT_735_mask = 1'h1;
  assign pht_0_5_MPORT_735_en = reset;
  assign pht_0_5_MPORT_737_data = 1'h0;
  assign pht_0_5_MPORT_737_addr = 6'h18;
  assign pht_0_5_MPORT_737_mask = 1'h1;
  assign pht_0_5_MPORT_737_en = reset;
  assign pht_0_5_MPORT_739_data = 1'h0;
  assign pht_0_5_MPORT_739_addr = 6'h19;
  assign pht_0_5_MPORT_739_mask = 1'h1;
  assign pht_0_5_MPORT_739_en = reset;
  assign pht_0_5_MPORT_741_data = 1'h0;
  assign pht_0_5_MPORT_741_addr = 6'h1a;
  assign pht_0_5_MPORT_741_mask = 1'h1;
  assign pht_0_5_MPORT_741_en = reset;
  assign pht_0_5_MPORT_743_data = 1'h0;
  assign pht_0_5_MPORT_743_addr = 6'h1b;
  assign pht_0_5_MPORT_743_mask = 1'h1;
  assign pht_0_5_MPORT_743_en = reset;
  assign pht_0_5_MPORT_745_data = 1'h0;
  assign pht_0_5_MPORT_745_addr = 6'h1c;
  assign pht_0_5_MPORT_745_mask = 1'h1;
  assign pht_0_5_MPORT_745_en = reset;
  assign pht_0_5_MPORT_747_data = 1'h0;
  assign pht_0_5_MPORT_747_addr = 6'h1d;
  assign pht_0_5_MPORT_747_mask = 1'h1;
  assign pht_0_5_MPORT_747_en = reset;
  assign pht_0_5_MPORT_749_data = 1'h0;
  assign pht_0_5_MPORT_749_addr = 6'h1e;
  assign pht_0_5_MPORT_749_mask = 1'h1;
  assign pht_0_5_MPORT_749_en = reset;
  assign pht_0_5_MPORT_751_data = 1'h0;
  assign pht_0_5_MPORT_751_addr = 6'h1f;
  assign pht_0_5_MPORT_751_mask = 1'h1;
  assign pht_0_5_MPORT_751_en = reset;
  assign pht_0_5_MPORT_753_data = 1'h0;
  assign pht_0_5_MPORT_753_addr = 6'h20;
  assign pht_0_5_MPORT_753_mask = 1'h1;
  assign pht_0_5_MPORT_753_en = reset;
  assign pht_0_5_MPORT_755_data = 1'h0;
  assign pht_0_5_MPORT_755_addr = 6'h21;
  assign pht_0_5_MPORT_755_mask = 1'h1;
  assign pht_0_5_MPORT_755_en = reset;
  assign pht_0_5_MPORT_757_data = 1'h0;
  assign pht_0_5_MPORT_757_addr = 6'h22;
  assign pht_0_5_MPORT_757_mask = 1'h1;
  assign pht_0_5_MPORT_757_en = reset;
  assign pht_0_5_MPORT_759_data = 1'h0;
  assign pht_0_5_MPORT_759_addr = 6'h23;
  assign pht_0_5_MPORT_759_mask = 1'h1;
  assign pht_0_5_MPORT_759_en = reset;
  assign pht_0_5_MPORT_761_data = 1'h0;
  assign pht_0_5_MPORT_761_addr = 6'h24;
  assign pht_0_5_MPORT_761_mask = 1'h1;
  assign pht_0_5_MPORT_761_en = reset;
  assign pht_0_5_MPORT_763_data = 1'h0;
  assign pht_0_5_MPORT_763_addr = 6'h25;
  assign pht_0_5_MPORT_763_mask = 1'h1;
  assign pht_0_5_MPORT_763_en = reset;
  assign pht_0_5_MPORT_765_data = 1'h0;
  assign pht_0_5_MPORT_765_addr = 6'h26;
  assign pht_0_5_MPORT_765_mask = 1'h1;
  assign pht_0_5_MPORT_765_en = reset;
  assign pht_0_5_MPORT_767_data = 1'h0;
  assign pht_0_5_MPORT_767_addr = 6'h27;
  assign pht_0_5_MPORT_767_mask = 1'h1;
  assign pht_0_5_MPORT_767_en = reset;
  assign pht_0_5_MPORT_769_data = 1'h0;
  assign pht_0_5_MPORT_769_addr = 6'h28;
  assign pht_0_5_MPORT_769_mask = 1'h1;
  assign pht_0_5_MPORT_769_en = reset;
  assign pht_0_5_MPORT_771_data = 1'h0;
  assign pht_0_5_MPORT_771_addr = 6'h29;
  assign pht_0_5_MPORT_771_mask = 1'h1;
  assign pht_0_5_MPORT_771_en = reset;
  assign pht_0_5_MPORT_773_data = 1'h0;
  assign pht_0_5_MPORT_773_addr = 6'h2a;
  assign pht_0_5_MPORT_773_mask = 1'h1;
  assign pht_0_5_MPORT_773_en = reset;
  assign pht_0_5_MPORT_775_data = 1'h0;
  assign pht_0_5_MPORT_775_addr = 6'h2b;
  assign pht_0_5_MPORT_775_mask = 1'h1;
  assign pht_0_5_MPORT_775_en = reset;
  assign pht_0_5_MPORT_777_data = 1'h0;
  assign pht_0_5_MPORT_777_addr = 6'h2c;
  assign pht_0_5_MPORT_777_mask = 1'h1;
  assign pht_0_5_MPORT_777_en = reset;
  assign pht_0_5_MPORT_779_data = 1'h0;
  assign pht_0_5_MPORT_779_addr = 6'h2d;
  assign pht_0_5_MPORT_779_mask = 1'h1;
  assign pht_0_5_MPORT_779_en = reset;
  assign pht_0_5_MPORT_781_data = 1'h0;
  assign pht_0_5_MPORT_781_addr = 6'h2e;
  assign pht_0_5_MPORT_781_mask = 1'h1;
  assign pht_0_5_MPORT_781_en = reset;
  assign pht_0_5_MPORT_783_data = 1'h0;
  assign pht_0_5_MPORT_783_addr = 6'h2f;
  assign pht_0_5_MPORT_783_mask = 1'h1;
  assign pht_0_5_MPORT_783_en = reset;
  assign pht_0_5_MPORT_785_data = 1'h0;
  assign pht_0_5_MPORT_785_addr = 6'h30;
  assign pht_0_5_MPORT_785_mask = 1'h1;
  assign pht_0_5_MPORT_785_en = reset;
  assign pht_0_5_MPORT_787_data = 1'h0;
  assign pht_0_5_MPORT_787_addr = 6'h31;
  assign pht_0_5_MPORT_787_mask = 1'h1;
  assign pht_0_5_MPORT_787_en = reset;
  assign pht_0_5_MPORT_789_data = 1'h0;
  assign pht_0_5_MPORT_789_addr = 6'h32;
  assign pht_0_5_MPORT_789_mask = 1'h1;
  assign pht_0_5_MPORT_789_en = reset;
  assign pht_0_5_MPORT_791_data = 1'h0;
  assign pht_0_5_MPORT_791_addr = 6'h33;
  assign pht_0_5_MPORT_791_mask = 1'h1;
  assign pht_0_5_MPORT_791_en = reset;
  assign pht_0_5_MPORT_793_data = 1'h0;
  assign pht_0_5_MPORT_793_addr = 6'h34;
  assign pht_0_5_MPORT_793_mask = 1'h1;
  assign pht_0_5_MPORT_793_en = reset;
  assign pht_0_5_MPORT_795_data = 1'h0;
  assign pht_0_5_MPORT_795_addr = 6'h35;
  assign pht_0_5_MPORT_795_mask = 1'h1;
  assign pht_0_5_MPORT_795_en = reset;
  assign pht_0_5_MPORT_797_data = 1'h0;
  assign pht_0_5_MPORT_797_addr = 6'h36;
  assign pht_0_5_MPORT_797_mask = 1'h1;
  assign pht_0_5_MPORT_797_en = reset;
  assign pht_0_5_MPORT_799_data = 1'h0;
  assign pht_0_5_MPORT_799_addr = 6'h37;
  assign pht_0_5_MPORT_799_mask = 1'h1;
  assign pht_0_5_MPORT_799_en = reset;
  assign pht_0_5_MPORT_801_data = 1'h0;
  assign pht_0_5_MPORT_801_addr = 6'h38;
  assign pht_0_5_MPORT_801_mask = 1'h1;
  assign pht_0_5_MPORT_801_en = reset;
  assign pht_0_5_MPORT_803_data = 1'h0;
  assign pht_0_5_MPORT_803_addr = 6'h39;
  assign pht_0_5_MPORT_803_mask = 1'h1;
  assign pht_0_5_MPORT_803_en = reset;
  assign pht_0_5_MPORT_805_data = 1'h0;
  assign pht_0_5_MPORT_805_addr = 6'h3a;
  assign pht_0_5_MPORT_805_mask = 1'h1;
  assign pht_0_5_MPORT_805_en = reset;
  assign pht_0_5_MPORT_807_data = 1'h0;
  assign pht_0_5_MPORT_807_addr = 6'h3b;
  assign pht_0_5_MPORT_807_mask = 1'h1;
  assign pht_0_5_MPORT_807_en = reset;
  assign pht_0_5_MPORT_809_data = 1'h0;
  assign pht_0_5_MPORT_809_addr = 6'h3c;
  assign pht_0_5_MPORT_809_mask = 1'h1;
  assign pht_0_5_MPORT_809_en = reset;
  assign pht_0_5_MPORT_811_data = 1'h0;
  assign pht_0_5_MPORT_811_addr = 6'h3d;
  assign pht_0_5_MPORT_811_mask = 1'h1;
  assign pht_0_5_MPORT_811_en = reset;
  assign pht_0_5_MPORT_813_data = 1'h0;
  assign pht_0_5_MPORT_813_addr = 6'h3e;
  assign pht_0_5_MPORT_813_mask = 1'h1;
  assign pht_0_5_MPORT_813_en = reset;
  assign pht_0_5_MPORT_815_data = 1'h0;
  assign pht_0_5_MPORT_815_addr = 6'h3f;
  assign pht_0_5_MPORT_815_mask = 1'h1;
  assign pht_0_5_MPORT_815_en = reset;
//   assign pht_0_6_MPORT_29_en = pht_0_6_MPORT_29_en_pipe_0;
  assign pht_0_6_MPORT_29_addr = pht_0_6_MPORT_29_addr_pipe_0;
  assign pht_0_6_MPORT_29_data = pht_0_6[pht_0_6_MPORT_29_addr]; // @[PatternHistoryTable.scala 26:28]
  assign pht_0_6_MPORT_45_data = pht_wdata_w[0];
  assign pht_0_6_MPORT_45_addr = REG_50;
  assign pht_0_6_MPORT_45_mask = 1'h1;
  assign pht_0_6_MPORT_45_en = REG_29 & REG_48;
  assign pht_0_6_MPORT_817_data = 1'h0;
  assign pht_0_6_MPORT_817_addr = 6'h0;
  assign pht_0_6_MPORT_817_mask = 1'h1;
  assign pht_0_6_MPORT_817_en = reset;
  assign pht_0_6_MPORT_819_data = 1'h0;
  assign pht_0_6_MPORT_819_addr = 6'h1;
  assign pht_0_6_MPORT_819_mask = 1'h1;
  assign pht_0_6_MPORT_819_en = reset;
  assign pht_0_6_MPORT_821_data = 1'h0;
  assign pht_0_6_MPORT_821_addr = 6'h2;
  assign pht_0_6_MPORT_821_mask = 1'h1;
  assign pht_0_6_MPORT_821_en = reset;
  assign pht_0_6_MPORT_823_data = 1'h0;
  assign pht_0_6_MPORT_823_addr = 6'h3;
  assign pht_0_6_MPORT_823_mask = 1'h1;
  assign pht_0_6_MPORT_823_en = reset;
  assign pht_0_6_MPORT_825_data = 1'h0;
  assign pht_0_6_MPORT_825_addr = 6'h4;
  assign pht_0_6_MPORT_825_mask = 1'h1;
  assign pht_0_6_MPORT_825_en = reset;
  assign pht_0_6_MPORT_827_data = 1'h0;
  assign pht_0_6_MPORT_827_addr = 6'h5;
  assign pht_0_6_MPORT_827_mask = 1'h1;
  assign pht_0_6_MPORT_827_en = reset;
  assign pht_0_6_MPORT_829_data = 1'h0;
  assign pht_0_6_MPORT_829_addr = 6'h6;
  assign pht_0_6_MPORT_829_mask = 1'h1;
  assign pht_0_6_MPORT_829_en = reset;
  assign pht_0_6_MPORT_831_data = 1'h0;
  assign pht_0_6_MPORT_831_addr = 6'h7;
  assign pht_0_6_MPORT_831_mask = 1'h1;
  assign pht_0_6_MPORT_831_en = reset;
  assign pht_0_6_MPORT_833_data = 1'h0;
  assign pht_0_6_MPORT_833_addr = 6'h8;
  assign pht_0_6_MPORT_833_mask = 1'h1;
  assign pht_0_6_MPORT_833_en = reset;
  assign pht_0_6_MPORT_835_data = 1'h0;
  assign pht_0_6_MPORT_835_addr = 6'h9;
  assign pht_0_6_MPORT_835_mask = 1'h1;
  assign pht_0_6_MPORT_835_en = reset;
  assign pht_0_6_MPORT_837_data = 1'h0;
  assign pht_0_6_MPORT_837_addr = 6'ha;
  assign pht_0_6_MPORT_837_mask = 1'h1;
  assign pht_0_6_MPORT_837_en = reset;
  assign pht_0_6_MPORT_839_data = 1'h0;
  assign pht_0_6_MPORT_839_addr = 6'hb;
  assign pht_0_6_MPORT_839_mask = 1'h1;
  assign pht_0_6_MPORT_839_en = reset;
  assign pht_0_6_MPORT_841_data = 1'h0;
  assign pht_0_6_MPORT_841_addr = 6'hc;
  assign pht_0_6_MPORT_841_mask = 1'h1;
  assign pht_0_6_MPORT_841_en = reset;
  assign pht_0_6_MPORT_843_data = 1'h0;
  assign pht_0_6_MPORT_843_addr = 6'hd;
  assign pht_0_6_MPORT_843_mask = 1'h1;
  assign pht_0_6_MPORT_843_en = reset;
  assign pht_0_6_MPORT_845_data = 1'h0;
  assign pht_0_6_MPORT_845_addr = 6'he;
  assign pht_0_6_MPORT_845_mask = 1'h1;
  assign pht_0_6_MPORT_845_en = reset;
  assign pht_0_6_MPORT_847_data = 1'h0;
  assign pht_0_6_MPORT_847_addr = 6'hf;
  assign pht_0_6_MPORT_847_mask = 1'h1;
  assign pht_0_6_MPORT_847_en = reset;
  assign pht_0_6_MPORT_849_data = 1'h0;
  assign pht_0_6_MPORT_849_addr = 6'h10;
  assign pht_0_6_MPORT_849_mask = 1'h1;
  assign pht_0_6_MPORT_849_en = reset;
  assign pht_0_6_MPORT_851_data = 1'h0;
  assign pht_0_6_MPORT_851_addr = 6'h11;
  assign pht_0_6_MPORT_851_mask = 1'h1;
  assign pht_0_6_MPORT_851_en = reset;
  assign pht_0_6_MPORT_853_data = 1'h0;
  assign pht_0_6_MPORT_853_addr = 6'h12;
  assign pht_0_6_MPORT_853_mask = 1'h1;
  assign pht_0_6_MPORT_853_en = reset;
  assign pht_0_6_MPORT_855_data = 1'h0;
  assign pht_0_6_MPORT_855_addr = 6'h13;
  assign pht_0_6_MPORT_855_mask = 1'h1;
  assign pht_0_6_MPORT_855_en = reset;
  assign pht_0_6_MPORT_857_data = 1'h0;
  assign pht_0_6_MPORT_857_addr = 6'h14;
  assign pht_0_6_MPORT_857_mask = 1'h1;
  assign pht_0_6_MPORT_857_en = reset;
  assign pht_0_6_MPORT_859_data = 1'h0;
  assign pht_0_6_MPORT_859_addr = 6'h15;
  assign pht_0_6_MPORT_859_mask = 1'h1;
  assign pht_0_6_MPORT_859_en = reset;
  assign pht_0_6_MPORT_861_data = 1'h0;
  assign pht_0_6_MPORT_861_addr = 6'h16;
  assign pht_0_6_MPORT_861_mask = 1'h1;
  assign pht_0_6_MPORT_861_en = reset;
  assign pht_0_6_MPORT_863_data = 1'h0;
  assign pht_0_6_MPORT_863_addr = 6'h17;
  assign pht_0_6_MPORT_863_mask = 1'h1;
  assign pht_0_6_MPORT_863_en = reset;
  assign pht_0_6_MPORT_865_data = 1'h0;
  assign pht_0_6_MPORT_865_addr = 6'h18;
  assign pht_0_6_MPORT_865_mask = 1'h1;
  assign pht_0_6_MPORT_865_en = reset;
  assign pht_0_6_MPORT_867_data = 1'h0;
  assign pht_0_6_MPORT_867_addr = 6'h19;
  assign pht_0_6_MPORT_867_mask = 1'h1;
  assign pht_0_6_MPORT_867_en = reset;
  assign pht_0_6_MPORT_869_data = 1'h0;
  assign pht_0_6_MPORT_869_addr = 6'h1a;
  assign pht_0_6_MPORT_869_mask = 1'h1;
  assign pht_0_6_MPORT_869_en = reset;
  assign pht_0_6_MPORT_871_data = 1'h0;
  assign pht_0_6_MPORT_871_addr = 6'h1b;
  assign pht_0_6_MPORT_871_mask = 1'h1;
  assign pht_0_6_MPORT_871_en = reset;
  assign pht_0_6_MPORT_873_data = 1'h0;
  assign pht_0_6_MPORT_873_addr = 6'h1c;
  assign pht_0_6_MPORT_873_mask = 1'h1;
  assign pht_0_6_MPORT_873_en = reset;
  assign pht_0_6_MPORT_875_data = 1'h0;
  assign pht_0_6_MPORT_875_addr = 6'h1d;
  assign pht_0_6_MPORT_875_mask = 1'h1;
  assign pht_0_6_MPORT_875_en = reset;
  assign pht_0_6_MPORT_877_data = 1'h0;
  assign pht_0_6_MPORT_877_addr = 6'h1e;
  assign pht_0_6_MPORT_877_mask = 1'h1;
  assign pht_0_6_MPORT_877_en = reset;
  assign pht_0_6_MPORT_879_data = 1'h0;
  assign pht_0_6_MPORT_879_addr = 6'h1f;
  assign pht_0_6_MPORT_879_mask = 1'h1;
  assign pht_0_6_MPORT_879_en = reset;
  assign pht_0_6_MPORT_881_data = 1'h0;
  assign pht_0_6_MPORT_881_addr = 6'h20;
  assign pht_0_6_MPORT_881_mask = 1'h1;
  assign pht_0_6_MPORT_881_en = reset;
  assign pht_0_6_MPORT_883_data = 1'h0;
  assign pht_0_6_MPORT_883_addr = 6'h21;
  assign pht_0_6_MPORT_883_mask = 1'h1;
  assign pht_0_6_MPORT_883_en = reset;
  assign pht_0_6_MPORT_885_data = 1'h0;
  assign pht_0_6_MPORT_885_addr = 6'h22;
  assign pht_0_6_MPORT_885_mask = 1'h1;
  assign pht_0_6_MPORT_885_en = reset;
  assign pht_0_6_MPORT_887_data = 1'h0;
  assign pht_0_6_MPORT_887_addr = 6'h23;
  assign pht_0_6_MPORT_887_mask = 1'h1;
  assign pht_0_6_MPORT_887_en = reset;
  assign pht_0_6_MPORT_889_data = 1'h0;
  assign pht_0_6_MPORT_889_addr = 6'h24;
  assign pht_0_6_MPORT_889_mask = 1'h1;
  assign pht_0_6_MPORT_889_en = reset;
  assign pht_0_6_MPORT_891_data = 1'h0;
  assign pht_0_6_MPORT_891_addr = 6'h25;
  assign pht_0_6_MPORT_891_mask = 1'h1;
  assign pht_0_6_MPORT_891_en = reset;
  assign pht_0_6_MPORT_893_data = 1'h0;
  assign pht_0_6_MPORT_893_addr = 6'h26;
  assign pht_0_6_MPORT_893_mask = 1'h1;
  assign pht_0_6_MPORT_893_en = reset;
  assign pht_0_6_MPORT_895_data = 1'h0;
  assign pht_0_6_MPORT_895_addr = 6'h27;
  assign pht_0_6_MPORT_895_mask = 1'h1;
  assign pht_0_6_MPORT_895_en = reset;
  assign pht_0_6_MPORT_897_data = 1'h0;
  assign pht_0_6_MPORT_897_addr = 6'h28;
  assign pht_0_6_MPORT_897_mask = 1'h1;
  assign pht_0_6_MPORT_897_en = reset;
  assign pht_0_6_MPORT_899_data = 1'h0;
  assign pht_0_6_MPORT_899_addr = 6'h29;
  assign pht_0_6_MPORT_899_mask = 1'h1;
  assign pht_0_6_MPORT_899_en = reset;
  assign pht_0_6_MPORT_901_data = 1'h0;
  assign pht_0_6_MPORT_901_addr = 6'h2a;
  assign pht_0_6_MPORT_901_mask = 1'h1;
  assign pht_0_6_MPORT_901_en = reset;
  assign pht_0_6_MPORT_903_data = 1'h0;
  assign pht_0_6_MPORT_903_addr = 6'h2b;
  assign pht_0_6_MPORT_903_mask = 1'h1;
  assign pht_0_6_MPORT_903_en = reset;
  assign pht_0_6_MPORT_905_data = 1'h0;
  assign pht_0_6_MPORT_905_addr = 6'h2c;
  assign pht_0_6_MPORT_905_mask = 1'h1;
  assign pht_0_6_MPORT_905_en = reset;
  assign pht_0_6_MPORT_907_data = 1'h0;
  assign pht_0_6_MPORT_907_addr = 6'h2d;
  assign pht_0_6_MPORT_907_mask = 1'h1;
  assign pht_0_6_MPORT_907_en = reset;
  assign pht_0_6_MPORT_909_data = 1'h0;
  assign pht_0_6_MPORT_909_addr = 6'h2e;
  assign pht_0_6_MPORT_909_mask = 1'h1;
  assign pht_0_6_MPORT_909_en = reset;
  assign pht_0_6_MPORT_911_data = 1'h0;
  assign pht_0_6_MPORT_911_addr = 6'h2f;
  assign pht_0_6_MPORT_911_mask = 1'h1;
  assign pht_0_6_MPORT_911_en = reset;
  assign pht_0_6_MPORT_913_data = 1'h0;
  assign pht_0_6_MPORT_913_addr = 6'h30;
  assign pht_0_6_MPORT_913_mask = 1'h1;
  assign pht_0_6_MPORT_913_en = reset;
  assign pht_0_6_MPORT_915_data = 1'h0;
  assign pht_0_6_MPORT_915_addr = 6'h31;
  assign pht_0_6_MPORT_915_mask = 1'h1;
  assign pht_0_6_MPORT_915_en = reset;
  assign pht_0_6_MPORT_917_data = 1'h0;
  assign pht_0_6_MPORT_917_addr = 6'h32;
  assign pht_0_6_MPORT_917_mask = 1'h1;
  assign pht_0_6_MPORT_917_en = reset;
  assign pht_0_6_MPORT_919_data = 1'h0;
  assign pht_0_6_MPORT_919_addr = 6'h33;
  assign pht_0_6_MPORT_919_mask = 1'h1;
  assign pht_0_6_MPORT_919_en = reset;
  assign pht_0_6_MPORT_921_data = 1'h0;
  assign pht_0_6_MPORT_921_addr = 6'h34;
  assign pht_0_6_MPORT_921_mask = 1'h1;
  assign pht_0_6_MPORT_921_en = reset;
  assign pht_0_6_MPORT_923_data = 1'h0;
  assign pht_0_6_MPORT_923_addr = 6'h35;
  assign pht_0_6_MPORT_923_mask = 1'h1;
  assign pht_0_6_MPORT_923_en = reset;
  assign pht_0_6_MPORT_925_data = 1'h0;
  assign pht_0_6_MPORT_925_addr = 6'h36;
  assign pht_0_6_MPORT_925_mask = 1'h1;
  assign pht_0_6_MPORT_925_en = reset;
  assign pht_0_6_MPORT_927_data = 1'h0;
  assign pht_0_6_MPORT_927_addr = 6'h37;
  assign pht_0_6_MPORT_927_mask = 1'h1;
  assign pht_0_6_MPORT_927_en = reset;
  assign pht_0_6_MPORT_929_data = 1'h0;
  assign pht_0_6_MPORT_929_addr = 6'h38;
  assign pht_0_6_MPORT_929_mask = 1'h1;
  assign pht_0_6_MPORT_929_en = reset;
  assign pht_0_6_MPORT_931_data = 1'h0;
  assign pht_0_6_MPORT_931_addr = 6'h39;
  assign pht_0_6_MPORT_931_mask = 1'h1;
  assign pht_0_6_MPORT_931_en = reset;
  assign pht_0_6_MPORT_933_data = 1'h0;
  assign pht_0_6_MPORT_933_addr = 6'h3a;
  assign pht_0_6_MPORT_933_mask = 1'h1;
  assign pht_0_6_MPORT_933_en = reset;
  assign pht_0_6_MPORT_935_data = 1'h0;
  assign pht_0_6_MPORT_935_addr = 6'h3b;
  assign pht_0_6_MPORT_935_mask = 1'h1;
  assign pht_0_6_MPORT_935_en = reset;
  assign pht_0_6_MPORT_937_data = 1'h0;
  assign pht_0_6_MPORT_937_addr = 6'h3c;
  assign pht_0_6_MPORT_937_mask = 1'h1;
  assign pht_0_6_MPORT_937_en = reset;
  assign pht_0_6_MPORT_939_data = 1'h0;
  assign pht_0_6_MPORT_939_addr = 6'h3d;
  assign pht_0_6_MPORT_939_mask = 1'h1;
  assign pht_0_6_MPORT_939_en = reset;
  assign pht_0_6_MPORT_941_data = 1'h0;
  assign pht_0_6_MPORT_941_addr = 6'h3e;
  assign pht_0_6_MPORT_941_mask = 1'h1;
  assign pht_0_6_MPORT_941_en = reset;
  assign pht_0_6_MPORT_943_data = 1'h0;
  assign pht_0_6_MPORT_943_addr = 6'h3f;
  assign pht_0_6_MPORT_943_mask = 1'h1;
  assign pht_0_6_MPORT_943_en = reset;
//   assign pht_0_7_MPORT_31_en = pht_0_7_MPORT_31_en_pipe_0;
  assign pht_0_7_MPORT_31_addr = pht_0_7_MPORT_31_addr_pipe_0;
  assign pht_0_7_MPORT_31_data = pht_0_7[pht_0_7_MPORT_31_addr]; // @[PatternHistoryTable.scala 26:28]
  assign pht_0_7_MPORT_47_data = pht_wdata_w[0];
  assign pht_0_7_MPORT_47_addr = REG_53;
  assign pht_0_7_MPORT_47_mask = 1'h1;
  assign pht_0_7_MPORT_47_en = REG_29 & REG_51;
  assign pht_0_7_MPORT_945_data = 1'h0;
  assign pht_0_7_MPORT_945_addr = 6'h0;
  assign pht_0_7_MPORT_945_mask = 1'h1;
  assign pht_0_7_MPORT_945_en = reset;
  assign pht_0_7_MPORT_947_data = 1'h0;
  assign pht_0_7_MPORT_947_addr = 6'h1;
  assign pht_0_7_MPORT_947_mask = 1'h1;
  assign pht_0_7_MPORT_947_en = reset;
  assign pht_0_7_MPORT_949_data = 1'h0;
  assign pht_0_7_MPORT_949_addr = 6'h2;
  assign pht_0_7_MPORT_949_mask = 1'h1;
  assign pht_0_7_MPORT_949_en = reset;
  assign pht_0_7_MPORT_951_data = 1'h0;
  assign pht_0_7_MPORT_951_addr = 6'h3;
  assign pht_0_7_MPORT_951_mask = 1'h1;
  assign pht_0_7_MPORT_951_en = reset;
  assign pht_0_7_MPORT_953_data = 1'h0;
  assign pht_0_7_MPORT_953_addr = 6'h4;
  assign pht_0_7_MPORT_953_mask = 1'h1;
  assign pht_0_7_MPORT_953_en = reset;
  assign pht_0_7_MPORT_955_data = 1'h0;
  assign pht_0_7_MPORT_955_addr = 6'h5;
  assign pht_0_7_MPORT_955_mask = 1'h1;
  assign pht_0_7_MPORT_955_en = reset;
  assign pht_0_7_MPORT_957_data = 1'h0;
  assign pht_0_7_MPORT_957_addr = 6'h6;
  assign pht_0_7_MPORT_957_mask = 1'h1;
  assign pht_0_7_MPORT_957_en = reset;
  assign pht_0_7_MPORT_959_data = 1'h0;
  assign pht_0_7_MPORT_959_addr = 6'h7;
  assign pht_0_7_MPORT_959_mask = 1'h1;
  assign pht_0_7_MPORT_959_en = reset;
  assign pht_0_7_MPORT_961_data = 1'h0;
  assign pht_0_7_MPORT_961_addr = 6'h8;
  assign pht_0_7_MPORT_961_mask = 1'h1;
  assign pht_0_7_MPORT_961_en = reset;
  assign pht_0_7_MPORT_963_data = 1'h0;
  assign pht_0_7_MPORT_963_addr = 6'h9;
  assign pht_0_7_MPORT_963_mask = 1'h1;
  assign pht_0_7_MPORT_963_en = reset;
  assign pht_0_7_MPORT_965_data = 1'h0;
  assign pht_0_7_MPORT_965_addr = 6'ha;
  assign pht_0_7_MPORT_965_mask = 1'h1;
  assign pht_0_7_MPORT_965_en = reset;
  assign pht_0_7_MPORT_967_data = 1'h0;
  assign pht_0_7_MPORT_967_addr = 6'hb;
  assign pht_0_7_MPORT_967_mask = 1'h1;
  assign pht_0_7_MPORT_967_en = reset;
  assign pht_0_7_MPORT_969_data = 1'h0;
  assign pht_0_7_MPORT_969_addr = 6'hc;
  assign pht_0_7_MPORT_969_mask = 1'h1;
  assign pht_0_7_MPORT_969_en = reset;
  assign pht_0_7_MPORT_971_data = 1'h0;
  assign pht_0_7_MPORT_971_addr = 6'hd;
  assign pht_0_7_MPORT_971_mask = 1'h1;
  assign pht_0_7_MPORT_971_en = reset;
  assign pht_0_7_MPORT_973_data = 1'h0;
  assign pht_0_7_MPORT_973_addr = 6'he;
  assign pht_0_7_MPORT_973_mask = 1'h1;
  assign pht_0_7_MPORT_973_en = reset;
  assign pht_0_7_MPORT_975_data = 1'h0;
  assign pht_0_7_MPORT_975_addr = 6'hf;
  assign pht_0_7_MPORT_975_mask = 1'h1;
  assign pht_0_7_MPORT_975_en = reset;
  assign pht_0_7_MPORT_977_data = 1'h0;
  assign pht_0_7_MPORT_977_addr = 6'h10;
  assign pht_0_7_MPORT_977_mask = 1'h1;
  assign pht_0_7_MPORT_977_en = reset;
  assign pht_0_7_MPORT_979_data = 1'h0;
  assign pht_0_7_MPORT_979_addr = 6'h11;
  assign pht_0_7_MPORT_979_mask = 1'h1;
  assign pht_0_7_MPORT_979_en = reset;
  assign pht_0_7_MPORT_981_data = 1'h0;
  assign pht_0_7_MPORT_981_addr = 6'h12;
  assign pht_0_7_MPORT_981_mask = 1'h1;
  assign pht_0_7_MPORT_981_en = reset;
  assign pht_0_7_MPORT_983_data = 1'h0;
  assign pht_0_7_MPORT_983_addr = 6'h13;
  assign pht_0_7_MPORT_983_mask = 1'h1;
  assign pht_0_7_MPORT_983_en = reset;
  assign pht_0_7_MPORT_985_data = 1'h0;
  assign pht_0_7_MPORT_985_addr = 6'h14;
  assign pht_0_7_MPORT_985_mask = 1'h1;
  assign pht_0_7_MPORT_985_en = reset;
  assign pht_0_7_MPORT_987_data = 1'h0;
  assign pht_0_7_MPORT_987_addr = 6'h15;
  assign pht_0_7_MPORT_987_mask = 1'h1;
  assign pht_0_7_MPORT_987_en = reset;
  assign pht_0_7_MPORT_989_data = 1'h0;
  assign pht_0_7_MPORT_989_addr = 6'h16;
  assign pht_0_7_MPORT_989_mask = 1'h1;
  assign pht_0_7_MPORT_989_en = reset;
  assign pht_0_7_MPORT_991_data = 1'h0;
  assign pht_0_7_MPORT_991_addr = 6'h17;
  assign pht_0_7_MPORT_991_mask = 1'h1;
  assign pht_0_7_MPORT_991_en = reset;
  assign pht_0_7_MPORT_993_data = 1'h0;
  assign pht_0_7_MPORT_993_addr = 6'h18;
  assign pht_0_7_MPORT_993_mask = 1'h1;
  assign pht_0_7_MPORT_993_en = reset;
  assign pht_0_7_MPORT_995_data = 1'h0;
  assign pht_0_7_MPORT_995_addr = 6'h19;
  assign pht_0_7_MPORT_995_mask = 1'h1;
  assign pht_0_7_MPORT_995_en = reset;
  assign pht_0_7_MPORT_997_data = 1'h0;
  assign pht_0_7_MPORT_997_addr = 6'h1a;
  assign pht_0_7_MPORT_997_mask = 1'h1;
  assign pht_0_7_MPORT_997_en = reset;
  assign pht_0_7_MPORT_999_data = 1'h0;
  assign pht_0_7_MPORT_999_addr = 6'h1b;
  assign pht_0_7_MPORT_999_mask = 1'h1;
  assign pht_0_7_MPORT_999_en = reset;
  assign pht_0_7_MPORT_1001_data = 1'h0;
  assign pht_0_7_MPORT_1001_addr = 6'h1c;
  assign pht_0_7_MPORT_1001_mask = 1'h1;
  assign pht_0_7_MPORT_1001_en = reset;
  assign pht_0_7_MPORT_1003_data = 1'h0;
  assign pht_0_7_MPORT_1003_addr = 6'h1d;
  assign pht_0_7_MPORT_1003_mask = 1'h1;
  assign pht_0_7_MPORT_1003_en = reset;
  assign pht_0_7_MPORT_1005_data = 1'h0;
  assign pht_0_7_MPORT_1005_addr = 6'h1e;
  assign pht_0_7_MPORT_1005_mask = 1'h1;
  assign pht_0_7_MPORT_1005_en = reset;
  assign pht_0_7_MPORT_1007_data = 1'h0;
  assign pht_0_7_MPORT_1007_addr = 6'h1f;
  assign pht_0_7_MPORT_1007_mask = 1'h1;
  assign pht_0_7_MPORT_1007_en = reset;
  assign pht_0_7_MPORT_1009_data = 1'h0;
  assign pht_0_7_MPORT_1009_addr = 6'h20;
  assign pht_0_7_MPORT_1009_mask = 1'h1;
  assign pht_0_7_MPORT_1009_en = reset;
  assign pht_0_7_MPORT_1011_data = 1'h0;
  assign pht_0_7_MPORT_1011_addr = 6'h21;
  assign pht_0_7_MPORT_1011_mask = 1'h1;
  assign pht_0_7_MPORT_1011_en = reset;
  assign pht_0_7_MPORT_1013_data = 1'h0;
  assign pht_0_7_MPORT_1013_addr = 6'h22;
  assign pht_0_7_MPORT_1013_mask = 1'h1;
  assign pht_0_7_MPORT_1013_en = reset;
  assign pht_0_7_MPORT_1015_data = 1'h0;
  assign pht_0_7_MPORT_1015_addr = 6'h23;
  assign pht_0_7_MPORT_1015_mask = 1'h1;
  assign pht_0_7_MPORT_1015_en = reset;
  assign pht_0_7_MPORT_1017_data = 1'h0;
  assign pht_0_7_MPORT_1017_addr = 6'h24;
  assign pht_0_7_MPORT_1017_mask = 1'h1;
  assign pht_0_7_MPORT_1017_en = reset;
  assign pht_0_7_MPORT_1019_data = 1'h0;
  assign pht_0_7_MPORT_1019_addr = 6'h25;
  assign pht_0_7_MPORT_1019_mask = 1'h1;
  assign pht_0_7_MPORT_1019_en = reset;
  assign pht_0_7_MPORT_1021_data = 1'h0;
  assign pht_0_7_MPORT_1021_addr = 6'h26;
  assign pht_0_7_MPORT_1021_mask = 1'h1;
  assign pht_0_7_MPORT_1021_en = reset;
  assign pht_0_7_MPORT_1023_data = 1'h0;
  assign pht_0_7_MPORT_1023_addr = 6'h27;
  assign pht_0_7_MPORT_1023_mask = 1'h1;
  assign pht_0_7_MPORT_1023_en = reset;
  assign pht_0_7_MPORT_1025_data = 1'h0;
  assign pht_0_7_MPORT_1025_addr = 6'h28;
  assign pht_0_7_MPORT_1025_mask = 1'h1;
  assign pht_0_7_MPORT_1025_en = reset;
  assign pht_0_7_MPORT_1027_data = 1'h0;
  assign pht_0_7_MPORT_1027_addr = 6'h29;
  assign pht_0_7_MPORT_1027_mask = 1'h1;
  assign pht_0_7_MPORT_1027_en = reset;
  assign pht_0_7_MPORT_1029_data = 1'h0;
  assign pht_0_7_MPORT_1029_addr = 6'h2a;
  assign pht_0_7_MPORT_1029_mask = 1'h1;
  assign pht_0_7_MPORT_1029_en = reset;
  assign pht_0_7_MPORT_1031_data = 1'h0;
  assign pht_0_7_MPORT_1031_addr = 6'h2b;
  assign pht_0_7_MPORT_1031_mask = 1'h1;
  assign pht_0_7_MPORT_1031_en = reset;
  assign pht_0_7_MPORT_1033_data = 1'h0;
  assign pht_0_7_MPORT_1033_addr = 6'h2c;
  assign pht_0_7_MPORT_1033_mask = 1'h1;
  assign pht_0_7_MPORT_1033_en = reset;
  assign pht_0_7_MPORT_1035_data = 1'h0;
  assign pht_0_7_MPORT_1035_addr = 6'h2d;
  assign pht_0_7_MPORT_1035_mask = 1'h1;
  assign pht_0_7_MPORT_1035_en = reset;
  assign pht_0_7_MPORT_1037_data = 1'h0;
  assign pht_0_7_MPORT_1037_addr = 6'h2e;
  assign pht_0_7_MPORT_1037_mask = 1'h1;
  assign pht_0_7_MPORT_1037_en = reset;
  assign pht_0_7_MPORT_1039_data = 1'h0;
  assign pht_0_7_MPORT_1039_addr = 6'h2f;
  assign pht_0_7_MPORT_1039_mask = 1'h1;
  assign pht_0_7_MPORT_1039_en = reset;
  assign pht_0_7_MPORT_1041_data = 1'h0;
  assign pht_0_7_MPORT_1041_addr = 6'h30;
  assign pht_0_7_MPORT_1041_mask = 1'h1;
  assign pht_0_7_MPORT_1041_en = reset;
  assign pht_0_7_MPORT_1043_data = 1'h0;
  assign pht_0_7_MPORT_1043_addr = 6'h31;
  assign pht_0_7_MPORT_1043_mask = 1'h1;
  assign pht_0_7_MPORT_1043_en = reset;
  assign pht_0_7_MPORT_1045_data = 1'h0;
  assign pht_0_7_MPORT_1045_addr = 6'h32;
  assign pht_0_7_MPORT_1045_mask = 1'h1;
  assign pht_0_7_MPORT_1045_en = reset;
  assign pht_0_7_MPORT_1047_data = 1'h0;
  assign pht_0_7_MPORT_1047_addr = 6'h33;
  assign pht_0_7_MPORT_1047_mask = 1'h1;
  assign pht_0_7_MPORT_1047_en = reset;
  assign pht_0_7_MPORT_1049_data = 1'h0;
  assign pht_0_7_MPORT_1049_addr = 6'h34;
  assign pht_0_7_MPORT_1049_mask = 1'h1;
  assign pht_0_7_MPORT_1049_en = reset;
  assign pht_0_7_MPORT_1051_data = 1'h0;
  assign pht_0_7_MPORT_1051_addr = 6'h35;
  assign pht_0_7_MPORT_1051_mask = 1'h1;
  assign pht_0_7_MPORT_1051_en = reset;
  assign pht_0_7_MPORT_1053_data = 1'h0;
  assign pht_0_7_MPORT_1053_addr = 6'h36;
  assign pht_0_7_MPORT_1053_mask = 1'h1;
  assign pht_0_7_MPORT_1053_en = reset;
  assign pht_0_7_MPORT_1055_data = 1'h0;
  assign pht_0_7_MPORT_1055_addr = 6'h37;
  assign pht_0_7_MPORT_1055_mask = 1'h1;
  assign pht_0_7_MPORT_1055_en = reset;
  assign pht_0_7_MPORT_1057_data = 1'h0;
  assign pht_0_7_MPORT_1057_addr = 6'h38;
  assign pht_0_7_MPORT_1057_mask = 1'h1;
  assign pht_0_7_MPORT_1057_en = reset;
  assign pht_0_7_MPORT_1059_data = 1'h0;
  assign pht_0_7_MPORT_1059_addr = 6'h39;
  assign pht_0_7_MPORT_1059_mask = 1'h1;
  assign pht_0_7_MPORT_1059_en = reset;
  assign pht_0_7_MPORT_1061_data = 1'h0;
  assign pht_0_7_MPORT_1061_addr = 6'h3a;
  assign pht_0_7_MPORT_1061_mask = 1'h1;
  assign pht_0_7_MPORT_1061_en = reset;
  assign pht_0_7_MPORT_1063_data = 1'h0;
  assign pht_0_7_MPORT_1063_addr = 6'h3b;
  assign pht_0_7_MPORT_1063_mask = 1'h1;
  assign pht_0_7_MPORT_1063_en = reset;
  assign pht_0_7_MPORT_1065_data = 1'h0;
  assign pht_0_7_MPORT_1065_addr = 6'h3c;
  assign pht_0_7_MPORT_1065_mask = 1'h1;
  assign pht_0_7_MPORT_1065_en = reset;
  assign pht_0_7_MPORT_1067_data = 1'h0;
  assign pht_0_7_MPORT_1067_addr = 6'h3d;
  assign pht_0_7_MPORT_1067_mask = 1'h1;
  assign pht_0_7_MPORT_1067_en = reset;
  assign pht_0_7_MPORT_1069_data = 1'h0;
  assign pht_0_7_MPORT_1069_addr = 6'h3e;
  assign pht_0_7_MPORT_1069_mask = 1'h1;
  assign pht_0_7_MPORT_1069_en = reset;
  assign pht_0_7_MPORT_1071_data = 1'h0;
  assign pht_0_7_MPORT_1071_addr = 6'h3f;
  assign pht_0_7_MPORT_1071_mask = 1'h1;
  assign pht_0_7_MPORT_1071_en = reset;
  assign io_rdirect_0 = REG_7 == 3'h7 ? pht_1_7_MPORT_7_data : _GEN_17; // @[PatternHistoryTable.scala 42:44 43:23]
  assign io_rdirect_1 = REG_15 == 3'h7 ? pht_1_7_MPORT_15_data : _GEN_34; // @[PatternHistoryTable.scala 42:44 43:23]
  always @(posedge clock) begin
    if (pht_1_0_MPORT_32_en & pht_1_0_MPORT_32_mask) begin
      pht_1_0[pht_1_0_MPORT_32_addr] <= pht_1_0_MPORT_32_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_48_en & pht_1_0_MPORT_48_mask) begin
      pht_1_0[pht_1_0_MPORT_48_addr] <= pht_1_0_MPORT_48_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_50_en & pht_1_0_MPORT_50_mask) begin
      pht_1_0[pht_1_0_MPORT_50_addr] <= pht_1_0_MPORT_50_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_52_en & pht_1_0_MPORT_52_mask) begin
      pht_1_0[pht_1_0_MPORT_52_addr] <= pht_1_0_MPORT_52_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_54_en & pht_1_0_MPORT_54_mask) begin
      pht_1_0[pht_1_0_MPORT_54_addr] <= pht_1_0_MPORT_54_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_56_en & pht_1_0_MPORT_56_mask) begin
      pht_1_0[pht_1_0_MPORT_56_addr] <= pht_1_0_MPORT_56_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_58_en & pht_1_0_MPORT_58_mask) begin
      pht_1_0[pht_1_0_MPORT_58_addr] <= pht_1_0_MPORT_58_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_60_en & pht_1_0_MPORT_60_mask) begin
      pht_1_0[pht_1_0_MPORT_60_addr] <= pht_1_0_MPORT_60_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_62_en & pht_1_0_MPORT_62_mask) begin
      pht_1_0[pht_1_0_MPORT_62_addr] <= pht_1_0_MPORT_62_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_64_en & pht_1_0_MPORT_64_mask) begin
      pht_1_0[pht_1_0_MPORT_64_addr] <= pht_1_0_MPORT_64_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_66_en & pht_1_0_MPORT_66_mask) begin
      pht_1_0[pht_1_0_MPORT_66_addr] <= pht_1_0_MPORT_66_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_68_en & pht_1_0_MPORT_68_mask) begin
      pht_1_0[pht_1_0_MPORT_68_addr] <= pht_1_0_MPORT_68_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_70_en & pht_1_0_MPORT_70_mask) begin
      pht_1_0[pht_1_0_MPORT_70_addr] <= pht_1_0_MPORT_70_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_72_en & pht_1_0_MPORT_72_mask) begin
      pht_1_0[pht_1_0_MPORT_72_addr] <= pht_1_0_MPORT_72_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_74_en & pht_1_0_MPORT_74_mask) begin
      pht_1_0[pht_1_0_MPORT_74_addr] <= pht_1_0_MPORT_74_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_76_en & pht_1_0_MPORT_76_mask) begin
      pht_1_0[pht_1_0_MPORT_76_addr] <= pht_1_0_MPORT_76_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_78_en & pht_1_0_MPORT_78_mask) begin
      pht_1_0[pht_1_0_MPORT_78_addr] <= pht_1_0_MPORT_78_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_80_en & pht_1_0_MPORT_80_mask) begin
      pht_1_0[pht_1_0_MPORT_80_addr] <= pht_1_0_MPORT_80_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_82_en & pht_1_0_MPORT_82_mask) begin
      pht_1_0[pht_1_0_MPORT_82_addr] <= pht_1_0_MPORT_82_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_84_en & pht_1_0_MPORT_84_mask) begin
      pht_1_0[pht_1_0_MPORT_84_addr] <= pht_1_0_MPORT_84_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_86_en & pht_1_0_MPORT_86_mask) begin
      pht_1_0[pht_1_0_MPORT_86_addr] <= pht_1_0_MPORT_86_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_88_en & pht_1_0_MPORT_88_mask) begin
      pht_1_0[pht_1_0_MPORT_88_addr] <= pht_1_0_MPORT_88_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_90_en & pht_1_0_MPORT_90_mask) begin
      pht_1_0[pht_1_0_MPORT_90_addr] <= pht_1_0_MPORT_90_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_92_en & pht_1_0_MPORT_92_mask) begin
      pht_1_0[pht_1_0_MPORT_92_addr] <= pht_1_0_MPORT_92_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_94_en & pht_1_0_MPORT_94_mask) begin
      pht_1_0[pht_1_0_MPORT_94_addr] <= pht_1_0_MPORT_94_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_96_en & pht_1_0_MPORT_96_mask) begin
      pht_1_0[pht_1_0_MPORT_96_addr] <= pht_1_0_MPORT_96_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_98_en & pht_1_0_MPORT_98_mask) begin
      pht_1_0[pht_1_0_MPORT_98_addr] <= pht_1_0_MPORT_98_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_100_en & pht_1_0_MPORT_100_mask) begin
      pht_1_0[pht_1_0_MPORT_100_addr] <= pht_1_0_MPORT_100_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_102_en & pht_1_0_MPORT_102_mask) begin
      pht_1_0[pht_1_0_MPORT_102_addr] <= pht_1_0_MPORT_102_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_104_en & pht_1_0_MPORT_104_mask) begin
      pht_1_0[pht_1_0_MPORT_104_addr] <= pht_1_0_MPORT_104_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_106_en & pht_1_0_MPORT_106_mask) begin
      pht_1_0[pht_1_0_MPORT_106_addr] <= pht_1_0_MPORT_106_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_108_en & pht_1_0_MPORT_108_mask) begin
      pht_1_0[pht_1_0_MPORT_108_addr] <= pht_1_0_MPORT_108_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_110_en & pht_1_0_MPORT_110_mask) begin
      pht_1_0[pht_1_0_MPORT_110_addr] <= pht_1_0_MPORT_110_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_112_en & pht_1_0_MPORT_112_mask) begin
      pht_1_0[pht_1_0_MPORT_112_addr] <= pht_1_0_MPORT_112_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_114_en & pht_1_0_MPORT_114_mask) begin
      pht_1_0[pht_1_0_MPORT_114_addr] <= pht_1_0_MPORT_114_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_116_en & pht_1_0_MPORT_116_mask) begin
      pht_1_0[pht_1_0_MPORT_116_addr] <= pht_1_0_MPORT_116_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_118_en & pht_1_0_MPORT_118_mask) begin
      pht_1_0[pht_1_0_MPORT_118_addr] <= pht_1_0_MPORT_118_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_120_en & pht_1_0_MPORT_120_mask) begin
      pht_1_0[pht_1_0_MPORT_120_addr] <= pht_1_0_MPORT_120_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_122_en & pht_1_0_MPORT_122_mask) begin
      pht_1_0[pht_1_0_MPORT_122_addr] <= pht_1_0_MPORT_122_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_124_en & pht_1_0_MPORT_124_mask) begin
      pht_1_0[pht_1_0_MPORT_124_addr] <= pht_1_0_MPORT_124_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_126_en & pht_1_0_MPORT_126_mask) begin
      pht_1_0[pht_1_0_MPORT_126_addr] <= pht_1_0_MPORT_126_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_128_en & pht_1_0_MPORT_128_mask) begin
      pht_1_0[pht_1_0_MPORT_128_addr] <= pht_1_0_MPORT_128_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_130_en & pht_1_0_MPORT_130_mask) begin
      pht_1_0[pht_1_0_MPORT_130_addr] <= pht_1_0_MPORT_130_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_132_en & pht_1_0_MPORT_132_mask) begin
      pht_1_0[pht_1_0_MPORT_132_addr] <= pht_1_0_MPORT_132_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_134_en & pht_1_0_MPORT_134_mask) begin
      pht_1_0[pht_1_0_MPORT_134_addr] <= pht_1_0_MPORT_134_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_136_en & pht_1_0_MPORT_136_mask) begin
      pht_1_0[pht_1_0_MPORT_136_addr] <= pht_1_0_MPORT_136_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_138_en & pht_1_0_MPORT_138_mask) begin
      pht_1_0[pht_1_0_MPORT_138_addr] <= pht_1_0_MPORT_138_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_140_en & pht_1_0_MPORT_140_mask) begin
      pht_1_0[pht_1_0_MPORT_140_addr] <= pht_1_0_MPORT_140_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_142_en & pht_1_0_MPORT_142_mask) begin
      pht_1_0[pht_1_0_MPORT_142_addr] <= pht_1_0_MPORT_142_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_144_en & pht_1_0_MPORT_144_mask) begin
      pht_1_0[pht_1_0_MPORT_144_addr] <= pht_1_0_MPORT_144_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_146_en & pht_1_0_MPORT_146_mask) begin
      pht_1_0[pht_1_0_MPORT_146_addr] <= pht_1_0_MPORT_146_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_148_en & pht_1_0_MPORT_148_mask) begin
      pht_1_0[pht_1_0_MPORT_148_addr] <= pht_1_0_MPORT_148_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_150_en & pht_1_0_MPORT_150_mask) begin
      pht_1_0[pht_1_0_MPORT_150_addr] <= pht_1_0_MPORT_150_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_152_en & pht_1_0_MPORT_152_mask) begin
      pht_1_0[pht_1_0_MPORT_152_addr] <= pht_1_0_MPORT_152_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_154_en & pht_1_0_MPORT_154_mask) begin
      pht_1_0[pht_1_0_MPORT_154_addr] <= pht_1_0_MPORT_154_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_156_en & pht_1_0_MPORT_156_mask) begin
      pht_1_0[pht_1_0_MPORT_156_addr] <= pht_1_0_MPORT_156_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_158_en & pht_1_0_MPORT_158_mask) begin
      pht_1_0[pht_1_0_MPORT_158_addr] <= pht_1_0_MPORT_158_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_160_en & pht_1_0_MPORT_160_mask) begin
      pht_1_0[pht_1_0_MPORT_160_addr] <= pht_1_0_MPORT_160_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_162_en & pht_1_0_MPORT_162_mask) begin
      pht_1_0[pht_1_0_MPORT_162_addr] <= pht_1_0_MPORT_162_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_164_en & pht_1_0_MPORT_164_mask) begin
      pht_1_0[pht_1_0_MPORT_164_addr] <= pht_1_0_MPORT_164_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_166_en & pht_1_0_MPORT_166_mask) begin
      pht_1_0[pht_1_0_MPORT_166_addr] <= pht_1_0_MPORT_166_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_168_en & pht_1_0_MPORT_168_mask) begin
      pht_1_0[pht_1_0_MPORT_168_addr] <= pht_1_0_MPORT_168_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_170_en & pht_1_0_MPORT_170_mask) begin
      pht_1_0[pht_1_0_MPORT_170_addr] <= pht_1_0_MPORT_170_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_172_en & pht_1_0_MPORT_172_mask) begin
      pht_1_0[pht_1_0_MPORT_172_addr] <= pht_1_0_MPORT_172_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_0_MPORT_174_en & pht_1_0_MPORT_174_mask) begin
      pht_1_0[pht_1_0_MPORT_174_addr] <= pht_1_0_MPORT_174_data; // @[PatternHistoryTable.scala 21:28]
    end
//     pht_1_0_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_0_MPORT_addr_pipe_0 <= io_raddr_0;
    end
//     pht_1_0_MPORT_8_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_0_MPORT_8_addr_pipe_0 <= io_raddr_1;
    end
//     pht_1_0_MPORT_16_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_0_MPORT_16_addr_pipe_0 <= io_waddr;
    end
    if (pht_1_1_MPORT_34_en & pht_1_1_MPORT_34_mask) begin
      pht_1_1[pht_1_1_MPORT_34_addr] <= pht_1_1_MPORT_34_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_176_en & pht_1_1_MPORT_176_mask) begin
      pht_1_1[pht_1_1_MPORT_176_addr] <= pht_1_1_MPORT_176_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_178_en & pht_1_1_MPORT_178_mask) begin
      pht_1_1[pht_1_1_MPORT_178_addr] <= pht_1_1_MPORT_178_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_180_en & pht_1_1_MPORT_180_mask) begin
      pht_1_1[pht_1_1_MPORT_180_addr] <= pht_1_1_MPORT_180_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_182_en & pht_1_1_MPORT_182_mask) begin
      pht_1_1[pht_1_1_MPORT_182_addr] <= pht_1_1_MPORT_182_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_184_en & pht_1_1_MPORT_184_mask) begin
      pht_1_1[pht_1_1_MPORT_184_addr] <= pht_1_1_MPORT_184_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_186_en & pht_1_1_MPORT_186_mask) begin
      pht_1_1[pht_1_1_MPORT_186_addr] <= pht_1_1_MPORT_186_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_188_en & pht_1_1_MPORT_188_mask) begin
      pht_1_1[pht_1_1_MPORT_188_addr] <= pht_1_1_MPORT_188_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_190_en & pht_1_1_MPORT_190_mask) begin
      pht_1_1[pht_1_1_MPORT_190_addr] <= pht_1_1_MPORT_190_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_192_en & pht_1_1_MPORT_192_mask) begin
      pht_1_1[pht_1_1_MPORT_192_addr] <= pht_1_1_MPORT_192_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_194_en & pht_1_1_MPORT_194_mask) begin
      pht_1_1[pht_1_1_MPORT_194_addr] <= pht_1_1_MPORT_194_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_196_en & pht_1_1_MPORT_196_mask) begin
      pht_1_1[pht_1_1_MPORT_196_addr] <= pht_1_1_MPORT_196_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_198_en & pht_1_1_MPORT_198_mask) begin
      pht_1_1[pht_1_1_MPORT_198_addr] <= pht_1_1_MPORT_198_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_200_en & pht_1_1_MPORT_200_mask) begin
      pht_1_1[pht_1_1_MPORT_200_addr] <= pht_1_1_MPORT_200_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_202_en & pht_1_1_MPORT_202_mask) begin
      pht_1_1[pht_1_1_MPORT_202_addr] <= pht_1_1_MPORT_202_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_204_en & pht_1_1_MPORT_204_mask) begin
      pht_1_1[pht_1_1_MPORT_204_addr] <= pht_1_1_MPORT_204_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_206_en & pht_1_1_MPORT_206_mask) begin
      pht_1_1[pht_1_1_MPORT_206_addr] <= pht_1_1_MPORT_206_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_208_en & pht_1_1_MPORT_208_mask) begin
      pht_1_1[pht_1_1_MPORT_208_addr] <= pht_1_1_MPORT_208_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_210_en & pht_1_1_MPORT_210_mask) begin
      pht_1_1[pht_1_1_MPORT_210_addr] <= pht_1_1_MPORT_210_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_212_en & pht_1_1_MPORT_212_mask) begin
      pht_1_1[pht_1_1_MPORT_212_addr] <= pht_1_1_MPORT_212_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_214_en & pht_1_1_MPORT_214_mask) begin
      pht_1_1[pht_1_1_MPORT_214_addr] <= pht_1_1_MPORT_214_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_216_en & pht_1_1_MPORT_216_mask) begin
      pht_1_1[pht_1_1_MPORT_216_addr] <= pht_1_1_MPORT_216_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_218_en & pht_1_1_MPORT_218_mask) begin
      pht_1_1[pht_1_1_MPORT_218_addr] <= pht_1_1_MPORT_218_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_220_en & pht_1_1_MPORT_220_mask) begin
      pht_1_1[pht_1_1_MPORT_220_addr] <= pht_1_1_MPORT_220_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_222_en & pht_1_1_MPORT_222_mask) begin
      pht_1_1[pht_1_1_MPORT_222_addr] <= pht_1_1_MPORT_222_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_224_en & pht_1_1_MPORT_224_mask) begin
      pht_1_1[pht_1_1_MPORT_224_addr] <= pht_1_1_MPORT_224_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_226_en & pht_1_1_MPORT_226_mask) begin
      pht_1_1[pht_1_1_MPORT_226_addr] <= pht_1_1_MPORT_226_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_228_en & pht_1_1_MPORT_228_mask) begin
      pht_1_1[pht_1_1_MPORT_228_addr] <= pht_1_1_MPORT_228_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_230_en & pht_1_1_MPORT_230_mask) begin
      pht_1_1[pht_1_1_MPORT_230_addr] <= pht_1_1_MPORT_230_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_232_en & pht_1_1_MPORT_232_mask) begin
      pht_1_1[pht_1_1_MPORT_232_addr] <= pht_1_1_MPORT_232_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_234_en & pht_1_1_MPORT_234_mask) begin
      pht_1_1[pht_1_1_MPORT_234_addr] <= pht_1_1_MPORT_234_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_236_en & pht_1_1_MPORT_236_mask) begin
      pht_1_1[pht_1_1_MPORT_236_addr] <= pht_1_1_MPORT_236_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_238_en & pht_1_1_MPORT_238_mask) begin
      pht_1_1[pht_1_1_MPORT_238_addr] <= pht_1_1_MPORT_238_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_240_en & pht_1_1_MPORT_240_mask) begin
      pht_1_1[pht_1_1_MPORT_240_addr] <= pht_1_1_MPORT_240_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_242_en & pht_1_1_MPORT_242_mask) begin
      pht_1_1[pht_1_1_MPORT_242_addr] <= pht_1_1_MPORT_242_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_244_en & pht_1_1_MPORT_244_mask) begin
      pht_1_1[pht_1_1_MPORT_244_addr] <= pht_1_1_MPORT_244_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_246_en & pht_1_1_MPORT_246_mask) begin
      pht_1_1[pht_1_1_MPORT_246_addr] <= pht_1_1_MPORT_246_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_248_en & pht_1_1_MPORT_248_mask) begin
      pht_1_1[pht_1_1_MPORT_248_addr] <= pht_1_1_MPORT_248_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_250_en & pht_1_1_MPORT_250_mask) begin
      pht_1_1[pht_1_1_MPORT_250_addr] <= pht_1_1_MPORT_250_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_252_en & pht_1_1_MPORT_252_mask) begin
      pht_1_1[pht_1_1_MPORT_252_addr] <= pht_1_1_MPORT_252_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_254_en & pht_1_1_MPORT_254_mask) begin
      pht_1_1[pht_1_1_MPORT_254_addr] <= pht_1_1_MPORT_254_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_256_en & pht_1_1_MPORT_256_mask) begin
      pht_1_1[pht_1_1_MPORT_256_addr] <= pht_1_1_MPORT_256_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_258_en & pht_1_1_MPORT_258_mask) begin
      pht_1_1[pht_1_1_MPORT_258_addr] <= pht_1_1_MPORT_258_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_260_en & pht_1_1_MPORT_260_mask) begin
      pht_1_1[pht_1_1_MPORT_260_addr] <= pht_1_1_MPORT_260_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_262_en & pht_1_1_MPORT_262_mask) begin
      pht_1_1[pht_1_1_MPORT_262_addr] <= pht_1_1_MPORT_262_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_264_en & pht_1_1_MPORT_264_mask) begin
      pht_1_1[pht_1_1_MPORT_264_addr] <= pht_1_1_MPORT_264_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_266_en & pht_1_1_MPORT_266_mask) begin
      pht_1_1[pht_1_1_MPORT_266_addr] <= pht_1_1_MPORT_266_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_268_en & pht_1_1_MPORT_268_mask) begin
      pht_1_1[pht_1_1_MPORT_268_addr] <= pht_1_1_MPORT_268_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_270_en & pht_1_1_MPORT_270_mask) begin
      pht_1_1[pht_1_1_MPORT_270_addr] <= pht_1_1_MPORT_270_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_272_en & pht_1_1_MPORT_272_mask) begin
      pht_1_1[pht_1_1_MPORT_272_addr] <= pht_1_1_MPORT_272_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_274_en & pht_1_1_MPORT_274_mask) begin
      pht_1_1[pht_1_1_MPORT_274_addr] <= pht_1_1_MPORT_274_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_276_en & pht_1_1_MPORT_276_mask) begin
      pht_1_1[pht_1_1_MPORT_276_addr] <= pht_1_1_MPORT_276_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_278_en & pht_1_1_MPORT_278_mask) begin
      pht_1_1[pht_1_1_MPORT_278_addr] <= pht_1_1_MPORT_278_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_280_en & pht_1_1_MPORT_280_mask) begin
      pht_1_1[pht_1_1_MPORT_280_addr] <= pht_1_1_MPORT_280_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_282_en & pht_1_1_MPORT_282_mask) begin
      pht_1_1[pht_1_1_MPORT_282_addr] <= pht_1_1_MPORT_282_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_284_en & pht_1_1_MPORT_284_mask) begin
      pht_1_1[pht_1_1_MPORT_284_addr] <= pht_1_1_MPORT_284_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_286_en & pht_1_1_MPORT_286_mask) begin
      pht_1_1[pht_1_1_MPORT_286_addr] <= pht_1_1_MPORT_286_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_288_en & pht_1_1_MPORT_288_mask) begin
      pht_1_1[pht_1_1_MPORT_288_addr] <= pht_1_1_MPORT_288_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_290_en & pht_1_1_MPORT_290_mask) begin
      pht_1_1[pht_1_1_MPORT_290_addr] <= pht_1_1_MPORT_290_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_292_en & pht_1_1_MPORT_292_mask) begin
      pht_1_1[pht_1_1_MPORT_292_addr] <= pht_1_1_MPORT_292_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_294_en & pht_1_1_MPORT_294_mask) begin
      pht_1_1[pht_1_1_MPORT_294_addr] <= pht_1_1_MPORT_294_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_296_en & pht_1_1_MPORT_296_mask) begin
      pht_1_1[pht_1_1_MPORT_296_addr] <= pht_1_1_MPORT_296_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_298_en & pht_1_1_MPORT_298_mask) begin
      pht_1_1[pht_1_1_MPORT_298_addr] <= pht_1_1_MPORT_298_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_300_en & pht_1_1_MPORT_300_mask) begin
      pht_1_1[pht_1_1_MPORT_300_addr] <= pht_1_1_MPORT_300_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_1_MPORT_302_en & pht_1_1_MPORT_302_mask) begin
      pht_1_1[pht_1_1_MPORT_302_addr] <= pht_1_1_MPORT_302_data; // @[PatternHistoryTable.scala 21:28]
    end
//     pht_1_1_MPORT_1_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_1_MPORT_1_addr_pipe_0 <= io_raddr_0;
    end
//     pht_1_1_MPORT_9_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_1_MPORT_9_addr_pipe_0 <= io_raddr_1;
    end
//     pht_1_1_MPORT_18_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_1_MPORT_18_addr_pipe_0 <= io_waddr;
    end
    if (pht_1_2_MPORT_36_en & pht_1_2_MPORT_36_mask) begin
      pht_1_2[pht_1_2_MPORT_36_addr] <= pht_1_2_MPORT_36_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_304_en & pht_1_2_MPORT_304_mask) begin
      pht_1_2[pht_1_2_MPORT_304_addr] <= pht_1_2_MPORT_304_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_306_en & pht_1_2_MPORT_306_mask) begin
      pht_1_2[pht_1_2_MPORT_306_addr] <= pht_1_2_MPORT_306_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_308_en & pht_1_2_MPORT_308_mask) begin
      pht_1_2[pht_1_2_MPORT_308_addr] <= pht_1_2_MPORT_308_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_310_en & pht_1_2_MPORT_310_mask) begin
      pht_1_2[pht_1_2_MPORT_310_addr] <= pht_1_2_MPORT_310_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_312_en & pht_1_2_MPORT_312_mask) begin
      pht_1_2[pht_1_2_MPORT_312_addr] <= pht_1_2_MPORT_312_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_314_en & pht_1_2_MPORT_314_mask) begin
      pht_1_2[pht_1_2_MPORT_314_addr] <= pht_1_2_MPORT_314_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_316_en & pht_1_2_MPORT_316_mask) begin
      pht_1_2[pht_1_2_MPORT_316_addr] <= pht_1_2_MPORT_316_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_318_en & pht_1_2_MPORT_318_mask) begin
      pht_1_2[pht_1_2_MPORT_318_addr] <= pht_1_2_MPORT_318_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_320_en & pht_1_2_MPORT_320_mask) begin
      pht_1_2[pht_1_2_MPORT_320_addr] <= pht_1_2_MPORT_320_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_322_en & pht_1_2_MPORT_322_mask) begin
      pht_1_2[pht_1_2_MPORT_322_addr] <= pht_1_2_MPORT_322_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_324_en & pht_1_2_MPORT_324_mask) begin
      pht_1_2[pht_1_2_MPORT_324_addr] <= pht_1_2_MPORT_324_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_326_en & pht_1_2_MPORT_326_mask) begin
      pht_1_2[pht_1_2_MPORT_326_addr] <= pht_1_2_MPORT_326_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_328_en & pht_1_2_MPORT_328_mask) begin
      pht_1_2[pht_1_2_MPORT_328_addr] <= pht_1_2_MPORT_328_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_330_en & pht_1_2_MPORT_330_mask) begin
      pht_1_2[pht_1_2_MPORT_330_addr] <= pht_1_2_MPORT_330_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_332_en & pht_1_2_MPORT_332_mask) begin
      pht_1_2[pht_1_2_MPORT_332_addr] <= pht_1_2_MPORT_332_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_334_en & pht_1_2_MPORT_334_mask) begin
      pht_1_2[pht_1_2_MPORT_334_addr] <= pht_1_2_MPORT_334_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_336_en & pht_1_2_MPORT_336_mask) begin
      pht_1_2[pht_1_2_MPORT_336_addr] <= pht_1_2_MPORT_336_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_338_en & pht_1_2_MPORT_338_mask) begin
      pht_1_2[pht_1_2_MPORT_338_addr] <= pht_1_2_MPORT_338_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_340_en & pht_1_2_MPORT_340_mask) begin
      pht_1_2[pht_1_2_MPORT_340_addr] <= pht_1_2_MPORT_340_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_342_en & pht_1_2_MPORT_342_mask) begin
      pht_1_2[pht_1_2_MPORT_342_addr] <= pht_1_2_MPORT_342_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_344_en & pht_1_2_MPORT_344_mask) begin
      pht_1_2[pht_1_2_MPORT_344_addr] <= pht_1_2_MPORT_344_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_346_en & pht_1_2_MPORT_346_mask) begin
      pht_1_2[pht_1_2_MPORT_346_addr] <= pht_1_2_MPORT_346_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_348_en & pht_1_2_MPORT_348_mask) begin
      pht_1_2[pht_1_2_MPORT_348_addr] <= pht_1_2_MPORT_348_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_350_en & pht_1_2_MPORT_350_mask) begin
      pht_1_2[pht_1_2_MPORT_350_addr] <= pht_1_2_MPORT_350_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_352_en & pht_1_2_MPORT_352_mask) begin
      pht_1_2[pht_1_2_MPORT_352_addr] <= pht_1_2_MPORT_352_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_354_en & pht_1_2_MPORT_354_mask) begin
      pht_1_2[pht_1_2_MPORT_354_addr] <= pht_1_2_MPORT_354_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_356_en & pht_1_2_MPORT_356_mask) begin
      pht_1_2[pht_1_2_MPORT_356_addr] <= pht_1_2_MPORT_356_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_358_en & pht_1_2_MPORT_358_mask) begin
      pht_1_2[pht_1_2_MPORT_358_addr] <= pht_1_2_MPORT_358_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_360_en & pht_1_2_MPORT_360_mask) begin
      pht_1_2[pht_1_2_MPORT_360_addr] <= pht_1_2_MPORT_360_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_362_en & pht_1_2_MPORT_362_mask) begin
      pht_1_2[pht_1_2_MPORT_362_addr] <= pht_1_2_MPORT_362_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_364_en & pht_1_2_MPORT_364_mask) begin
      pht_1_2[pht_1_2_MPORT_364_addr] <= pht_1_2_MPORT_364_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_366_en & pht_1_2_MPORT_366_mask) begin
      pht_1_2[pht_1_2_MPORT_366_addr] <= pht_1_2_MPORT_366_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_368_en & pht_1_2_MPORT_368_mask) begin
      pht_1_2[pht_1_2_MPORT_368_addr] <= pht_1_2_MPORT_368_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_370_en & pht_1_2_MPORT_370_mask) begin
      pht_1_2[pht_1_2_MPORT_370_addr] <= pht_1_2_MPORT_370_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_372_en & pht_1_2_MPORT_372_mask) begin
      pht_1_2[pht_1_2_MPORT_372_addr] <= pht_1_2_MPORT_372_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_374_en & pht_1_2_MPORT_374_mask) begin
      pht_1_2[pht_1_2_MPORT_374_addr] <= pht_1_2_MPORT_374_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_376_en & pht_1_2_MPORT_376_mask) begin
      pht_1_2[pht_1_2_MPORT_376_addr] <= pht_1_2_MPORT_376_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_378_en & pht_1_2_MPORT_378_mask) begin
      pht_1_2[pht_1_2_MPORT_378_addr] <= pht_1_2_MPORT_378_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_380_en & pht_1_2_MPORT_380_mask) begin
      pht_1_2[pht_1_2_MPORT_380_addr] <= pht_1_2_MPORT_380_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_382_en & pht_1_2_MPORT_382_mask) begin
      pht_1_2[pht_1_2_MPORT_382_addr] <= pht_1_2_MPORT_382_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_384_en & pht_1_2_MPORT_384_mask) begin
      pht_1_2[pht_1_2_MPORT_384_addr] <= pht_1_2_MPORT_384_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_386_en & pht_1_2_MPORT_386_mask) begin
      pht_1_2[pht_1_2_MPORT_386_addr] <= pht_1_2_MPORT_386_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_388_en & pht_1_2_MPORT_388_mask) begin
      pht_1_2[pht_1_2_MPORT_388_addr] <= pht_1_2_MPORT_388_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_390_en & pht_1_2_MPORT_390_mask) begin
      pht_1_2[pht_1_2_MPORT_390_addr] <= pht_1_2_MPORT_390_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_392_en & pht_1_2_MPORT_392_mask) begin
      pht_1_2[pht_1_2_MPORT_392_addr] <= pht_1_2_MPORT_392_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_394_en & pht_1_2_MPORT_394_mask) begin
      pht_1_2[pht_1_2_MPORT_394_addr] <= pht_1_2_MPORT_394_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_396_en & pht_1_2_MPORT_396_mask) begin
      pht_1_2[pht_1_2_MPORT_396_addr] <= pht_1_2_MPORT_396_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_398_en & pht_1_2_MPORT_398_mask) begin
      pht_1_2[pht_1_2_MPORT_398_addr] <= pht_1_2_MPORT_398_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_400_en & pht_1_2_MPORT_400_mask) begin
      pht_1_2[pht_1_2_MPORT_400_addr] <= pht_1_2_MPORT_400_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_402_en & pht_1_2_MPORT_402_mask) begin
      pht_1_2[pht_1_2_MPORT_402_addr] <= pht_1_2_MPORT_402_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_404_en & pht_1_2_MPORT_404_mask) begin
      pht_1_2[pht_1_2_MPORT_404_addr] <= pht_1_2_MPORT_404_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_406_en & pht_1_2_MPORT_406_mask) begin
      pht_1_2[pht_1_2_MPORT_406_addr] <= pht_1_2_MPORT_406_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_408_en & pht_1_2_MPORT_408_mask) begin
      pht_1_2[pht_1_2_MPORT_408_addr] <= pht_1_2_MPORT_408_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_410_en & pht_1_2_MPORT_410_mask) begin
      pht_1_2[pht_1_2_MPORT_410_addr] <= pht_1_2_MPORT_410_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_412_en & pht_1_2_MPORT_412_mask) begin
      pht_1_2[pht_1_2_MPORT_412_addr] <= pht_1_2_MPORT_412_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_414_en & pht_1_2_MPORT_414_mask) begin
      pht_1_2[pht_1_2_MPORT_414_addr] <= pht_1_2_MPORT_414_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_416_en & pht_1_2_MPORT_416_mask) begin
      pht_1_2[pht_1_2_MPORT_416_addr] <= pht_1_2_MPORT_416_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_418_en & pht_1_2_MPORT_418_mask) begin
      pht_1_2[pht_1_2_MPORT_418_addr] <= pht_1_2_MPORT_418_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_420_en & pht_1_2_MPORT_420_mask) begin
      pht_1_2[pht_1_2_MPORT_420_addr] <= pht_1_2_MPORT_420_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_422_en & pht_1_2_MPORT_422_mask) begin
      pht_1_2[pht_1_2_MPORT_422_addr] <= pht_1_2_MPORT_422_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_424_en & pht_1_2_MPORT_424_mask) begin
      pht_1_2[pht_1_2_MPORT_424_addr] <= pht_1_2_MPORT_424_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_426_en & pht_1_2_MPORT_426_mask) begin
      pht_1_2[pht_1_2_MPORT_426_addr] <= pht_1_2_MPORT_426_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_428_en & pht_1_2_MPORT_428_mask) begin
      pht_1_2[pht_1_2_MPORT_428_addr] <= pht_1_2_MPORT_428_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_2_MPORT_430_en & pht_1_2_MPORT_430_mask) begin
      pht_1_2[pht_1_2_MPORT_430_addr] <= pht_1_2_MPORT_430_data; // @[PatternHistoryTable.scala 21:28]
    end
//     pht_1_2_MPORT_2_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_2_MPORT_2_addr_pipe_0 <= io_raddr_0;
    end
//     pht_1_2_MPORT_10_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_2_MPORT_10_addr_pipe_0 <= io_raddr_1;
    end
//     pht_1_2_MPORT_20_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_2_MPORT_20_addr_pipe_0 <= io_waddr;
    end
    if (pht_1_3_MPORT_38_en & pht_1_3_MPORT_38_mask) begin
      pht_1_3[pht_1_3_MPORT_38_addr] <= pht_1_3_MPORT_38_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_432_en & pht_1_3_MPORT_432_mask) begin
      pht_1_3[pht_1_3_MPORT_432_addr] <= pht_1_3_MPORT_432_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_434_en & pht_1_3_MPORT_434_mask) begin
      pht_1_3[pht_1_3_MPORT_434_addr] <= pht_1_3_MPORT_434_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_436_en & pht_1_3_MPORT_436_mask) begin
      pht_1_3[pht_1_3_MPORT_436_addr] <= pht_1_3_MPORT_436_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_438_en & pht_1_3_MPORT_438_mask) begin
      pht_1_3[pht_1_3_MPORT_438_addr] <= pht_1_3_MPORT_438_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_440_en & pht_1_3_MPORT_440_mask) begin
      pht_1_3[pht_1_3_MPORT_440_addr] <= pht_1_3_MPORT_440_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_442_en & pht_1_3_MPORT_442_mask) begin
      pht_1_3[pht_1_3_MPORT_442_addr] <= pht_1_3_MPORT_442_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_444_en & pht_1_3_MPORT_444_mask) begin
      pht_1_3[pht_1_3_MPORT_444_addr] <= pht_1_3_MPORT_444_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_446_en & pht_1_3_MPORT_446_mask) begin
      pht_1_3[pht_1_3_MPORT_446_addr] <= pht_1_3_MPORT_446_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_448_en & pht_1_3_MPORT_448_mask) begin
      pht_1_3[pht_1_3_MPORT_448_addr] <= pht_1_3_MPORT_448_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_450_en & pht_1_3_MPORT_450_mask) begin
      pht_1_3[pht_1_3_MPORT_450_addr] <= pht_1_3_MPORT_450_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_452_en & pht_1_3_MPORT_452_mask) begin
      pht_1_3[pht_1_3_MPORT_452_addr] <= pht_1_3_MPORT_452_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_454_en & pht_1_3_MPORT_454_mask) begin
      pht_1_3[pht_1_3_MPORT_454_addr] <= pht_1_3_MPORT_454_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_456_en & pht_1_3_MPORT_456_mask) begin
      pht_1_3[pht_1_3_MPORT_456_addr] <= pht_1_3_MPORT_456_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_458_en & pht_1_3_MPORT_458_mask) begin
      pht_1_3[pht_1_3_MPORT_458_addr] <= pht_1_3_MPORT_458_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_460_en & pht_1_3_MPORT_460_mask) begin
      pht_1_3[pht_1_3_MPORT_460_addr] <= pht_1_3_MPORT_460_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_462_en & pht_1_3_MPORT_462_mask) begin
      pht_1_3[pht_1_3_MPORT_462_addr] <= pht_1_3_MPORT_462_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_464_en & pht_1_3_MPORT_464_mask) begin
      pht_1_3[pht_1_3_MPORT_464_addr] <= pht_1_3_MPORT_464_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_466_en & pht_1_3_MPORT_466_mask) begin
      pht_1_3[pht_1_3_MPORT_466_addr] <= pht_1_3_MPORT_466_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_468_en & pht_1_3_MPORT_468_mask) begin
      pht_1_3[pht_1_3_MPORT_468_addr] <= pht_1_3_MPORT_468_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_470_en & pht_1_3_MPORT_470_mask) begin
      pht_1_3[pht_1_3_MPORT_470_addr] <= pht_1_3_MPORT_470_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_472_en & pht_1_3_MPORT_472_mask) begin
      pht_1_3[pht_1_3_MPORT_472_addr] <= pht_1_3_MPORT_472_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_474_en & pht_1_3_MPORT_474_mask) begin
      pht_1_3[pht_1_3_MPORT_474_addr] <= pht_1_3_MPORT_474_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_476_en & pht_1_3_MPORT_476_mask) begin
      pht_1_3[pht_1_3_MPORT_476_addr] <= pht_1_3_MPORT_476_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_478_en & pht_1_3_MPORT_478_mask) begin
      pht_1_3[pht_1_3_MPORT_478_addr] <= pht_1_3_MPORT_478_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_480_en & pht_1_3_MPORT_480_mask) begin
      pht_1_3[pht_1_3_MPORT_480_addr] <= pht_1_3_MPORT_480_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_482_en & pht_1_3_MPORT_482_mask) begin
      pht_1_3[pht_1_3_MPORT_482_addr] <= pht_1_3_MPORT_482_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_484_en & pht_1_3_MPORT_484_mask) begin
      pht_1_3[pht_1_3_MPORT_484_addr] <= pht_1_3_MPORT_484_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_486_en & pht_1_3_MPORT_486_mask) begin
      pht_1_3[pht_1_3_MPORT_486_addr] <= pht_1_3_MPORT_486_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_488_en & pht_1_3_MPORT_488_mask) begin
      pht_1_3[pht_1_3_MPORT_488_addr] <= pht_1_3_MPORT_488_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_490_en & pht_1_3_MPORT_490_mask) begin
      pht_1_3[pht_1_3_MPORT_490_addr] <= pht_1_3_MPORT_490_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_492_en & pht_1_3_MPORT_492_mask) begin
      pht_1_3[pht_1_3_MPORT_492_addr] <= pht_1_3_MPORT_492_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_494_en & pht_1_3_MPORT_494_mask) begin
      pht_1_3[pht_1_3_MPORT_494_addr] <= pht_1_3_MPORT_494_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_496_en & pht_1_3_MPORT_496_mask) begin
      pht_1_3[pht_1_3_MPORT_496_addr] <= pht_1_3_MPORT_496_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_498_en & pht_1_3_MPORT_498_mask) begin
      pht_1_3[pht_1_3_MPORT_498_addr] <= pht_1_3_MPORT_498_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_500_en & pht_1_3_MPORT_500_mask) begin
      pht_1_3[pht_1_3_MPORT_500_addr] <= pht_1_3_MPORT_500_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_502_en & pht_1_3_MPORT_502_mask) begin
      pht_1_3[pht_1_3_MPORT_502_addr] <= pht_1_3_MPORT_502_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_504_en & pht_1_3_MPORT_504_mask) begin
      pht_1_3[pht_1_3_MPORT_504_addr] <= pht_1_3_MPORT_504_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_506_en & pht_1_3_MPORT_506_mask) begin
      pht_1_3[pht_1_3_MPORT_506_addr] <= pht_1_3_MPORT_506_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_508_en & pht_1_3_MPORT_508_mask) begin
      pht_1_3[pht_1_3_MPORT_508_addr] <= pht_1_3_MPORT_508_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_510_en & pht_1_3_MPORT_510_mask) begin
      pht_1_3[pht_1_3_MPORT_510_addr] <= pht_1_3_MPORT_510_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_512_en & pht_1_3_MPORT_512_mask) begin
      pht_1_3[pht_1_3_MPORT_512_addr] <= pht_1_3_MPORT_512_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_514_en & pht_1_3_MPORT_514_mask) begin
      pht_1_3[pht_1_3_MPORT_514_addr] <= pht_1_3_MPORT_514_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_516_en & pht_1_3_MPORT_516_mask) begin
      pht_1_3[pht_1_3_MPORT_516_addr] <= pht_1_3_MPORT_516_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_518_en & pht_1_3_MPORT_518_mask) begin
      pht_1_3[pht_1_3_MPORT_518_addr] <= pht_1_3_MPORT_518_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_520_en & pht_1_3_MPORT_520_mask) begin
      pht_1_3[pht_1_3_MPORT_520_addr] <= pht_1_3_MPORT_520_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_522_en & pht_1_3_MPORT_522_mask) begin
      pht_1_3[pht_1_3_MPORT_522_addr] <= pht_1_3_MPORT_522_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_524_en & pht_1_3_MPORT_524_mask) begin
      pht_1_3[pht_1_3_MPORT_524_addr] <= pht_1_3_MPORT_524_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_526_en & pht_1_3_MPORT_526_mask) begin
      pht_1_3[pht_1_3_MPORT_526_addr] <= pht_1_3_MPORT_526_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_528_en & pht_1_3_MPORT_528_mask) begin
      pht_1_3[pht_1_3_MPORT_528_addr] <= pht_1_3_MPORT_528_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_530_en & pht_1_3_MPORT_530_mask) begin
      pht_1_3[pht_1_3_MPORT_530_addr] <= pht_1_3_MPORT_530_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_532_en & pht_1_3_MPORT_532_mask) begin
      pht_1_3[pht_1_3_MPORT_532_addr] <= pht_1_3_MPORT_532_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_534_en & pht_1_3_MPORT_534_mask) begin
      pht_1_3[pht_1_3_MPORT_534_addr] <= pht_1_3_MPORT_534_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_536_en & pht_1_3_MPORT_536_mask) begin
      pht_1_3[pht_1_3_MPORT_536_addr] <= pht_1_3_MPORT_536_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_538_en & pht_1_3_MPORT_538_mask) begin
      pht_1_3[pht_1_3_MPORT_538_addr] <= pht_1_3_MPORT_538_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_540_en & pht_1_3_MPORT_540_mask) begin
      pht_1_3[pht_1_3_MPORT_540_addr] <= pht_1_3_MPORT_540_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_542_en & pht_1_3_MPORT_542_mask) begin
      pht_1_3[pht_1_3_MPORT_542_addr] <= pht_1_3_MPORT_542_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_544_en & pht_1_3_MPORT_544_mask) begin
      pht_1_3[pht_1_3_MPORT_544_addr] <= pht_1_3_MPORT_544_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_546_en & pht_1_3_MPORT_546_mask) begin
      pht_1_3[pht_1_3_MPORT_546_addr] <= pht_1_3_MPORT_546_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_548_en & pht_1_3_MPORT_548_mask) begin
      pht_1_3[pht_1_3_MPORT_548_addr] <= pht_1_3_MPORT_548_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_550_en & pht_1_3_MPORT_550_mask) begin
      pht_1_3[pht_1_3_MPORT_550_addr] <= pht_1_3_MPORT_550_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_552_en & pht_1_3_MPORT_552_mask) begin
      pht_1_3[pht_1_3_MPORT_552_addr] <= pht_1_3_MPORT_552_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_554_en & pht_1_3_MPORT_554_mask) begin
      pht_1_3[pht_1_3_MPORT_554_addr] <= pht_1_3_MPORT_554_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_556_en & pht_1_3_MPORT_556_mask) begin
      pht_1_3[pht_1_3_MPORT_556_addr] <= pht_1_3_MPORT_556_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_3_MPORT_558_en & pht_1_3_MPORT_558_mask) begin
      pht_1_3[pht_1_3_MPORT_558_addr] <= pht_1_3_MPORT_558_data; // @[PatternHistoryTable.scala 21:28]
    end
//     pht_1_3_MPORT_3_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_3_MPORT_3_addr_pipe_0 <= io_raddr_0;
    end
//     pht_1_3_MPORT_11_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_3_MPORT_11_addr_pipe_0 <= io_raddr_1;
    end
//     pht_1_3_MPORT_22_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_3_MPORT_22_addr_pipe_0 <= io_waddr;
    end
    if (pht_1_4_MPORT_40_en & pht_1_4_MPORT_40_mask) begin
      pht_1_4[pht_1_4_MPORT_40_addr] <= pht_1_4_MPORT_40_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_560_en & pht_1_4_MPORT_560_mask) begin
      pht_1_4[pht_1_4_MPORT_560_addr] <= pht_1_4_MPORT_560_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_562_en & pht_1_4_MPORT_562_mask) begin
      pht_1_4[pht_1_4_MPORT_562_addr] <= pht_1_4_MPORT_562_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_564_en & pht_1_4_MPORT_564_mask) begin
      pht_1_4[pht_1_4_MPORT_564_addr] <= pht_1_4_MPORT_564_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_566_en & pht_1_4_MPORT_566_mask) begin
      pht_1_4[pht_1_4_MPORT_566_addr] <= pht_1_4_MPORT_566_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_568_en & pht_1_4_MPORT_568_mask) begin
      pht_1_4[pht_1_4_MPORT_568_addr] <= pht_1_4_MPORT_568_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_570_en & pht_1_4_MPORT_570_mask) begin
      pht_1_4[pht_1_4_MPORT_570_addr] <= pht_1_4_MPORT_570_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_572_en & pht_1_4_MPORT_572_mask) begin
      pht_1_4[pht_1_4_MPORT_572_addr] <= pht_1_4_MPORT_572_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_574_en & pht_1_4_MPORT_574_mask) begin
      pht_1_4[pht_1_4_MPORT_574_addr] <= pht_1_4_MPORT_574_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_576_en & pht_1_4_MPORT_576_mask) begin
      pht_1_4[pht_1_4_MPORT_576_addr] <= pht_1_4_MPORT_576_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_578_en & pht_1_4_MPORT_578_mask) begin
      pht_1_4[pht_1_4_MPORT_578_addr] <= pht_1_4_MPORT_578_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_580_en & pht_1_4_MPORT_580_mask) begin
      pht_1_4[pht_1_4_MPORT_580_addr] <= pht_1_4_MPORT_580_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_582_en & pht_1_4_MPORT_582_mask) begin
      pht_1_4[pht_1_4_MPORT_582_addr] <= pht_1_4_MPORT_582_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_584_en & pht_1_4_MPORT_584_mask) begin
      pht_1_4[pht_1_4_MPORT_584_addr] <= pht_1_4_MPORT_584_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_586_en & pht_1_4_MPORT_586_mask) begin
      pht_1_4[pht_1_4_MPORT_586_addr] <= pht_1_4_MPORT_586_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_588_en & pht_1_4_MPORT_588_mask) begin
      pht_1_4[pht_1_4_MPORT_588_addr] <= pht_1_4_MPORT_588_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_590_en & pht_1_4_MPORT_590_mask) begin
      pht_1_4[pht_1_4_MPORT_590_addr] <= pht_1_4_MPORT_590_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_592_en & pht_1_4_MPORT_592_mask) begin
      pht_1_4[pht_1_4_MPORT_592_addr] <= pht_1_4_MPORT_592_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_594_en & pht_1_4_MPORT_594_mask) begin
      pht_1_4[pht_1_4_MPORT_594_addr] <= pht_1_4_MPORT_594_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_596_en & pht_1_4_MPORT_596_mask) begin
      pht_1_4[pht_1_4_MPORT_596_addr] <= pht_1_4_MPORT_596_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_598_en & pht_1_4_MPORT_598_mask) begin
      pht_1_4[pht_1_4_MPORT_598_addr] <= pht_1_4_MPORT_598_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_600_en & pht_1_4_MPORT_600_mask) begin
      pht_1_4[pht_1_4_MPORT_600_addr] <= pht_1_4_MPORT_600_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_602_en & pht_1_4_MPORT_602_mask) begin
      pht_1_4[pht_1_4_MPORT_602_addr] <= pht_1_4_MPORT_602_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_604_en & pht_1_4_MPORT_604_mask) begin
      pht_1_4[pht_1_4_MPORT_604_addr] <= pht_1_4_MPORT_604_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_606_en & pht_1_4_MPORT_606_mask) begin
      pht_1_4[pht_1_4_MPORT_606_addr] <= pht_1_4_MPORT_606_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_608_en & pht_1_4_MPORT_608_mask) begin
      pht_1_4[pht_1_4_MPORT_608_addr] <= pht_1_4_MPORT_608_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_610_en & pht_1_4_MPORT_610_mask) begin
      pht_1_4[pht_1_4_MPORT_610_addr] <= pht_1_4_MPORT_610_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_612_en & pht_1_4_MPORT_612_mask) begin
      pht_1_4[pht_1_4_MPORT_612_addr] <= pht_1_4_MPORT_612_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_614_en & pht_1_4_MPORT_614_mask) begin
      pht_1_4[pht_1_4_MPORT_614_addr] <= pht_1_4_MPORT_614_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_616_en & pht_1_4_MPORT_616_mask) begin
      pht_1_4[pht_1_4_MPORT_616_addr] <= pht_1_4_MPORT_616_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_618_en & pht_1_4_MPORT_618_mask) begin
      pht_1_4[pht_1_4_MPORT_618_addr] <= pht_1_4_MPORT_618_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_620_en & pht_1_4_MPORT_620_mask) begin
      pht_1_4[pht_1_4_MPORT_620_addr] <= pht_1_4_MPORT_620_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_622_en & pht_1_4_MPORT_622_mask) begin
      pht_1_4[pht_1_4_MPORT_622_addr] <= pht_1_4_MPORT_622_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_624_en & pht_1_4_MPORT_624_mask) begin
      pht_1_4[pht_1_4_MPORT_624_addr] <= pht_1_4_MPORT_624_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_626_en & pht_1_4_MPORT_626_mask) begin
      pht_1_4[pht_1_4_MPORT_626_addr] <= pht_1_4_MPORT_626_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_628_en & pht_1_4_MPORT_628_mask) begin
      pht_1_4[pht_1_4_MPORT_628_addr] <= pht_1_4_MPORT_628_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_630_en & pht_1_4_MPORT_630_mask) begin
      pht_1_4[pht_1_4_MPORT_630_addr] <= pht_1_4_MPORT_630_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_632_en & pht_1_4_MPORT_632_mask) begin
      pht_1_4[pht_1_4_MPORT_632_addr] <= pht_1_4_MPORT_632_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_634_en & pht_1_4_MPORT_634_mask) begin
      pht_1_4[pht_1_4_MPORT_634_addr] <= pht_1_4_MPORT_634_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_636_en & pht_1_4_MPORT_636_mask) begin
      pht_1_4[pht_1_4_MPORT_636_addr] <= pht_1_4_MPORT_636_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_638_en & pht_1_4_MPORT_638_mask) begin
      pht_1_4[pht_1_4_MPORT_638_addr] <= pht_1_4_MPORT_638_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_640_en & pht_1_4_MPORT_640_mask) begin
      pht_1_4[pht_1_4_MPORT_640_addr] <= pht_1_4_MPORT_640_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_642_en & pht_1_4_MPORT_642_mask) begin
      pht_1_4[pht_1_4_MPORT_642_addr] <= pht_1_4_MPORT_642_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_644_en & pht_1_4_MPORT_644_mask) begin
      pht_1_4[pht_1_4_MPORT_644_addr] <= pht_1_4_MPORT_644_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_646_en & pht_1_4_MPORT_646_mask) begin
      pht_1_4[pht_1_4_MPORT_646_addr] <= pht_1_4_MPORT_646_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_648_en & pht_1_4_MPORT_648_mask) begin
      pht_1_4[pht_1_4_MPORT_648_addr] <= pht_1_4_MPORT_648_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_650_en & pht_1_4_MPORT_650_mask) begin
      pht_1_4[pht_1_4_MPORT_650_addr] <= pht_1_4_MPORT_650_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_652_en & pht_1_4_MPORT_652_mask) begin
      pht_1_4[pht_1_4_MPORT_652_addr] <= pht_1_4_MPORT_652_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_654_en & pht_1_4_MPORT_654_mask) begin
      pht_1_4[pht_1_4_MPORT_654_addr] <= pht_1_4_MPORT_654_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_656_en & pht_1_4_MPORT_656_mask) begin
      pht_1_4[pht_1_4_MPORT_656_addr] <= pht_1_4_MPORT_656_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_658_en & pht_1_4_MPORT_658_mask) begin
      pht_1_4[pht_1_4_MPORT_658_addr] <= pht_1_4_MPORT_658_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_660_en & pht_1_4_MPORT_660_mask) begin
      pht_1_4[pht_1_4_MPORT_660_addr] <= pht_1_4_MPORT_660_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_662_en & pht_1_4_MPORT_662_mask) begin
      pht_1_4[pht_1_4_MPORT_662_addr] <= pht_1_4_MPORT_662_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_664_en & pht_1_4_MPORT_664_mask) begin
      pht_1_4[pht_1_4_MPORT_664_addr] <= pht_1_4_MPORT_664_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_666_en & pht_1_4_MPORT_666_mask) begin
      pht_1_4[pht_1_4_MPORT_666_addr] <= pht_1_4_MPORT_666_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_668_en & pht_1_4_MPORT_668_mask) begin
      pht_1_4[pht_1_4_MPORT_668_addr] <= pht_1_4_MPORT_668_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_670_en & pht_1_4_MPORT_670_mask) begin
      pht_1_4[pht_1_4_MPORT_670_addr] <= pht_1_4_MPORT_670_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_672_en & pht_1_4_MPORT_672_mask) begin
      pht_1_4[pht_1_4_MPORT_672_addr] <= pht_1_4_MPORT_672_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_674_en & pht_1_4_MPORT_674_mask) begin
      pht_1_4[pht_1_4_MPORT_674_addr] <= pht_1_4_MPORT_674_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_676_en & pht_1_4_MPORT_676_mask) begin
      pht_1_4[pht_1_4_MPORT_676_addr] <= pht_1_4_MPORT_676_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_678_en & pht_1_4_MPORT_678_mask) begin
      pht_1_4[pht_1_4_MPORT_678_addr] <= pht_1_4_MPORT_678_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_680_en & pht_1_4_MPORT_680_mask) begin
      pht_1_4[pht_1_4_MPORT_680_addr] <= pht_1_4_MPORT_680_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_682_en & pht_1_4_MPORT_682_mask) begin
      pht_1_4[pht_1_4_MPORT_682_addr] <= pht_1_4_MPORT_682_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_684_en & pht_1_4_MPORT_684_mask) begin
      pht_1_4[pht_1_4_MPORT_684_addr] <= pht_1_4_MPORT_684_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_4_MPORT_686_en & pht_1_4_MPORT_686_mask) begin
      pht_1_4[pht_1_4_MPORT_686_addr] <= pht_1_4_MPORT_686_data; // @[PatternHistoryTable.scala 21:28]
    end
//     pht_1_4_MPORT_4_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_4_MPORT_4_addr_pipe_0 <= io_raddr_0;
    end
//     pht_1_4_MPORT_12_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_4_MPORT_12_addr_pipe_0 <= io_raddr_1;
    end
//     pht_1_4_MPORT_24_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_4_MPORT_24_addr_pipe_0 <= io_waddr;
    end
    if (pht_1_5_MPORT_42_en & pht_1_5_MPORT_42_mask) begin
      pht_1_5[pht_1_5_MPORT_42_addr] <= pht_1_5_MPORT_42_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_688_en & pht_1_5_MPORT_688_mask) begin
      pht_1_5[pht_1_5_MPORT_688_addr] <= pht_1_5_MPORT_688_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_690_en & pht_1_5_MPORT_690_mask) begin
      pht_1_5[pht_1_5_MPORT_690_addr] <= pht_1_5_MPORT_690_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_692_en & pht_1_5_MPORT_692_mask) begin
      pht_1_5[pht_1_5_MPORT_692_addr] <= pht_1_5_MPORT_692_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_694_en & pht_1_5_MPORT_694_mask) begin
      pht_1_5[pht_1_5_MPORT_694_addr] <= pht_1_5_MPORT_694_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_696_en & pht_1_5_MPORT_696_mask) begin
      pht_1_5[pht_1_5_MPORT_696_addr] <= pht_1_5_MPORT_696_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_698_en & pht_1_5_MPORT_698_mask) begin
      pht_1_5[pht_1_5_MPORT_698_addr] <= pht_1_5_MPORT_698_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_700_en & pht_1_5_MPORT_700_mask) begin
      pht_1_5[pht_1_5_MPORT_700_addr] <= pht_1_5_MPORT_700_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_702_en & pht_1_5_MPORT_702_mask) begin
      pht_1_5[pht_1_5_MPORT_702_addr] <= pht_1_5_MPORT_702_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_704_en & pht_1_5_MPORT_704_mask) begin
      pht_1_5[pht_1_5_MPORT_704_addr] <= pht_1_5_MPORT_704_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_706_en & pht_1_5_MPORT_706_mask) begin
      pht_1_5[pht_1_5_MPORT_706_addr] <= pht_1_5_MPORT_706_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_708_en & pht_1_5_MPORT_708_mask) begin
      pht_1_5[pht_1_5_MPORT_708_addr] <= pht_1_5_MPORT_708_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_710_en & pht_1_5_MPORT_710_mask) begin
      pht_1_5[pht_1_5_MPORT_710_addr] <= pht_1_5_MPORT_710_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_712_en & pht_1_5_MPORT_712_mask) begin
      pht_1_5[pht_1_5_MPORT_712_addr] <= pht_1_5_MPORT_712_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_714_en & pht_1_5_MPORT_714_mask) begin
      pht_1_5[pht_1_5_MPORT_714_addr] <= pht_1_5_MPORT_714_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_716_en & pht_1_5_MPORT_716_mask) begin
      pht_1_5[pht_1_5_MPORT_716_addr] <= pht_1_5_MPORT_716_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_718_en & pht_1_5_MPORT_718_mask) begin
      pht_1_5[pht_1_5_MPORT_718_addr] <= pht_1_5_MPORT_718_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_720_en & pht_1_5_MPORT_720_mask) begin
      pht_1_5[pht_1_5_MPORT_720_addr] <= pht_1_5_MPORT_720_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_722_en & pht_1_5_MPORT_722_mask) begin
      pht_1_5[pht_1_5_MPORT_722_addr] <= pht_1_5_MPORT_722_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_724_en & pht_1_5_MPORT_724_mask) begin
      pht_1_5[pht_1_5_MPORT_724_addr] <= pht_1_5_MPORT_724_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_726_en & pht_1_5_MPORT_726_mask) begin
      pht_1_5[pht_1_5_MPORT_726_addr] <= pht_1_5_MPORT_726_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_728_en & pht_1_5_MPORT_728_mask) begin
      pht_1_5[pht_1_5_MPORT_728_addr] <= pht_1_5_MPORT_728_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_730_en & pht_1_5_MPORT_730_mask) begin
      pht_1_5[pht_1_5_MPORT_730_addr] <= pht_1_5_MPORT_730_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_732_en & pht_1_5_MPORT_732_mask) begin
      pht_1_5[pht_1_5_MPORT_732_addr] <= pht_1_5_MPORT_732_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_734_en & pht_1_5_MPORT_734_mask) begin
      pht_1_5[pht_1_5_MPORT_734_addr] <= pht_1_5_MPORT_734_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_736_en & pht_1_5_MPORT_736_mask) begin
      pht_1_5[pht_1_5_MPORT_736_addr] <= pht_1_5_MPORT_736_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_738_en & pht_1_5_MPORT_738_mask) begin
      pht_1_5[pht_1_5_MPORT_738_addr] <= pht_1_5_MPORT_738_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_740_en & pht_1_5_MPORT_740_mask) begin
      pht_1_5[pht_1_5_MPORT_740_addr] <= pht_1_5_MPORT_740_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_742_en & pht_1_5_MPORT_742_mask) begin
      pht_1_5[pht_1_5_MPORT_742_addr] <= pht_1_5_MPORT_742_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_744_en & pht_1_5_MPORT_744_mask) begin
      pht_1_5[pht_1_5_MPORT_744_addr] <= pht_1_5_MPORT_744_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_746_en & pht_1_5_MPORT_746_mask) begin
      pht_1_5[pht_1_5_MPORT_746_addr] <= pht_1_5_MPORT_746_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_748_en & pht_1_5_MPORT_748_mask) begin
      pht_1_5[pht_1_5_MPORT_748_addr] <= pht_1_5_MPORT_748_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_750_en & pht_1_5_MPORT_750_mask) begin
      pht_1_5[pht_1_5_MPORT_750_addr] <= pht_1_5_MPORT_750_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_752_en & pht_1_5_MPORT_752_mask) begin
      pht_1_5[pht_1_5_MPORT_752_addr] <= pht_1_5_MPORT_752_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_754_en & pht_1_5_MPORT_754_mask) begin
      pht_1_5[pht_1_5_MPORT_754_addr] <= pht_1_5_MPORT_754_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_756_en & pht_1_5_MPORT_756_mask) begin
      pht_1_5[pht_1_5_MPORT_756_addr] <= pht_1_5_MPORT_756_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_758_en & pht_1_5_MPORT_758_mask) begin
      pht_1_5[pht_1_5_MPORT_758_addr] <= pht_1_5_MPORT_758_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_760_en & pht_1_5_MPORT_760_mask) begin
      pht_1_5[pht_1_5_MPORT_760_addr] <= pht_1_5_MPORT_760_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_762_en & pht_1_5_MPORT_762_mask) begin
      pht_1_5[pht_1_5_MPORT_762_addr] <= pht_1_5_MPORT_762_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_764_en & pht_1_5_MPORT_764_mask) begin
      pht_1_5[pht_1_5_MPORT_764_addr] <= pht_1_5_MPORT_764_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_766_en & pht_1_5_MPORT_766_mask) begin
      pht_1_5[pht_1_5_MPORT_766_addr] <= pht_1_5_MPORT_766_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_768_en & pht_1_5_MPORT_768_mask) begin
      pht_1_5[pht_1_5_MPORT_768_addr] <= pht_1_5_MPORT_768_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_770_en & pht_1_5_MPORT_770_mask) begin
      pht_1_5[pht_1_5_MPORT_770_addr] <= pht_1_5_MPORT_770_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_772_en & pht_1_5_MPORT_772_mask) begin
      pht_1_5[pht_1_5_MPORT_772_addr] <= pht_1_5_MPORT_772_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_774_en & pht_1_5_MPORT_774_mask) begin
      pht_1_5[pht_1_5_MPORT_774_addr] <= pht_1_5_MPORT_774_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_776_en & pht_1_5_MPORT_776_mask) begin
      pht_1_5[pht_1_5_MPORT_776_addr] <= pht_1_5_MPORT_776_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_778_en & pht_1_5_MPORT_778_mask) begin
      pht_1_5[pht_1_5_MPORT_778_addr] <= pht_1_5_MPORT_778_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_780_en & pht_1_5_MPORT_780_mask) begin
      pht_1_5[pht_1_5_MPORT_780_addr] <= pht_1_5_MPORT_780_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_782_en & pht_1_5_MPORT_782_mask) begin
      pht_1_5[pht_1_5_MPORT_782_addr] <= pht_1_5_MPORT_782_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_784_en & pht_1_5_MPORT_784_mask) begin
      pht_1_5[pht_1_5_MPORT_784_addr] <= pht_1_5_MPORT_784_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_786_en & pht_1_5_MPORT_786_mask) begin
      pht_1_5[pht_1_5_MPORT_786_addr] <= pht_1_5_MPORT_786_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_788_en & pht_1_5_MPORT_788_mask) begin
      pht_1_5[pht_1_5_MPORT_788_addr] <= pht_1_5_MPORT_788_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_790_en & pht_1_5_MPORT_790_mask) begin
      pht_1_5[pht_1_5_MPORT_790_addr] <= pht_1_5_MPORT_790_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_792_en & pht_1_5_MPORT_792_mask) begin
      pht_1_5[pht_1_5_MPORT_792_addr] <= pht_1_5_MPORT_792_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_794_en & pht_1_5_MPORT_794_mask) begin
      pht_1_5[pht_1_5_MPORT_794_addr] <= pht_1_5_MPORT_794_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_796_en & pht_1_5_MPORT_796_mask) begin
      pht_1_5[pht_1_5_MPORT_796_addr] <= pht_1_5_MPORT_796_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_798_en & pht_1_5_MPORT_798_mask) begin
      pht_1_5[pht_1_5_MPORT_798_addr] <= pht_1_5_MPORT_798_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_800_en & pht_1_5_MPORT_800_mask) begin
      pht_1_5[pht_1_5_MPORT_800_addr] <= pht_1_5_MPORT_800_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_802_en & pht_1_5_MPORT_802_mask) begin
      pht_1_5[pht_1_5_MPORT_802_addr] <= pht_1_5_MPORT_802_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_804_en & pht_1_5_MPORT_804_mask) begin
      pht_1_5[pht_1_5_MPORT_804_addr] <= pht_1_5_MPORT_804_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_806_en & pht_1_5_MPORT_806_mask) begin
      pht_1_5[pht_1_5_MPORT_806_addr] <= pht_1_5_MPORT_806_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_808_en & pht_1_5_MPORT_808_mask) begin
      pht_1_5[pht_1_5_MPORT_808_addr] <= pht_1_5_MPORT_808_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_810_en & pht_1_5_MPORT_810_mask) begin
      pht_1_5[pht_1_5_MPORT_810_addr] <= pht_1_5_MPORT_810_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_812_en & pht_1_5_MPORT_812_mask) begin
      pht_1_5[pht_1_5_MPORT_812_addr] <= pht_1_5_MPORT_812_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_5_MPORT_814_en & pht_1_5_MPORT_814_mask) begin
      pht_1_5[pht_1_5_MPORT_814_addr] <= pht_1_5_MPORT_814_data; // @[PatternHistoryTable.scala 21:28]
    end
//     pht_1_5_MPORT_5_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_5_MPORT_5_addr_pipe_0 <= io_raddr_0;
    end
//     pht_1_5_MPORT_13_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_5_MPORT_13_addr_pipe_0 <= io_raddr_1;
    end
//     pht_1_5_MPORT_26_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_5_MPORT_26_addr_pipe_0 <= io_waddr;
    end
    if (pht_1_6_MPORT_44_en & pht_1_6_MPORT_44_mask) begin
      pht_1_6[pht_1_6_MPORT_44_addr] <= pht_1_6_MPORT_44_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_816_en & pht_1_6_MPORT_816_mask) begin
      pht_1_6[pht_1_6_MPORT_816_addr] <= pht_1_6_MPORT_816_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_818_en & pht_1_6_MPORT_818_mask) begin
      pht_1_6[pht_1_6_MPORT_818_addr] <= pht_1_6_MPORT_818_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_820_en & pht_1_6_MPORT_820_mask) begin
      pht_1_6[pht_1_6_MPORT_820_addr] <= pht_1_6_MPORT_820_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_822_en & pht_1_6_MPORT_822_mask) begin
      pht_1_6[pht_1_6_MPORT_822_addr] <= pht_1_6_MPORT_822_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_824_en & pht_1_6_MPORT_824_mask) begin
      pht_1_6[pht_1_6_MPORT_824_addr] <= pht_1_6_MPORT_824_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_826_en & pht_1_6_MPORT_826_mask) begin
      pht_1_6[pht_1_6_MPORT_826_addr] <= pht_1_6_MPORT_826_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_828_en & pht_1_6_MPORT_828_mask) begin
      pht_1_6[pht_1_6_MPORT_828_addr] <= pht_1_6_MPORT_828_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_830_en & pht_1_6_MPORT_830_mask) begin
      pht_1_6[pht_1_6_MPORT_830_addr] <= pht_1_6_MPORT_830_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_832_en & pht_1_6_MPORT_832_mask) begin
      pht_1_6[pht_1_6_MPORT_832_addr] <= pht_1_6_MPORT_832_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_834_en & pht_1_6_MPORT_834_mask) begin
      pht_1_6[pht_1_6_MPORT_834_addr] <= pht_1_6_MPORT_834_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_836_en & pht_1_6_MPORT_836_mask) begin
      pht_1_6[pht_1_6_MPORT_836_addr] <= pht_1_6_MPORT_836_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_838_en & pht_1_6_MPORT_838_mask) begin
      pht_1_6[pht_1_6_MPORT_838_addr] <= pht_1_6_MPORT_838_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_840_en & pht_1_6_MPORT_840_mask) begin
      pht_1_6[pht_1_6_MPORT_840_addr] <= pht_1_6_MPORT_840_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_842_en & pht_1_6_MPORT_842_mask) begin
      pht_1_6[pht_1_6_MPORT_842_addr] <= pht_1_6_MPORT_842_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_844_en & pht_1_6_MPORT_844_mask) begin
      pht_1_6[pht_1_6_MPORT_844_addr] <= pht_1_6_MPORT_844_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_846_en & pht_1_6_MPORT_846_mask) begin
      pht_1_6[pht_1_6_MPORT_846_addr] <= pht_1_6_MPORT_846_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_848_en & pht_1_6_MPORT_848_mask) begin
      pht_1_6[pht_1_6_MPORT_848_addr] <= pht_1_6_MPORT_848_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_850_en & pht_1_6_MPORT_850_mask) begin
      pht_1_6[pht_1_6_MPORT_850_addr] <= pht_1_6_MPORT_850_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_852_en & pht_1_6_MPORT_852_mask) begin
      pht_1_6[pht_1_6_MPORT_852_addr] <= pht_1_6_MPORT_852_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_854_en & pht_1_6_MPORT_854_mask) begin
      pht_1_6[pht_1_6_MPORT_854_addr] <= pht_1_6_MPORT_854_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_856_en & pht_1_6_MPORT_856_mask) begin
      pht_1_6[pht_1_6_MPORT_856_addr] <= pht_1_6_MPORT_856_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_858_en & pht_1_6_MPORT_858_mask) begin
      pht_1_6[pht_1_6_MPORT_858_addr] <= pht_1_6_MPORT_858_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_860_en & pht_1_6_MPORT_860_mask) begin
      pht_1_6[pht_1_6_MPORT_860_addr] <= pht_1_6_MPORT_860_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_862_en & pht_1_6_MPORT_862_mask) begin
      pht_1_6[pht_1_6_MPORT_862_addr] <= pht_1_6_MPORT_862_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_864_en & pht_1_6_MPORT_864_mask) begin
      pht_1_6[pht_1_6_MPORT_864_addr] <= pht_1_6_MPORT_864_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_866_en & pht_1_6_MPORT_866_mask) begin
      pht_1_6[pht_1_6_MPORT_866_addr] <= pht_1_6_MPORT_866_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_868_en & pht_1_6_MPORT_868_mask) begin
      pht_1_6[pht_1_6_MPORT_868_addr] <= pht_1_6_MPORT_868_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_870_en & pht_1_6_MPORT_870_mask) begin
      pht_1_6[pht_1_6_MPORT_870_addr] <= pht_1_6_MPORT_870_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_872_en & pht_1_6_MPORT_872_mask) begin
      pht_1_6[pht_1_6_MPORT_872_addr] <= pht_1_6_MPORT_872_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_874_en & pht_1_6_MPORT_874_mask) begin
      pht_1_6[pht_1_6_MPORT_874_addr] <= pht_1_6_MPORT_874_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_876_en & pht_1_6_MPORT_876_mask) begin
      pht_1_6[pht_1_6_MPORT_876_addr] <= pht_1_6_MPORT_876_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_878_en & pht_1_6_MPORT_878_mask) begin
      pht_1_6[pht_1_6_MPORT_878_addr] <= pht_1_6_MPORT_878_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_880_en & pht_1_6_MPORT_880_mask) begin
      pht_1_6[pht_1_6_MPORT_880_addr] <= pht_1_6_MPORT_880_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_882_en & pht_1_6_MPORT_882_mask) begin
      pht_1_6[pht_1_6_MPORT_882_addr] <= pht_1_6_MPORT_882_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_884_en & pht_1_6_MPORT_884_mask) begin
      pht_1_6[pht_1_6_MPORT_884_addr] <= pht_1_6_MPORT_884_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_886_en & pht_1_6_MPORT_886_mask) begin
      pht_1_6[pht_1_6_MPORT_886_addr] <= pht_1_6_MPORT_886_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_888_en & pht_1_6_MPORT_888_mask) begin
      pht_1_6[pht_1_6_MPORT_888_addr] <= pht_1_6_MPORT_888_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_890_en & pht_1_6_MPORT_890_mask) begin
      pht_1_6[pht_1_6_MPORT_890_addr] <= pht_1_6_MPORT_890_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_892_en & pht_1_6_MPORT_892_mask) begin
      pht_1_6[pht_1_6_MPORT_892_addr] <= pht_1_6_MPORT_892_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_894_en & pht_1_6_MPORT_894_mask) begin
      pht_1_6[pht_1_6_MPORT_894_addr] <= pht_1_6_MPORT_894_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_896_en & pht_1_6_MPORT_896_mask) begin
      pht_1_6[pht_1_6_MPORT_896_addr] <= pht_1_6_MPORT_896_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_898_en & pht_1_6_MPORT_898_mask) begin
      pht_1_6[pht_1_6_MPORT_898_addr] <= pht_1_6_MPORT_898_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_900_en & pht_1_6_MPORT_900_mask) begin
      pht_1_6[pht_1_6_MPORT_900_addr] <= pht_1_6_MPORT_900_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_902_en & pht_1_6_MPORT_902_mask) begin
      pht_1_6[pht_1_6_MPORT_902_addr] <= pht_1_6_MPORT_902_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_904_en & pht_1_6_MPORT_904_mask) begin
      pht_1_6[pht_1_6_MPORT_904_addr] <= pht_1_6_MPORT_904_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_906_en & pht_1_6_MPORT_906_mask) begin
      pht_1_6[pht_1_6_MPORT_906_addr] <= pht_1_6_MPORT_906_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_908_en & pht_1_6_MPORT_908_mask) begin
      pht_1_6[pht_1_6_MPORT_908_addr] <= pht_1_6_MPORT_908_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_910_en & pht_1_6_MPORT_910_mask) begin
      pht_1_6[pht_1_6_MPORT_910_addr] <= pht_1_6_MPORT_910_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_912_en & pht_1_6_MPORT_912_mask) begin
      pht_1_6[pht_1_6_MPORT_912_addr] <= pht_1_6_MPORT_912_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_914_en & pht_1_6_MPORT_914_mask) begin
      pht_1_6[pht_1_6_MPORT_914_addr] <= pht_1_6_MPORT_914_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_916_en & pht_1_6_MPORT_916_mask) begin
      pht_1_6[pht_1_6_MPORT_916_addr] <= pht_1_6_MPORT_916_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_918_en & pht_1_6_MPORT_918_mask) begin
      pht_1_6[pht_1_6_MPORT_918_addr] <= pht_1_6_MPORT_918_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_920_en & pht_1_6_MPORT_920_mask) begin
      pht_1_6[pht_1_6_MPORT_920_addr] <= pht_1_6_MPORT_920_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_922_en & pht_1_6_MPORT_922_mask) begin
      pht_1_6[pht_1_6_MPORT_922_addr] <= pht_1_6_MPORT_922_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_924_en & pht_1_6_MPORT_924_mask) begin
      pht_1_6[pht_1_6_MPORT_924_addr] <= pht_1_6_MPORT_924_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_926_en & pht_1_6_MPORT_926_mask) begin
      pht_1_6[pht_1_6_MPORT_926_addr] <= pht_1_6_MPORT_926_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_928_en & pht_1_6_MPORT_928_mask) begin
      pht_1_6[pht_1_6_MPORT_928_addr] <= pht_1_6_MPORT_928_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_930_en & pht_1_6_MPORT_930_mask) begin
      pht_1_6[pht_1_6_MPORT_930_addr] <= pht_1_6_MPORT_930_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_932_en & pht_1_6_MPORT_932_mask) begin
      pht_1_6[pht_1_6_MPORT_932_addr] <= pht_1_6_MPORT_932_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_934_en & pht_1_6_MPORT_934_mask) begin
      pht_1_6[pht_1_6_MPORT_934_addr] <= pht_1_6_MPORT_934_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_936_en & pht_1_6_MPORT_936_mask) begin
      pht_1_6[pht_1_6_MPORT_936_addr] <= pht_1_6_MPORT_936_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_938_en & pht_1_6_MPORT_938_mask) begin
      pht_1_6[pht_1_6_MPORT_938_addr] <= pht_1_6_MPORT_938_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_940_en & pht_1_6_MPORT_940_mask) begin
      pht_1_6[pht_1_6_MPORT_940_addr] <= pht_1_6_MPORT_940_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_6_MPORT_942_en & pht_1_6_MPORT_942_mask) begin
      pht_1_6[pht_1_6_MPORT_942_addr] <= pht_1_6_MPORT_942_data; // @[PatternHistoryTable.scala 21:28]
    end
//     pht_1_6_MPORT_6_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_6_MPORT_6_addr_pipe_0 <= io_raddr_0;
    end
//     pht_1_6_MPORT_14_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_6_MPORT_14_addr_pipe_0 <= io_raddr_1;
    end
//     pht_1_6_MPORT_28_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_6_MPORT_28_addr_pipe_0 <= io_waddr;
    end
    if (pht_1_7_MPORT_46_en & pht_1_7_MPORT_46_mask) begin
      pht_1_7[pht_1_7_MPORT_46_addr] <= pht_1_7_MPORT_46_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_944_en & pht_1_7_MPORT_944_mask) begin
      pht_1_7[pht_1_7_MPORT_944_addr] <= pht_1_7_MPORT_944_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_946_en & pht_1_7_MPORT_946_mask) begin
      pht_1_7[pht_1_7_MPORT_946_addr] <= pht_1_7_MPORT_946_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_948_en & pht_1_7_MPORT_948_mask) begin
      pht_1_7[pht_1_7_MPORT_948_addr] <= pht_1_7_MPORT_948_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_950_en & pht_1_7_MPORT_950_mask) begin
      pht_1_7[pht_1_7_MPORT_950_addr] <= pht_1_7_MPORT_950_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_952_en & pht_1_7_MPORT_952_mask) begin
      pht_1_7[pht_1_7_MPORT_952_addr] <= pht_1_7_MPORT_952_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_954_en & pht_1_7_MPORT_954_mask) begin
      pht_1_7[pht_1_7_MPORT_954_addr] <= pht_1_7_MPORT_954_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_956_en & pht_1_7_MPORT_956_mask) begin
      pht_1_7[pht_1_7_MPORT_956_addr] <= pht_1_7_MPORT_956_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_958_en & pht_1_7_MPORT_958_mask) begin
      pht_1_7[pht_1_7_MPORT_958_addr] <= pht_1_7_MPORT_958_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_960_en & pht_1_7_MPORT_960_mask) begin
      pht_1_7[pht_1_7_MPORT_960_addr] <= pht_1_7_MPORT_960_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_962_en & pht_1_7_MPORT_962_mask) begin
      pht_1_7[pht_1_7_MPORT_962_addr] <= pht_1_7_MPORT_962_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_964_en & pht_1_7_MPORT_964_mask) begin
      pht_1_7[pht_1_7_MPORT_964_addr] <= pht_1_7_MPORT_964_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_966_en & pht_1_7_MPORT_966_mask) begin
      pht_1_7[pht_1_7_MPORT_966_addr] <= pht_1_7_MPORT_966_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_968_en & pht_1_7_MPORT_968_mask) begin
      pht_1_7[pht_1_7_MPORT_968_addr] <= pht_1_7_MPORT_968_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_970_en & pht_1_7_MPORT_970_mask) begin
      pht_1_7[pht_1_7_MPORT_970_addr] <= pht_1_7_MPORT_970_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_972_en & pht_1_7_MPORT_972_mask) begin
      pht_1_7[pht_1_7_MPORT_972_addr] <= pht_1_7_MPORT_972_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_974_en & pht_1_7_MPORT_974_mask) begin
      pht_1_7[pht_1_7_MPORT_974_addr] <= pht_1_7_MPORT_974_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_976_en & pht_1_7_MPORT_976_mask) begin
      pht_1_7[pht_1_7_MPORT_976_addr] <= pht_1_7_MPORT_976_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_978_en & pht_1_7_MPORT_978_mask) begin
      pht_1_7[pht_1_7_MPORT_978_addr] <= pht_1_7_MPORT_978_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_980_en & pht_1_7_MPORT_980_mask) begin
      pht_1_7[pht_1_7_MPORT_980_addr] <= pht_1_7_MPORT_980_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_982_en & pht_1_7_MPORT_982_mask) begin
      pht_1_7[pht_1_7_MPORT_982_addr] <= pht_1_7_MPORT_982_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_984_en & pht_1_7_MPORT_984_mask) begin
      pht_1_7[pht_1_7_MPORT_984_addr] <= pht_1_7_MPORT_984_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_986_en & pht_1_7_MPORT_986_mask) begin
      pht_1_7[pht_1_7_MPORT_986_addr] <= pht_1_7_MPORT_986_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_988_en & pht_1_7_MPORT_988_mask) begin
      pht_1_7[pht_1_7_MPORT_988_addr] <= pht_1_7_MPORT_988_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_990_en & pht_1_7_MPORT_990_mask) begin
      pht_1_7[pht_1_7_MPORT_990_addr] <= pht_1_7_MPORT_990_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_992_en & pht_1_7_MPORT_992_mask) begin
      pht_1_7[pht_1_7_MPORT_992_addr] <= pht_1_7_MPORT_992_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_994_en & pht_1_7_MPORT_994_mask) begin
      pht_1_7[pht_1_7_MPORT_994_addr] <= pht_1_7_MPORT_994_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_996_en & pht_1_7_MPORT_996_mask) begin
      pht_1_7[pht_1_7_MPORT_996_addr] <= pht_1_7_MPORT_996_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_998_en & pht_1_7_MPORT_998_mask) begin
      pht_1_7[pht_1_7_MPORT_998_addr] <= pht_1_7_MPORT_998_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1000_en & pht_1_7_MPORT_1000_mask) begin
      pht_1_7[pht_1_7_MPORT_1000_addr] <= pht_1_7_MPORT_1000_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1002_en & pht_1_7_MPORT_1002_mask) begin
      pht_1_7[pht_1_7_MPORT_1002_addr] <= pht_1_7_MPORT_1002_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1004_en & pht_1_7_MPORT_1004_mask) begin
      pht_1_7[pht_1_7_MPORT_1004_addr] <= pht_1_7_MPORT_1004_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1006_en & pht_1_7_MPORT_1006_mask) begin
      pht_1_7[pht_1_7_MPORT_1006_addr] <= pht_1_7_MPORT_1006_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1008_en & pht_1_7_MPORT_1008_mask) begin
      pht_1_7[pht_1_7_MPORT_1008_addr] <= pht_1_7_MPORT_1008_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1010_en & pht_1_7_MPORT_1010_mask) begin
      pht_1_7[pht_1_7_MPORT_1010_addr] <= pht_1_7_MPORT_1010_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1012_en & pht_1_7_MPORT_1012_mask) begin
      pht_1_7[pht_1_7_MPORT_1012_addr] <= pht_1_7_MPORT_1012_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1014_en & pht_1_7_MPORT_1014_mask) begin
      pht_1_7[pht_1_7_MPORT_1014_addr] <= pht_1_7_MPORT_1014_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1016_en & pht_1_7_MPORT_1016_mask) begin
      pht_1_7[pht_1_7_MPORT_1016_addr] <= pht_1_7_MPORT_1016_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1018_en & pht_1_7_MPORT_1018_mask) begin
      pht_1_7[pht_1_7_MPORT_1018_addr] <= pht_1_7_MPORT_1018_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1020_en & pht_1_7_MPORT_1020_mask) begin
      pht_1_7[pht_1_7_MPORT_1020_addr] <= pht_1_7_MPORT_1020_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1022_en & pht_1_7_MPORT_1022_mask) begin
      pht_1_7[pht_1_7_MPORT_1022_addr] <= pht_1_7_MPORT_1022_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1024_en & pht_1_7_MPORT_1024_mask) begin
      pht_1_7[pht_1_7_MPORT_1024_addr] <= pht_1_7_MPORT_1024_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1026_en & pht_1_7_MPORT_1026_mask) begin
      pht_1_7[pht_1_7_MPORT_1026_addr] <= pht_1_7_MPORT_1026_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1028_en & pht_1_7_MPORT_1028_mask) begin
      pht_1_7[pht_1_7_MPORT_1028_addr] <= pht_1_7_MPORT_1028_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1030_en & pht_1_7_MPORT_1030_mask) begin
      pht_1_7[pht_1_7_MPORT_1030_addr] <= pht_1_7_MPORT_1030_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1032_en & pht_1_7_MPORT_1032_mask) begin
      pht_1_7[pht_1_7_MPORT_1032_addr] <= pht_1_7_MPORT_1032_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1034_en & pht_1_7_MPORT_1034_mask) begin
      pht_1_7[pht_1_7_MPORT_1034_addr] <= pht_1_7_MPORT_1034_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1036_en & pht_1_7_MPORT_1036_mask) begin
      pht_1_7[pht_1_7_MPORT_1036_addr] <= pht_1_7_MPORT_1036_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1038_en & pht_1_7_MPORT_1038_mask) begin
      pht_1_7[pht_1_7_MPORT_1038_addr] <= pht_1_7_MPORT_1038_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1040_en & pht_1_7_MPORT_1040_mask) begin
      pht_1_7[pht_1_7_MPORT_1040_addr] <= pht_1_7_MPORT_1040_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1042_en & pht_1_7_MPORT_1042_mask) begin
      pht_1_7[pht_1_7_MPORT_1042_addr] <= pht_1_7_MPORT_1042_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1044_en & pht_1_7_MPORT_1044_mask) begin
      pht_1_7[pht_1_7_MPORT_1044_addr] <= pht_1_7_MPORT_1044_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1046_en & pht_1_7_MPORT_1046_mask) begin
      pht_1_7[pht_1_7_MPORT_1046_addr] <= pht_1_7_MPORT_1046_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1048_en & pht_1_7_MPORT_1048_mask) begin
      pht_1_7[pht_1_7_MPORT_1048_addr] <= pht_1_7_MPORT_1048_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1050_en & pht_1_7_MPORT_1050_mask) begin
      pht_1_7[pht_1_7_MPORT_1050_addr] <= pht_1_7_MPORT_1050_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1052_en & pht_1_7_MPORT_1052_mask) begin
      pht_1_7[pht_1_7_MPORT_1052_addr] <= pht_1_7_MPORT_1052_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1054_en & pht_1_7_MPORT_1054_mask) begin
      pht_1_7[pht_1_7_MPORT_1054_addr] <= pht_1_7_MPORT_1054_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1056_en & pht_1_7_MPORT_1056_mask) begin
      pht_1_7[pht_1_7_MPORT_1056_addr] <= pht_1_7_MPORT_1056_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1058_en & pht_1_7_MPORT_1058_mask) begin
      pht_1_7[pht_1_7_MPORT_1058_addr] <= pht_1_7_MPORT_1058_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1060_en & pht_1_7_MPORT_1060_mask) begin
      pht_1_7[pht_1_7_MPORT_1060_addr] <= pht_1_7_MPORT_1060_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1062_en & pht_1_7_MPORT_1062_mask) begin
      pht_1_7[pht_1_7_MPORT_1062_addr] <= pht_1_7_MPORT_1062_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1064_en & pht_1_7_MPORT_1064_mask) begin
      pht_1_7[pht_1_7_MPORT_1064_addr] <= pht_1_7_MPORT_1064_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1066_en & pht_1_7_MPORT_1066_mask) begin
      pht_1_7[pht_1_7_MPORT_1066_addr] <= pht_1_7_MPORT_1066_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1068_en & pht_1_7_MPORT_1068_mask) begin
      pht_1_7[pht_1_7_MPORT_1068_addr] <= pht_1_7_MPORT_1068_data; // @[PatternHistoryTable.scala 21:28]
    end
    if (pht_1_7_MPORT_1070_en & pht_1_7_MPORT_1070_mask) begin
      pht_1_7[pht_1_7_MPORT_1070_addr] <= pht_1_7_MPORT_1070_data; // @[PatternHistoryTable.scala 21:28]
    end
//     pht_1_7_MPORT_7_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_7_MPORT_7_addr_pipe_0 <= io_raddr_0;
    end
//     pht_1_7_MPORT_15_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_7_MPORT_15_addr_pipe_0 <= io_raddr_1;
    end
//     pht_1_7_MPORT_30_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_1_7_MPORT_30_addr_pipe_0 <= io_waddr;
    end
    if (pht_0_0_MPORT_33_en & pht_0_0_MPORT_33_mask) begin
      pht_0_0[pht_0_0_MPORT_33_addr] <= pht_0_0_MPORT_33_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_49_en & pht_0_0_MPORT_49_mask) begin
      pht_0_0[pht_0_0_MPORT_49_addr] <= pht_0_0_MPORT_49_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_51_en & pht_0_0_MPORT_51_mask) begin
      pht_0_0[pht_0_0_MPORT_51_addr] <= pht_0_0_MPORT_51_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_53_en & pht_0_0_MPORT_53_mask) begin
      pht_0_0[pht_0_0_MPORT_53_addr] <= pht_0_0_MPORT_53_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_55_en & pht_0_0_MPORT_55_mask) begin
      pht_0_0[pht_0_0_MPORT_55_addr] <= pht_0_0_MPORT_55_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_57_en & pht_0_0_MPORT_57_mask) begin
      pht_0_0[pht_0_0_MPORT_57_addr] <= pht_0_0_MPORT_57_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_59_en & pht_0_0_MPORT_59_mask) begin
      pht_0_0[pht_0_0_MPORT_59_addr] <= pht_0_0_MPORT_59_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_61_en & pht_0_0_MPORT_61_mask) begin
      pht_0_0[pht_0_0_MPORT_61_addr] <= pht_0_0_MPORT_61_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_63_en & pht_0_0_MPORT_63_mask) begin
      pht_0_0[pht_0_0_MPORT_63_addr] <= pht_0_0_MPORT_63_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_65_en & pht_0_0_MPORT_65_mask) begin
      pht_0_0[pht_0_0_MPORT_65_addr] <= pht_0_0_MPORT_65_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_67_en & pht_0_0_MPORT_67_mask) begin
      pht_0_0[pht_0_0_MPORT_67_addr] <= pht_0_0_MPORT_67_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_69_en & pht_0_0_MPORT_69_mask) begin
      pht_0_0[pht_0_0_MPORT_69_addr] <= pht_0_0_MPORT_69_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_71_en & pht_0_0_MPORT_71_mask) begin
      pht_0_0[pht_0_0_MPORT_71_addr] <= pht_0_0_MPORT_71_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_73_en & pht_0_0_MPORT_73_mask) begin
      pht_0_0[pht_0_0_MPORT_73_addr] <= pht_0_0_MPORT_73_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_75_en & pht_0_0_MPORT_75_mask) begin
      pht_0_0[pht_0_0_MPORT_75_addr] <= pht_0_0_MPORT_75_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_77_en & pht_0_0_MPORT_77_mask) begin
      pht_0_0[pht_0_0_MPORT_77_addr] <= pht_0_0_MPORT_77_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_79_en & pht_0_0_MPORT_79_mask) begin
      pht_0_0[pht_0_0_MPORT_79_addr] <= pht_0_0_MPORT_79_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_81_en & pht_0_0_MPORT_81_mask) begin
      pht_0_0[pht_0_0_MPORT_81_addr] <= pht_0_0_MPORT_81_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_83_en & pht_0_0_MPORT_83_mask) begin
      pht_0_0[pht_0_0_MPORT_83_addr] <= pht_0_0_MPORT_83_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_85_en & pht_0_0_MPORT_85_mask) begin
      pht_0_0[pht_0_0_MPORT_85_addr] <= pht_0_0_MPORT_85_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_87_en & pht_0_0_MPORT_87_mask) begin
      pht_0_0[pht_0_0_MPORT_87_addr] <= pht_0_0_MPORT_87_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_89_en & pht_0_0_MPORT_89_mask) begin
      pht_0_0[pht_0_0_MPORT_89_addr] <= pht_0_0_MPORT_89_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_91_en & pht_0_0_MPORT_91_mask) begin
      pht_0_0[pht_0_0_MPORT_91_addr] <= pht_0_0_MPORT_91_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_93_en & pht_0_0_MPORT_93_mask) begin
      pht_0_0[pht_0_0_MPORT_93_addr] <= pht_0_0_MPORT_93_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_95_en & pht_0_0_MPORT_95_mask) begin
      pht_0_0[pht_0_0_MPORT_95_addr] <= pht_0_0_MPORT_95_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_97_en & pht_0_0_MPORT_97_mask) begin
      pht_0_0[pht_0_0_MPORT_97_addr] <= pht_0_0_MPORT_97_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_99_en & pht_0_0_MPORT_99_mask) begin
      pht_0_0[pht_0_0_MPORT_99_addr] <= pht_0_0_MPORT_99_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_101_en & pht_0_0_MPORT_101_mask) begin
      pht_0_0[pht_0_0_MPORT_101_addr] <= pht_0_0_MPORT_101_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_103_en & pht_0_0_MPORT_103_mask) begin
      pht_0_0[pht_0_0_MPORT_103_addr] <= pht_0_0_MPORT_103_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_105_en & pht_0_0_MPORT_105_mask) begin
      pht_0_0[pht_0_0_MPORT_105_addr] <= pht_0_0_MPORT_105_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_107_en & pht_0_0_MPORT_107_mask) begin
      pht_0_0[pht_0_0_MPORT_107_addr] <= pht_0_0_MPORT_107_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_109_en & pht_0_0_MPORT_109_mask) begin
      pht_0_0[pht_0_0_MPORT_109_addr] <= pht_0_0_MPORT_109_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_111_en & pht_0_0_MPORT_111_mask) begin
      pht_0_0[pht_0_0_MPORT_111_addr] <= pht_0_0_MPORT_111_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_113_en & pht_0_0_MPORT_113_mask) begin
      pht_0_0[pht_0_0_MPORT_113_addr] <= pht_0_0_MPORT_113_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_115_en & pht_0_0_MPORT_115_mask) begin
      pht_0_0[pht_0_0_MPORT_115_addr] <= pht_0_0_MPORT_115_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_117_en & pht_0_0_MPORT_117_mask) begin
      pht_0_0[pht_0_0_MPORT_117_addr] <= pht_0_0_MPORT_117_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_119_en & pht_0_0_MPORT_119_mask) begin
      pht_0_0[pht_0_0_MPORT_119_addr] <= pht_0_0_MPORT_119_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_121_en & pht_0_0_MPORT_121_mask) begin
      pht_0_0[pht_0_0_MPORT_121_addr] <= pht_0_0_MPORT_121_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_123_en & pht_0_0_MPORT_123_mask) begin
      pht_0_0[pht_0_0_MPORT_123_addr] <= pht_0_0_MPORT_123_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_125_en & pht_0_0_MPORT_125_mask) begin
      pht_0_0[pht_0_0_MPORT_125_addr] <= pht_0_0_MPORT_125_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_127_en & pht_0_0_MPORT_127_mask) begin
      pht_0_0[pht_0_0_MPORT_127_addr] <= pht_0_0_MPORT_127_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_129_en & pht_0_0_MPORT_129_mask) begin
      pht_0_0[pht_0_0_MPORT_129_addr] <= pht_0_0_MPORT_129_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_131_en & pht_0_0_MPORT_131_mask) begin
      pht_0_0[pht_0_0_MPORT_131_addr] <= pht_0_0_MPORT_131_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_133_en & pht_0_0_MPORT_133_mask) begin
      pht_0_0[pht_0_0_MPORT_133_addr] <= pht_0_0_MPORT_133_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_135_en & pht_0_0_MPORT_135_mask) begin
      pht_0_0[pht_0_0_MPORT_135_addr] <= pht_0_0_MPORT_135_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_137_en & pht_0_0_MPORT_137_mask) begin
      pht_0_0[pht_0_0_MPORT_137_addr] <= pht_0_0_MPORT_137_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_139_en & pht_0_0_MPORT_139_mask) begin
      pht_0_0[pht_0_0_MPORT_139_addr] <= pht_0_0_MPORT_139_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_141_en & pht_0_0_MPORT_141_mask) begin
      pht_0_0[pht_0_0_MPORT_141_addr] <= pht_0_0_MPORT_141_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_143_en & pht_0_0_MPORT_143_mask) begin
      pht_0_0[pht_0_0_MPORT_143_addr] <= pht_0_0_MPORT_143_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_145_en & pht_0_0_MPORT_145_mask) begin
      pht_0_0[pht_0_0_MPORT_145_addr] <= pht_0_0_MPORT_145_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_147_en & pht_0_0_MPORT_147_mask) begin
      pht_0_0[pht_0_0_MPORT_147_addr] <= pht_0_0_MPORT_147_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_149_en & pht_0_0_MPORT_149_mask) begin
      pht_0_0[pht_0_0_MPORT_149_addr] <= pht_0_0_MPORT_149_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_151_en & pht_0_0_MPORT_151_mask) begin
      pht_0_0[pht_0_0_MPORT_151_addr] <= pht_0_0_MPORT_151_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_153_en & pht_0_0_MPORT_153_mask) begin
      pht_0_0[pht_0_0_MPORT_153_addr] <= pht_0_0_MPORT_153_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_155_en & pht_0_0_MPORT_155_mask) begin
      pht_0_0[pht_0_0_MPORT_155_addr] <= pht_0_0_MPORT_155_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_157_en & pht_0_0_MPORT_157_mask) begin
      pht_0_0[pht_0_0_MPORT_157_addr] <= pht_0_0_MPORT_157_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_159_en & pht_0_0_MPORT_159_mask) begin
      pht_0_0[pht_0_0_MPORT_159_addr] <= pht_0_0_MPORT_159_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_161_en & pht_0_0_MPORT_161_mask) begin
      pht_0_0[pht_0_0_MPORT_161_addr] <= pht_0_0_MPORT_161_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_163_en & pht_0_0_MPORT_163_mask) begin
      pht_0_0[pht_0_0_MPORT_163_addr] <= pht_0_0_MPORT_163_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_165_en & pht_0_0_MPORT_165_mask) begin
      pht_0_0[pht_0_0_MPORT_165_addr] <= pht_0_0_MPORT_165_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_167_en & pht_0_0_MPORT_167_mask) begin
      pht_0_0[pht_0_0_MPORT_167_addr] <= pht_0_0_MPORT_167_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_169_en & pht_0_0_MPORT_169_mask) begin
      pht_0_0[pht_0_0_MPORT_169_addr] <= pht_0_0_MPORT_169_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_171_en & pht_0_0_MPORT_171_mask) begin
      pht_0_0[pht_0_0_MPORT_171_addr] <= pht_0_0_MPORT_171_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_173_en & pht_0_0_MPORT_173_mask) begin
      pht_0_0[pht_0_0_MPORT_173_addr] <= pht_0_0_MPORT_173_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_0_MPORT_175_en & pht_0_0_MPORT_175_mask) begin
      pht_0_0[pht_0_0_MPORT_175_addr] <= pht_0_0_MPORT_175_data; // @[PatternHistoryTable.scala 26:28]
    end
//     pht_0_0_MPORT_17_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_0_0_MPORT_17_addr_pipe_0 <= io_waddr;
    end
    if (pht_0_1_MPORT_35_en & pht_0_1_MPORT_35_mask) begin
      pht_0_1[pht_0_1_MPORT_35_addr] <= pht_0_1_MPORT_35_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_177_en & pht_0_1_MPORT_177_mask) begin
      pht_0_1[pht_0_1_MPORT_177_addr] <= pht_0_1_MPORT_177_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_179_en & pht_0_1_MPORT_179_mask) begin
      pht_0_1[pht_0_1_MPORT_179_addr] <= pht_0_1_MPORT_179_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_181_en & pht_0_1_MPORT_181_mask) begin
      pht_0_1[pht_0_1_MPORT_181_addr] <= pht_0_1_MPORT_181_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_183_en & pht_0_1_MPORT_183_mask) begin
      pht_0_1[pht_0_1_MPORT_183_addr] <= pht_0_1_MPORT_183_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_185_en & pht_0_1_MPORT_185_mask) begin
      pht_0_1[pht_0_1_MPORT_185_addr] <= pht_0_1_MPORT_185_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_187_en & pht_0_1_MPORT_187_mask) begin
      pht_0_1[pht_0_1_MPORT_187_addr] <= pht_0_1_MPORT_187_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_189_en & pht_0_1_MPORT_189_mask) begin
      pht_0_1[pht_0_1_MPORT_189_addr] <= pht_0_1_MPORT_189_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_191_en & pht_0_1_MPORT_191_mask) begin
      pht_0_1[pht_0_1_MPORT_191_addr] <= pht_0_1_MPORT_191_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_193_en & pht_0_1_MPORT_193_mask) begin
      pht_0_1[pht_0_1_MPORT_193_addr] <= pht_0_1_MPORT_193_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_195_en & pht_0_1_MPORT_195_mask) begin
      pht_0_1[pht_0_1_MPORT_195_addr] <= pht_0_1_MPORT_195_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_197_en & pht_0_1_MPORT_197_mask) begin
      pht_0_1[pht_0_1_MPORT_197_addr] <= pht_0_1_MPORT_197_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_199_en & pht_0_1_MPORT_199_mask) begin
      pht_0_1[pht_0_1_MPORT_199_addr] <= pht_0_1_MPORT_199_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_201_en & pht_0_1_MPORT_201_mask) begin
      pht_0_1[pht_0_1_MPORT_201_addr] <= pht_0_1_MPORT_201_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_203_en & pht_0_1_MPORT_203_mask) begin
      pht_0_1[pht_0_1_MPORT_203_addr] <= pht_0_1_MPORT_203_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_205_en & pht_0_1_MPORT_205_mask) begin
      pht_0_1[pht_0_1_MPORT_205_addr] <= pht_0_1_MPORT_205_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_207_en & pht_0_1_MPORT_207_mask) begin
      pht_0_1[pht_0_1_MPORT_207_addr] <= pht_0_1_MPORT_207_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_209_en & pht_0_1_MPORT_209_mask) begin
      pht_0_1[pht_0_1_MPORT_209_addr] <= pht_0_1_MPORT_209_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_211_en & pht_0_1_MPORT_211_mask) begin
      pht_0_1[pht_0_1_MPORT_211_addr] <= pht_0_1_MPORT_211_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_213_en & pht_0_1_MPORT_213_mask) begin
      pht_0_1[pht_0_1_MPORT_213_addr] <= pht_0_1_MPORT_213_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_215_en & pht_0_1_MPORT_215_mask) begin
      pht_0_1[pht_0_1_MPORT_215_addr] <= pht_0_1_MPORT_215_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_217_en & pht_0_1_MPORT_217_mask) begin
      pht_0_1[pht_0_1_MPORT_217_addr] <= pht_0_1_MPORT_217_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_219_en & pht_0_1_MPORT_219_mask) begin
      pht_0_1[pht_0_1_MPORT_219_addr] <= pht_0_1_MPORT_219_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_221_en & pht_0_1_MPORT_221_mask) begin
      pht_0_1[pht_0_1_MPORT_221_addr] <= pht_0_1_MPORT_221_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_223_en & pht_0_1_MPORT_223_mask) begin
      pht_0_1[pht_0_1_MPORT_223_addr] <= pht_0_1_MPORT_223_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_225_en & pht_0_1_MPORT_225_mask) begin
      pht_0_1[pht_0_1_MPORT_225_addr] <= pht_0_1_MPORT_225_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_227_en & pht_0_1_MPORT_227_mask) begin
      pht_0_1[pht_0_1_MPORT_227_addr] <= pht_0_1_MPORT_227_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_229_en & pht_0_1_MPORT_229_mask) begin
      pht_0_1[pht_0_1_MPORT_229_addr] <= pht_0_1_MPORT_229_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_231_en & pht_0_1_MPORT_231_mask) begin
      pht_0_1[pht_0_1_MPORT_231_addr] <= pht_0_1_MPORT_231_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_233_en & pht_0_1_MPORT_233_mask) begin
      pht_0_1[pht_0_1_MPORT_233_addr] <= pht_0_1_MPORT_233_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_235_en & pht_0_1_MPORT_235_mask) begin
      pht_0_1[pht_0_1_MPORT_235_addr] <= pht_0_1_MPORT_235_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_237_en & pht_0_1_MPORT_237_mask) begin
      pht_0_1[pht_0_1_MPORT_237_addr] <= pht_0_1_MPORT_237_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_239_en & pht_0_1_MPORT_239_mask) begin
      pht_0_1[pht_0_1_MPORT_239_addr] <= pht_0_1_MPORT_239_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_241_en & pht_0_1_MPORT_241_mask) begin
      pht_0_1[pht_0_1_MPORT_241_addr] <= pht_0_1_MPORT_241_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_243_en & pht_0_1_MPORT_243_mask) begin
      pht_0_1[pht_0_1_MPORT_243_addr] <= pht_0_1_MPORT_243_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_245_en & pht_0_1_MPORT_245_mask) begin
      pht_0_1[pht_0_1_MPORT_245_addr] <= pht_0_1_MPORT_245_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_247_en & pht_0_1_MPORT_247_mask) begin
      pht_0_1[pht_0_1_MPORT_247_addr] <= pht_0_1_MPORT_247_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_249_en & pht_0_1_MPORT_249_mask) begin
      pht_0_1[pht_0_1_MPORT_249_addr] <= pht_0_1_MPORT_249_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_251_en & pht_0_1_MPORT_251_mask) begin
      pht_0_1[pht_0_1_MPORT_251_addr] <= pht_0_1_MPORT_251_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_253_en & pht_0_1_MPORT_253_mask) begin
      pht_0_1[pht_0_1_MPORT_253_addr] <= pht_0_1_MPORT_253_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_255_en & pht_0_1_MPORT_255_mask) begin
      pht_0_1[pht_0_1_MPORT_255_addr] <= pht_0_1_MPORT_255_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_257_en & pht_0_1_MPORT_257_mask) begin
      pht_0_1[pht_0_1_MPORT_257_addr] <= pht_0_1_MPORT_257_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_259_en & pht_0_1_MPORT_259_mask) begin
      pht_0_1[pht_0_1_MPORT_259_addr] <= pht_0_1_MPORT_259_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_261_en & pht_0_1_MPORT_261_mask) begin
      pht_0_1[pht_0_1_MPORT_261_addr] <= pht_0_1_MPORT_261_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_263_en & pht_0_1_MPORT_263_mask) begin
      pht_0_1[pht_0_1_MPORT_263_addr] <= pht_0_1_MPORT_263_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_265_en & pht_0_1_MPORT_265_mask) begin
      pht_0_1[pht_0_1_MPORT_265_addr] <= pht_0_1_MPORT_265_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_267_en & pht_0_1_MPORT_267_mask) begin
      pht_0_1[pht_0_1_MPORT_267_addr] <= pht_0_1_MPORT_267_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_269_en & pht_0_1_MPORT_269_mask) begin
      pht_0_1[pht_0_1_MPORT_269_addr] <= pht_0_1_MPORT_269_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_271_en & pht_0_1_MPORT_271_mask) begin
      pht_0_1[pht_0_1_MPORT_271_addr] <= pht_0_1_MPORT_271_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_273_en & pht_0_1_MPORT_273_mask) begin
      pht_0_1[pht_0_1_MPORT_273_addr] <= pht_0_1_MPORT_273_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_275_en & pht_0_1_MPORT_275_mask) begin
      pht_0_1[pht_0_1_MPORT_275_addr] <= pht_0_1_MPORT_275_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_277_en & pht_0_1_MPORT_277_mask) begin
      pht_0_1[pht_0_1_MPORT_277_addr] <= pht_0_1_MPORT_277_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_279_en & pht_0_1_MPORT_279_mask) begin
      pht_0_1[pht_0_1_MPORT_279_addr] <= pht_0_1_MPORT_279_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_281_en & pht_0_1_MPORT_281_mask) begin
      pht_0_1[pht_0_1_MPORT_281_addr] <= pht_0_1_MPORT_281_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_283_en & pht_0_1_MPORT_283_mask) begin
      pht_0_1[pht_0_1_MPORT_283_addr] <= pht_0_1_MPORT_283_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_285_en & pht_0_1_MPORT_285_mask) begin
      pht_0_1[pht_0_1_MPORT_285_addr] <= pht_0_1_MPORT_285_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_287_en & pht_0_1_MPORT_287_mask) begin
      pht_0_1[pht_0_1_MPORT_287_addr] <= pht_0_1_MPORT_287_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_289_en & pht_0_1_MPORT_289_mask) begin
      pht_0_1[pht_0_1_MPORT_289_addr] <= pht_0_1_MPORT_289_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_291_en & pht_0_1_MPORT_291_mask) begin
      pht_0_1[pht_0_1_MPORT_291_addr] <= pht_0_1_MPORT_291_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_293_en & pht_0_1_MPORT_293_mask) begin
      pht_0_1[pht_0_1_MPORT_293_addr] <= pht_0_1_MPORT_293_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_295_en & pht_0_1_MPORT_295_mask) begin
      pht_0_1[pht_0_1_MPORT_295_addr] <= pht_0_1_MPORT_295_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_297_en & pht_0_1_MPORT_297_mask) begin
      pht_0_1[pht_0_1_MPORT_297_addr] <= pht_0_1_MPORT_297_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_299_en & pht_0_1_MPORT_299_mask) begin
      pht_0_1[pht_0_1_MPORT_299_addr] <= pht_0_1_MPORT_299_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_301_en & pht_0_1_MPORT_301_mask) begin
      pht_0_1[pht_0_1_MPORT_301_addr] <= pht_0_1_MPORT_301_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_1_MPORT_303_en & pht_0_1_MPORT_303_mask) begin
      pht_0_1[pht_0_1_MPORT_303_addr] <= pht_0_1_MPORT_303_data; // @[PatternHistoryTable.scala 26:28]
    end
//     pht_0_1_MPORT_19_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_0_1_MPORT_19_addr_pipe_0 <= io_waddr;
    end
    if (pht_0_2_MPORT_37_en & pht_0_2_MPORT_37_mask) begin
      pht_0_2[pht_0_2_MPORT_37_addr] <= pht_0_2_MPORT_37_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_305_en & pht_0_2_MPORT_305_mask) begin
      pht_0_2[pht_0_2_MPORT_305_addr] <= pht_0_2_MPORT_305_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_307_en & pht_0_2_MPORT_307_mask) begin
      pht_0_2[pht_0_2_MPORT_307_addr] <= pht_0_2_MPORT_307_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_309_en & pht_0_2_MPORT_309_mask) begin
      pht_0_2[pht_0_2_MPORT_309_addr] <= pht_0_2_MPORT_309_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_311_en & pht_0_2_MPORT_311_mask) begin
      pht_0_2[pht_0_2_MPORT_311_addr] <= pht_0_2_MPORT_311_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_313_en & pht_0_2_MPORT_313_mask) begin
      pht_0_2[pht_0_2_MPORT_313_addr] <= pht_0_2_MPORT_313_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_315_en & pht_0_2_MPORT_315_mask) begin
      pht_0_2[pht_0_2_MPORT_315_addr] <= pht_0_2_MPORT_315_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_317_en & pht_0_2_MPORT_317_mask) begin
      pht_0_2[pht_0_2_MPORT_317_addr] <= pht_0_2_MPORT_317_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_319_en & pht_0_2_MPORT_319_mask) begin
      pht_0_2[pht_0_2_MPORT_319_addr] <= pht_0_2_MPORT_319_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_321_en & pht_0_2_MPORT_321_mask) begin
      pht_0_2[pht_0_2_MPORT_321_addr] <= pht_0_2_MPORT_321_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_323_en & pht_0_2_MPORT_323_mask) begin
      pht_0_2[pht_0_2_MPORT_323_addr] <= pht_0_2_MPORT_323_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_325_en & pht_0_2_MPORT_325_mask) begin
      pht_0_2[pht_0_2_MPORT_325_addr] <= pht_0_2_MPORT_325_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_327_en & pht_0_2_MPORT_327_mask) begin
      pht_0_2[pht_0_2_MPORT_327_addr] <= pht_0_2_MPORT_327_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_329_en & pht_0_2_MPORT_329_mask) begin
      pht_0_2[pht_0_2_MPORT_329_addr] <= pht_0_2_MPORT_329_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_331_en & pht_0_2_MPORT_331_mask) begin
      pht_0_2[pht_0_2_MPORT_331_addr] <= pht_0_2_MPORT_331_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_333_en & pht_0_2_MPORT_333_mask) begin
      pht_0_2[pht_0_2_MPORT_333_addr] <= pht_0_2_MPORT_333_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_335_en & pht_0_2_MPORT_335_mask) begin
      pht_0_2[pht_0_2_MPORT_335_addr] <= pht_0_2_MPORT_335_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_337_en & pht_0_2_MPORT_337_mask) begin
      pht_0_2[pht_0_2_MPORT_337_addr] <= pht_0_2_MPORT_337_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_339_en & pht_0_2_MPORT_339_mask) begin
      pht_0_2[pht_0_2_MPORT_339_addr] <= pht_0_2_MPORT_339_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_341_en & pht_0_2_MPORT_341_mask) begin
      pht_0_2[pht_0_2_MPORT_341_addr] <= pht_0_2_MPORT_341_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_343_en & pht_0_2_MPORT_343_mask) begin
      pht_0_2[pht_0_2_MPORT_343_addr] <= pht_0_2_MPORT_343_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_345_en & pht_0_2_MPORT_345_mask) begin
      pht_0_2[pht_0_2_MPORT_345_addr] <= pht_0_2_MPORT_345_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_347_en & pht_0_2_MPORT_347_mask) begin
      pht_0_2[pht_0_2_MPORT_347_addr] <= pht_0_2_MPORT_347_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_349_en & pht_0_2_MPORT_349_mask) begin
      pht_0_2[pht_0_2_MPORT_349_addr] <= pht_0_2_MPORT_349_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_351_en & pht_0_2_MPORT_351_mask) begin
      pht_0_2[pht_0_2_MPORT_351_addr] <= pht_0_2_MPORT_351_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_353_en & pht_0_2_MPORT_353_mask) begin
      pht_0_2[pht_0_2_MPORT_353_addr] <= pht_0_2_MPORT_353_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_355_en & pht_0_2_MPORT_355_mask) begin
      pht_0_2[pht_0_2_MPORT_355_addr] <= pht_0_2_MPORT_355_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_357_en & pht_0_2_MPORT_357_mask) begin
      pht_0_2[pht_0_2_MPORT_357_addr] <= pht_0_2_MPORT_357_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_359_en & pht_0_2_MPORT_359_mask) begin
      pht_0_2[pht_0_2_MPORT_359_addr] <= pht_0_2_MPORT_359_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_361_en & pht_0_2_MPORT_361_mask) begin
      pht_0_2[pht_0_2_MPORT_361_addr] <= pht_0_2_MPORT_361_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_363_en & pht_0_2_MPORT_363_mask) begin
      pht_0_2[pht_0_2_MPORT_363_addr] <= pht_0_2_MPORT_363_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_365_en & pht_0_2_MPORT_365_mask) begin
      pht_0_2[pht_0_2_MPORT_365_addr] <= pht_0_2_MPORT_365_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_367_en & pht_0_2_MPORT_367_mask) begin
      pht_0_2[pht_0_2_MPORT_367_addr] <= pht_0_2_MPORT_367_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_369_en & pht_0_2_MPORT_369_mask) begin
      pht_0_2[pht_0_2_MPORT_369_addr] <= pht_0_2_MPORT_369_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_371_en & pht_0_2_MPORT_371_mask) begin
      pht_0_2[pht_0_2_MPORT_371_addr] <= pht_0_2_MPORT_371_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_373_en & pht_0_2_MPORT_373_mask) begin
      pht_0_2[pht_0_2_MPORT_373_addr] <= pht_0_2_MPORT_373_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_375_en & pht_0_2_MPORT_375_mask) begin
      pht_0_2[pht_0_2_MPORT_375_addr] <= pht_0_2_MPORT_375_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_377_en & pht_0_2_MPORT_377_mask) begin
      pht_0_2[pht_0_2_MPORT_377_addr] <= pht_0_2_MPORT_377_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_379_en & pht_0_2_MPORT_379_mask) begin
      pht_0_2[pht_0_2_MPORT_379_addr] <= pht_0_2_MPORT_379_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_381_en & pht_0_2_MPORT_381_mask) begin
      pht_0_2[pht_0_2_MPORT_381_addr] <= pht_0_2_MPORT_381_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_383_en & pht_0_2_MPORT_383_mask) begin
      pht_0_2[pht_0_2_MPORT_383_addr] <= pht_0_2_MPORT_383_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_385_en & pht_0_2_MPORT_385_mask) begin
      pht_0_2[pht_0_2_MPORT_385_addr] <= pht_0_2_MPORT_385_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_387_en & pht_0_2_MPORT_387_mask) begin
      pht_0_2[pht_0_2_MPORT_387_addr] <= pht_0_2_MPORT_387_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_389_en & pht_0_2_MPORT_389_mask) begin
      pht_0_2[pht_0_2_MPORT_389_addr] <= pht_0_2_MPORT_389_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_391_en & pht_0_2_MPORT_391_mask) begin
      pht_0_2[pht_0_2_MPORT_391_addr] <= pht_0_2_MPORT_391_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_393_en & pht_0_2_MPORT_393_mask) begin
      pht_0_2[pht_0_2_MPORT_393_addr] <= pht_0_2_MPORT_393_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_395_en & pht_0_2_MPORT_395_mask) begin
      pht_0_2[pht_0_2_MPORT_395_addr] <= pht_0_2_MPORT_395_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_397_en & pht_0_2_MPORT_397_mask) begin
      pht_0_2[pht_0_2_MPORT_397_addr] <= pht_0_2_MPORT_397_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_399_en & pht_0_2_MPORT_399_mask) begin
      pht_0_2[pht_0_2_MPORT_399_addr] <= pht_0_2_MPORT_399_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_401_en & pht_0_2_MPORT_401_mask) begin
      pht_0_2[pht_0_2_MPORT_401_addr] <= pht_0_2_MPORT_401_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_403_en & pht_0_2_MPORT_403_mask) begin
      pht_0_2[pht_0_2_MPORT_403_addr] <= pht_0_2_MPORT_403_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_405_en & pht_0_2_MPORT_405_mask) begin
      pht_0_2[pht_0_2_MPORT_405_addr] <= pht_0_2_MPORT_405_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_407_en & pht_0_2_MPORT_407_mask) begin
      pht_0_2[pht_0_2_MPORT_407_addr] <= pht_0_2_MPORT_407_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_409_en & pht_0_2_MPORT_409_mask) begin
      pht_0_2[pht_0_2_MPORT_409_addr] <= pht_0_2_MPORT_409_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_411_en & pht_0_2_MPORT_411_mask) begin
      pht_0_2[pht_0_2_MPORT_411_addr] <= pht_0_2_MPORT_411_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_413_en & pht_0_2_MPORT_413_mask) begin
      pht_0_2[pht_0_2_MPORT_413_addr] <= pht_0_2_MPORT_413_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_415_en & pht_0_2_MPORT_415_mask) begin
      pht_0_2[pht_0_2_MPORT_415_addr] <= pht_0_2_MPORT_415_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_417_en & pht_0_2_MPORT_417_mask) begin
      pht_0_2[pht_0_2_MPORT_417_addr] <= pht_0_2_MPORT_417_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_419_en & pht_0_2_MPORT_419_mask) begin
      pht_0_2[pht_0_2_MPORT_419_addr] <= pht_0_2_MPORT_419_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_421_en & pht_0_2_MPORT_421_mask) begin
      pht_0_2[pht_0_2_MPORT_421_addr] <= pht_0_2_MPORT_421_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_423_en & pht_0_2_MPORT_423_mask) begin
      pht_0_2[pht_0_2_MPORT_423_addr] <= pht_0_2_MPORT_423_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_425_en & pht_0_2_MPORT_425_mask) begin
      pht_0_2[pht_0_2_MPORT_425_addr] <= pht_0_2_MPORT_425_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_427_en & pht_0_2_MPORT_427_mask) begin
      pht_0_2[pht_0_2_MPORT_427_addr] <= pht_0_2_MPORT_427_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_429_en & pht_0_2_MPORT_429_mask) begin
      pht_0_2[pht_0_2_MPORT_429_addr] <= pht_0_2_MPORT_429_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_2_MPORT_431_en & pht_0_2_MPORT_431_mask) begin
      pht_0_2[pht_0_2_MPORT_431_addr] <= pht_0_2_MPORT_431_data; // @[PatternHistoryTable.scala 26:28]
    end
//     pht_0_2_MPORT_21_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_0_2_MPORT_21_addr_pipe_0 <= io_waddr;
    end
    if (pht_0_3_MPORT_39_en & pht_0_3_MPORT_39_mask) begin
      pht_0_3[pht_0_3_MPORT_39_addr] <= pht_0_3_MPORT_39_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_433_en & pht_0_3_MPORT_433_mask) begin
      pht_0_3[pht_0_3_MPORT_433_addr] <= pht_0_3_MPORT_433_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_435_en & pht_0_3_MPORT_435_mask) begin
      pht_0_3[pht_0_3_MPORT_435_addr] <= pht_0_3_MPORT_435_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_437_en & pht_0_3_MPORT_437_mask) begin
      pht_0_3[pht_0_3_MPORT_437_addr] <= pht_0_3_MPORT_437_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_439_en & pht_0_3_MPORT_439_mask) begin
      pht_0_3[pht_0_3_MPORT_439_addr] <= pht_0_3_MPORT_439_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_441_en & pht_0_3_MPORT_441_mask) begin
      pht_0_3[pht_0_3_MPORT_441_addr] <= pht_0_3_MPORT_441_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_443_en & pht_0_3_MPORT_443_mask) begin
      pht_0_3[pht_0_3_MPORT_443_addr] <= pht_0_3_MPORT_443_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_445_en & pht_0_3_MPORT_445_mask) begin
      pht_0_3[pht_0_3_MPORT_445_addr] <= pht_0_3_MPORT_445_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_447_en & pht_0_3_MPORT_447_mask) begin
      pht_0_3[pht_0_3_MPORT_447_addr] <= pht_0_3_MPORT_447_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_449_en & pht_0_3_MPORT_449_mask) begin
      pht_0_3[pht_0_3_MPORT_449_addr] <= pht_0_3_MPORT_449_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_451_en & pht_0_3_MPORT_451_mask) begin
      pht_0_3[pht_0_3_MPORT_451_addr] <= pht_0_3_MPORT_451_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_453_en & pht_0_3_MPORT_453_mask) begin
      pht_0_3[pht_0_3_MPORT_453_addr] <= pht_0_3_MPORT_453_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_455_en & pht_0_3_MPORT_455_mask) begin
      pht_0_3[pht_0_3_MPORT_455_addr] <= pht_0_3_MPORT_455_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_457_en & pht_0_3_MPORT_457_mask) begin
      pht_0_3[pht_0_3_MPORT_457_addr] <= pht_0_3_MPORT_457_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_459_en & pht_0_3_MPORT_459_mask) begin
      pht_0_3[pht_0_3_MPORT_459_addr] <= pht_0_3_MPORT_459_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_461_en & pht_0_3_MPORT_461_mask) begin
      pht_0_3[pht_0_3_MPORT_461_addr] <= pht_0_3_MPORT_461_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_463_en & pht_0_3_MPORT_463_mask) begin
      pht_0_3[pht_0_3_MPORT_463_addr] <= pht_0_3_MPORT_463_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_465_en & pht_0_3_MPORT_465_mask) begin
      pht_0_3[pht_0_3_MPORT_465_addr] <= pht_0_3_MPORT_465_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_467_en & pht_0_3_MPORT_467_mask) begin
      pht_0_3[pht_0_3_MPORT_467_addr] <= pht_0_3_MPORT_467_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_469_en & pht_0_3_MPORT_469_mask) begin
      pht_0_3[pht_0_3_MPORT_469_addr] <= pht_0_3_MPORT_469_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_471_en & pht_0_3_MPORT_471_mask) begin
      pht_0_3[pht_0_3_MPORT_471_addr] <= pht_0_3_MPORT_471_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_473_en & pht_0_3_MPORT_473_mask) begin
      pht_0_3[pht_0_3_MPORT_473_addr] <= pht_0_3_MPORT_473_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_475_en & pht_0_3_MPORT_475_mask) begin
      pht_0_3[pht_0_3_MPORT_475_addr] <= pht_0_3_MPORT_475_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_477_en & pht_0_3_MPORT_477_mask) begin
      pht_0_3[pht_0_3_MPORT_477_addr] <= pht_0_3_MPORT_477_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_479_en & pht_0_3_MPORT_479_mask) begin
      pht_0_3[pht_0_3_MPORT_479_addr] <= pht_0_3_MPORT_479_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_481_en & pht_0_3_MPORT_481_mask) begin
      pht_0_3[pht_0_3_MPORT_481_addr] <= pht_0_3_MPORT_481_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_483_en & pht_0_3_MPORT_483_mask) begin
      pht_0_3[pht_0_3_MPORT_483_addr] <= pht_0_3_MPORT_483_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_485_en & pht_0_3_MPORT_485_mask) begin
      pht_0_3[pht_0_3_MPORT_485_addr] <= pht_0_3_MPORT_485_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_487_en & pht_0_3_MPORT_487_mask) begin
      pht_0_3[pht_0_3_MPORT_487_addr] <= pht_0_3_MPORT_487_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_489_en & pht_0_3_MPORT_489_mask) begin
      pht_0_3[pht_0_3_MPORT_489_addr] <= pht_0_3_MPORT_489_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_491_en & pht_0_3_MPORT_491_mask) begin
      pht_0_3[pht_0_3_MPORT_491_addr] <= pht_0_3_MPORT_491_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_493_en & pht_0_3_MPORT_493_mask) begin
      pht_0_3[pht_0_3_MPORT_493_addr] <= pht_0_3_MPORT_493_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_495_en & pht_0_3_MPORT_495_mask) begin
      pht_0_3[pht_0_3_MPORT_495_addr] <= pht_0_3_MPORT_495_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_497_en & pht_0_3_MPORT_497_mask) begin
      pht_0_3[pht_0_3_MPORT_497_addr] <= pht_0_3_MPORT_497_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_499_en & pht_0_3_MPORT_499_mask) begin
      pht_0_3[pht_0_3_MPORT_499_addr] <= pht_0_3_MPORT_499_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_501_en & pht_0_3_MPORT_501_mask) begin
      pht_0_3[pht_0_3_MPORT_501_addr] <= pht_0_3_MPORT_501_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_503_en & pht_0_3_MPORT_503_mask) begin
      pht_0_3[pht_0_3_MPORT_503_addr] <= pht_0_3_MPORT_503_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_505_en & pht_0_3_MPORT_505_mask) begin
      pht_0_3[pht_0_3_MPORT_505_addr] <= pht_0_3_MPORT_505_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_507_en & pht_0_3_MPORT_507_mask) begin
      pht_0_3[pht_0_3_MPORT_507_addr] <= pht_0_3_MPORT_507_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_509_en & pht_0_3_MPORT_509_mask) begin
      pht_0_3[pht_0_3_MPORT_509_addr] <= pht_0_3_MPORT_509_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_511_en & pht_0_3_MPORT_511_mask) begin
      pht_0_3[pht_0_3_MPORT_511_addr] <= pht_0_3_MPORT_511_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_513_en & pht_0_3_MPORT_513_mask) begin
      pht_0_3[pht_0_3_MPORT_513_addr] <= pht_0_3_MPORT_513_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_515_en & pht_0_3_MPORT_515_mask) begin
      pht_0_3[pht_0_3_MPORT_515_addr] <= pht_0_3_MPORT_515_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_517_en & pht_0_3_MPORT_517_mask) begin
      pht_0_3[pht_0_3_MPORT_517_addr] <= pht_0_3_MPORT_517_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_519_en & pht_0_3_MPORT_519_mask) begin
      pht_0_3[pht_0_3_MPORT_519_addr] <= pht_0_3_MPORT_519_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_521_en & pht_0_3_MPORT_521_mask) begin
      pht_0_3[pht_0_3_MPORT_521_addr] <= pht_0_3_MPORT_521_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_523_en & pht_0_3_MPORT_523_mask) begin
      pht_0_3[pht_0_3_MPORT_523_addr] <= pht_0_3_MPORT_523_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_525_en & pht_0_3_MPORT_525_mask) begin
      pht_0_3[pht_0_3_MPORT_525_addr] <= pht_0_3_MPORT_525_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_527_en & pht_0_3_MPORT_527_mask) begin
      pht_0_3[pht_0_3_MPORT_527_addr] <= pht_0_3_MPORT_527_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_529_en & pht_0_3_MPORT_529_mask) begin
      pht_0_3[pht_0_3_MPORT_529_addr] <= pht_0_3_MPORT_529_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_531_en & pht_0_3_MPORT_531_mask) begin
      pht_0_3[pht_0_3_MPORT_531_addr] <= pht_0_3_MPORT_531_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_533_en & pht_0_3_MPORT_533_mask) begin
      pht_0_3[pht_0_3_MPORT_533_addr] <= pht_0_3_MPORT_533_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_535_en & pht_0_3_MPORT_535_mask) begin
      pht_0_3[pht_0_3_MPORT_535_addr] <= pht_0_3_MPORT_535_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_537_en & pht_0_3_MPORT_537_mask) begin
      pht_0_3[pht_0_3_MPORT_537_addr] <= pht_0_3_MPORT_537_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_539_en & pht_0_3_MPORT_539_mask) begin
      pht_0_3[pht_0_3_MPORT_539_addr] <= pht_0_3_MPORT_539_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_541_en & pht_0_3_MPORT_541_mask) begin
      pht_0_3[pht_0_3_MPORT_541_addr] <= pht_0_3_MPORT_541_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_543_en & pht_0_3_MPORT_543_mask) begin
      pht_0_3[pht_0_3_MPORT_543_addr] <= pht_0_3_MPORT_543_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_545_en & pht_0_3_MPORT_545_mask) begin
      pht_0_3[pht_0_3_MPORT_545_addr] <= pht_0_3_MPORT_545_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_547_en & pht_0_3_MPORT_547_mask) begin
      pht_0_3[pht_0_3_MPORT_547_addr] <= pht_0_3_MPORT_547_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_549_en & pht_0_3_MPORT_549_mask) begin
      pht_0_3[pht_0_3_MPORT_549_addr] <= pht_0_3_MPORT_549_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_551_en & pht_0_3_MPORT_551_mask) begin
      pht_0_3[pht_0_3_MPORT_551_addr] <= pht_0_3_MPORT_551_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_553_en & pht_0_3_MPORT_553_mask) begin
      pht_0_3[pht_0_3_MPORT_553_addr] <= pht_0_3_MPORT_553_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_555_en & pht_0_3_MPORT_555_mask) begin
      pht_0_3[pht_0_3_MPORT_555_addr] <= pht_0_3_MPORT_555_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_557_en & pht_0_3_MPORT_557_mask) begin
      pht_0_3[pht_0_3_MPORT_557_addr] <= pht_0_3_MPORT_557_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_3_MPORT_559_en & pht_0_3_MPORT_559_mask) begin
      pht_0_3[pht_0_3_MPORT_559_addr] <= pht_0_3_MPORT_559_data; // @[PatternHistoryTable.scala 26:28]
    end
//     pht_0_3_MPORT_23_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_0_3_MPORT_23_addr_pipe_0 <= io_waddr;
    end
    if (pht_0_4_MPORT_41_en & pht_0_4_MPORT_41_mask) begin
      pht_0_4[pht_0_4_MPORT_41_addr] <= pht_0_4_MPORT_41_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_561_en & pht_0_4_MPORT_561_mask) begin
      pht_0_4[pht_0_4_MPORT_561_addr] <= pht_0_4_MPORT_561_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_563_en & pht_0_4_MPORT_563_mask) begin
      pht_0_4[pht_0_4_MPORT_563_addr] <= pht_0_4_MPORT_563_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_565_en & pht_0_4_MPORT_565_mask) begin
      pht_0_4[pht_0_4_MPORT_565_addr] <= pht_0_4_MPORT_565_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_567_en & pht_0_4_MPORT_567_mask) begin
      pht_0_4[pht_0_4_MPORT_567_addr] <= pht_0_4_MPORT_567_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_569_en & pht_0_4_MPORT_569_mask) begin
      pht_0_4[pht_0_4_MPORT_569_addr] <= pht_0_4_MPORT_569_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_571_en & pht_0_4_MPORT_571_mask) begin
      pht_0_4[pht_0_4_MPORT_571_addr] <= pht_0_4_MPORT_571_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_573_en & pht_0_4_MPORT_573_mask) begin
      pht_0_4[pht_0_4_MPORT_573_addr] <= pht_0_4_MPORT_573_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_575_en & pht_0_4_MPORT_575_mask) begin
      pht_0_4[pht_0_4_MPORT_575_addr] <= pht_0_4_MPORT_575_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_577_en & pht_0_4_MPORT_577_mask) begin
      pht_0_4[pht_0_4_MPORT_577_addr] <= pht_0_4_MPORT_577_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_579_en & pht_0_4_MPORT_579_mask) begin
      pht_0_4[pht_0_4_MPORT_579_addr] <= pht_0_4_MPORT_579_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_581_en & pht_0_4_MPORT_581_mask) begin
      pht_0_4[pht_0_4_MPORT_581_addr] <= pht_0_4_MPORT_581_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_583_en & pht_0_4_MPORT_583_mask) begin
      pht_0_4[pht_0_4_MPORT_583_addr] <= pht_0_4_MPORT_583_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_585_en & pht_0_4_MPORT_585_mask) begin
      pht_0_4[pht_0_4_MPORT_585_addr] <= pht_0_4_MPORT_585_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_587_en & pht_0_4_MPORT_587_mask) begin
      pht_0_4[pht_0_4_MPORT_587_addr] <= pht_0_4_MPORT_587_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_589_en & pht_0_4_MPORT_589_mask) begin
      pht_0_4[pht_0_4_MPORT_589_addr] <= pht_0_4_MPORT_589_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_591_en & pht_0_4_MPORT_591_mask) begin
      pht_0_4[pht_0_4_MPORT_591_addr] <= pht_0_4_MPORT_591_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_593_en & pht_0_4_MPORT_593_mask) begin
      pht_0_4[pht_0_4_MPORT_593_addr] <= pht_0_4_MPORT_593_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_595_en & pht_0_4_MPORT_595_mask) begin
      pht_0_4[pht_0_4_MPORT_595_addr] <= pht_0_4_MPORT_595_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_597_en & pht_0_4_MPORT_597_mask) begin
      pht_0_4[pht_0_4_MPORT_597_addr] <= pht_0_4_MPORT_597_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_599_en & pht_0_4_MPORT_599_mask) begin
      pht_0_4[pht_0_4_MPORT_599_addr] <= pht_0_4_MPORT_599_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_601_en & pht_0_4_MPORT_601_mask) begin
      pht_0_4[pht_0_4_MPORT_601_addr] <= pht_0_4_MPORT_601_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_603_en & pht_0_4_MPORT_603_mask) begin
      pht_0_4[pht_0_4_MPORT_603_addr] <= pht_0_4_MPORT_603_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_605_en & pht_0_4_MPORT_605_mask) begin
      pht_0_4[pht_0_4_MPORT_605_addr] <= pht_0_4_MPORT_605_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_607_en & pht_0_4_MPORT_607_mask) begin
      pht_0_4[pht_0_4_MPORT_607_addr] <= pht_0_4_MPORT_607_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_609_en & pht_0_4_MPORT_609_mask) begin
      pht_0_4[pht_0_4_MPORT_609_addr] <= pht_0_4_MPORT_609_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_611_en & pht_0_4_MPORT_611_mask) begin
      pht_0_4[pht_0_4_MPORT_611_addr] <= pht_0_4_MPORT_611_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_613_en & pht_0_4_MPORT_613_mask) begin
      pht_0_4[pht_0_4_MPORT_613_addr] <= pht_0_4_MPORT_613_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_615_en & pht_0_4_MPORT_615_mask) begin
      pht_0_4[pht_0_4_MPORT_615_addr] <= pht_0_4_MPORT_615_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_617_en & pht_0_4_MPORT_617_mask) begin
      pht_0_4[pht_0_4_MPORT_617_addr] <= pht_0_4_MPORT_617_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_619_en & pht_0_4_MPORT_619_mask) begin
      pht_0_4[pht_0_4_MPORT_619_addr] <= pht_0_4_MPORT_619_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_621_en & pht_0_4_MPORT_621_mask) begin
      pht_0_4[pht_0_4_MPORT_621_addr] <= pht_0_4_MPORT_621_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_623_en & pht_0_4_MPORT_623_mask) begin
      pht_0_4[pht_0_4_MPORT_623_addr] <= pht_0_4_MPORT_623_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_625_en & pht_0_4_MPORT_625_mask) begin
      pht_0_4[pht_0_4_MPORT_625_addr] <= pht_0_4_MPORT_625_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_627_en & pht_0_4_MPORT_627_mask) begin
      pht_0_4[pht_0_4_MPORT_627_addr] <= pht_0_4_MPORT_627_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_629_en & pht_0_4_MPORT_629_mask) begin
      pht_0_4[pht_0_4_MPORT_629_addr] <= pht_0_4_MPORT_629_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_631_en & pht_0_4_MPORT_631_mask) begin
      pht_0_4[pht_0_4_MPORT_631_addr] <= pht_0_4_MPORT_631_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_633_en & pht_0_4_MPORT_633_mask) begin
      pht_0_4[pht_0_4_MPORT_633_addr] <= pht_0_4_MPORT_633_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_635_en & pht_0_4_MPORT_635_mask) begin
      pht_0_4[pht_0_4_MPORT_635_addr] <= pht_0_4_MPORT_635_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_637_en & pht_0_4_MPORT_637_mask) begin
      pht_0_4[pht_0_4_MPORT_637_addr] <= pht_0_4_MPORT_637_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_639_en & pht_0_4_MPORT_639_mask) begin
      pht_0_4[pht_0_4_MPORT_639_addr] <= pht_0_4_MPORT_639_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_641_en & pht_0_4_MPORT_641_mask) begin
      pht_0_4[pht_0_4_MPORT_641_addr] <= pht_0_4_MPORT_641_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_643_en & pht_0_4_MPORT_643_mask) begin
      pht_0_4[pht_0_4_MPORT_643_addr] <= pht_0_4_MPORT_643_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_645_en & pht_0_4_MPORT_645_mask) begin
      pht_0_4[pht_0_4_MPORT_645_addr] <= pht_0_4_MPORT_645_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_647_en & pht_0_4_MPORT_647_mask) begin
      pht_0_4[pht_0_4_MPORT_647_addr] <= pht_0_4_MPORT_647_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_649_en & pht_0_4_MPORT_649_mask) begin
      pht_0_4[pht_0_4_MPORT_649_addr] <= pht_0_4_MPORT_649_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_651_en & pht_0_4_MPORT_651_mask) begin
      pht_0_4[pht_0_4_MPORT_651_addr] <= pht_0_4_MPORT_651_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_653_en & pht_0_4_MPORT_653_mask) begin
      pht_0_4[pht_0_4_MPORT_653_addr] <= pht_0_4_MPORT_653_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_655_en & pht_0_4_MPORT_655_mask) begin
      pht_0_4[pht_0_4_MPORT_655_addr] <= pht_0_4_MPORT_655_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_657_en & pht_0_4_MPORT_657_mask) begin
      pht_0_4[pht_0_4_MPORT_657_addr] <= pht_0_4_MPORT_657_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_659_en & pht_0_4_MPORT_659_mask) begin
      pht_0_4[pht_0_4_MPORT_659_addr] <= pht_0_4_MPORT_659_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_661_en & pht_0_4_MPORT_661_mask) begin
      pht_0_4[pht_0_4_MPORT_661_addr] <= pht_0_4_MPORT_661_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_663_en & pht_0_4_MPORT_663_mask) begin
      pht_0_4[pht_0_4_MPORT_663_addr] <= pht_0_4_MPORT_663_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_665_en & pht_0_4_MPORT_665_mask) begin
      pht_0_4[pht_0_4_MPORT_665_addr] <= pht_0_4_MPORT_665_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_667_en & pht_0_4_MPORT_667_mask) begin
      pht_0_4[pht_0_4_MPORT_667_addr] <= pht_0_4_MPORT_667_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_669_en & pht_0_4_MPORT_669_mask) begin
      pht_0_4[pht_0_4_MPORT_669_addr] <= pht_0_4_MPORT_669_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_671_en & pht_0_4_MPORT_671_mask) begin
      pht_0_4[pht_0_4_MPORT_671_addr] <= pht_0_4_MPORT_671_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_673_en & pht_0_4_MPORT_673_mask) begin
      pht_0_4[pht_0_4_MPORT_673_addr] <= pht_0_4_MPORT_673_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_675_en & pht_0_4_MPORT_675_mask) begin
      pht_0_4[pht_0_4_MPORT_675_addr] <= pht_0_4_MPORT_675_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_677_en & pht_0_4_MPORT_677_mask) begin
      pht_0_4[pht_0_4_MPORT_677_addr] <= pht_0_4_MPORT_677_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_679_en & pht_0_4_MPORT_679_mask) begin
      pht_0_4[pht_0_4_MPORT_679_addr] <= pht_0_4_MPORT_679_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_681_en & pht_0_4_MPORT_681_mask) begin
      pht_0_4[pht_0_4_MPORT_681_addr] <= pht_0_4_MPORT_681_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_683_en & pht_0_4_MPORT_683_mask) begin
      pht_0_4[pht_0_4_MPORT_683_addr] <= pht_0_4_MPORT_683_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_685_en & pht_0_4_MPORT_685_mask) begin
      pht_0_4[pht_0_4_MPORT_685_addr] <= pht_0_4_MPORT_685_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_4_MPORT_687_en & pht_0_4_MPORT_687_mask) begin
      pht_0_4[pht_0_4_MPORT_687_addr] <= pht_0_4_MPORT_687_data; // @[PatternHistoryTable.scala 26:28]
    end
//     pht_0_4_MPORT_25_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_0_4_MPORT_25_addr_pipe_0 <= io_waddr;
    end
    if (pht_0_5_MPORT_43_en & pht_0_5_MPORT_43_mask) begin
      pht_0_5[pht_0_5_MPORT_43_addr] <= pht_0_5_MPORT_43_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_689_en & pht_0_5_MPORT_689_mask) begin
      pht_0_5[pht_0_5_MPORT_689_addr] <= pht_0_5_MPORT_689_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_691_en & pht_0_5_MPORT_691_mask) begin
      pht_0_5[pht_0_5_MPORT_691_addr] <= pht_0_5_MPORT_691_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_693_en & pht_0_5_MPORT_693_mask) begin
      pht_0_5[pht_0_5_MPORT_693_addr] <= pht_0_5_MPORT_693_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_695_en & pht_0_5_MPORT_695_mask) begin
      pht_0_5[pht_0_5_MPORT_695_addr] <= pht_0_5_MPORT_695_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_697_en & pht_0_5_MPORT_697_mask) begin
      pht_0_5[pht_0_5_MPORT_697_addr] <= pht_0_5_MPORT_697_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_699_en & pht_0_5_MPORT_699_mask) begin
      pht_0_5[pht_0_5_MPORT_699_addr] <= pht_0_5_MPORT_699_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_701_en & pht_0_5_MPORT_701_mask) begin
      pht_0_5[pht_0_5_MPORT_701_addr] <= pht_0_5_MPORT_701_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_703_en & pht_0_5_MPORT_703_mask) begin
      pht_0_5[pht_0_5_MPORT_703_addr] <= pht_0_5_MPORT_703_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_705_en & pht_0_5_MPORT_705_mask) begin
      pht_0_5[pht_0_5_MPORT_705_addr] <= pht_0_5_MPORT_705_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_707_en & pht_0_5_MPORT_707_mask) begin
      pht_0_5[pht_0_5_MPORT_707_addr] <= pht_0_5_MPORT_707_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_709_en & pht_0_5_MPORT_709_mask) begin
      pht_0_5[pht_0_5_MPORT_709_addr] <= pht_0_5_MPORT_709_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_711_en & pht_0_5_MPORT_711_mask) begin
      pht_0_5[pht_0_5_MPORT_711_addr] <= pht_0_5_MPORT_711_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_713_en & pht_0_5_MPORT_713_mask) begin
      pht_0_5[pht_0_5_MPORT_713_addr] <= pht_0_5_MPORT_713_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_715_en & pht_0_5_MPORT_715_mask) begin
      pht_0_5[pht_0_5_MPORT_715_addr] <= pht_0_5_MPORT_715_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_717_en & pht_0_5_MPORT_717_mask) begin
      pht_0_5[pht_0_5_MPORT_717_addr] <= pht_0_5_MPORT_717_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_719_en & pht_0_5_MPORT_719_mask) begin
      pht_0_5[pht_0_5_MPORT_719_addr] <= pht_0_5_MPORT_719_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_721_en & pht_0_5_MPORT_721_mask) begin
      pht_0_5[pht_0_5_MPORT_721_addr] <= pht_0_5_MPORT_721_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_723_en & pht_0_5_MPORT_723_mask) begin
      pht_0_5[pht_0_5_MPORT_723_addr] <= pht_0_5_MPORT_723_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_725_en & pht_0_5_MPORT_725_mask) begin
      pht_0_5[pht_0_5_MPORT_725_addr] <= pht_0_5_MPORT_725_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_727_en & pht_0_5_MPORT_727_mask) begin
      pht_0_5[pht_0_5_MPORT_727_addr] <= pht_0_5_MPORT_727_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_729_en & pht_0_5_MPORT_729_mask) begin
      pht_0_5[pht_0_5_MPORT_729_addr] <= pht_0_5_MPORT_729_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_731_en & pht_0_5_MPORT_731_mask) begin
      pht_0_5[pht_0_5_MPORT_731_addr] <= pht_0_5_MPORT_731_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_733_en & pht_0_5_MPORT_733_mask) begin
      pht_0_5[pht_0_5_MPORT_733_addr] <= pht_0_5_MPORT_733_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_735_en & pht_0_5_MPORT_735_mask) begin
      pht_0_5[pht_0_5_MPORT_735_addr] <= pht_0_5_MPORT_735_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_737_en & pht_0_5_MPORT_737_mask) begin
      pht_0_5[pht_0_5_MPORT_737_addr] <= pht_0_5_MPORT_737_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_739_en & pht_0_5_MPORT_739_mask) begin
      pht_0_5[pht_0_5_MPORT_739_addr] <= pht_0_5_MPORT_739_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_741_en & pht_0_5_MPORT_741_mask) begin
      pht_0_5[pht_0_5_MPORT_741_addr] <= pht_0_5_MPORT_741_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_743_en & pht_0_5_MPORT_743_mask) begin
      pht_0_5[pht_0_5_MPORT_743_addr] <= pht_0_5_MPORT_743_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_745_en & pht_0_5_MPORT_745_mask) begin
      pht_0_5[pht_0_5_MPORT_745_addr] <= pht_0_5_MPORT_745_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_747_en & pht_0_5_MPORT_747_mask) begin
      pht_0_5[pht_0_5_MPORT_747_addr] <= pht_0_5_MPORT_747_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_749_en & pht_0_5_MPORT_749_mask) begin
      pht_0_5[pht_0_5_MPORT_749_addr] <= pht_0_5_MPORT_749_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_751_en & pht_0_5_MPORT_751_mask) begin
      pht_0_5[pht_0_5_MPORT_751_addr] <= pht_0_5_MPORT_751_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_753_en & pht_0_5_MPORT_753_mask) begin
      pht_0_5[pht_0_5_MPORT_753_addr] <= pht_0_5_MPORT_753_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_755_en & pht_0_5_MPORT_755_mask) begin
      pht_0_5[pht_0_5_MPORT_755_addr] <= pht_0_5_MPORT_755_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_757_en & pht_0_5_MPORT_757_mask) begin
      pht_0_5[pht_0_5_MPORT_757_addr] <= pht_0_5_MPORT_757_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_759_en & pht_0_5_MPORT_759_mask) begin
      pht_0_5[pht_0_5_MPORT_759_addr] <= pht_0_5_MPORT_759_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_761_en & pht_0_5_MPORT_761_mask) begin
      pht_0_5[pht_0_5_MPORT_761_addr] <= pht_0_5_MPORT_761_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_763_en & pht_0_5_MPORT_763_mask) begin
      pht_0_5[pht_0_5_MPORT_763_addr] <= pht_0_5_MPORT_763_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_765_en & pht_0_5_MPORT_765_mask) begin
      pht_0_5[pht_0_5_MPORT_765_addr] <= pht_0_5_MPORT_765_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_767_en & pht_0_5_MPORT_767_mask) begin
      pht_0_5[pht_0_5_MPORT_767_addr] <= pht_0_5_MPORT_767_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_769_en & pht_0_5_MPORT_769_mask) begin
      pht_0_5[pht_0_5_MPORT_769_addr] <= pht_0_5_MPORT_769_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_771_en & pht_0_5_MPORT_771_mask) begin
      pht_0_5[pht_0_5_MPORT_771_addr] <= pht_0_5_MPORT_771_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_773_en & pht_0_5_MPORT_773_mask) begin
      pht_0_5[pht_0_5_MPORT_773_addr] <= pht_0_5_MPORT_773_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_775_en & pht_0_5_MPORT_775_mask) begin
      pht_0_5[pht_0_5_MPORT_775_addr] <= pht_0_5_MPORT_775_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_777_en & pht_0_5_MPORT_777_mask) begin
      pht_0_5[pht_0_5_MPORT_777_addr] <= pht_0_5_MPORT_777_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_779_en & pht_0_5_MPORT_779_mask) begin
      pht_0_5[pht_0_5_MPORT_779_addr] <= pht_0_5_MPORT_779_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_781_en & pht_0_5_MPORT_781_mask) begin
      pht_0_5[pht_0_5_MPORT_781_addr] <= pht_0_5_MPORT_781_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_783_en & pht_0_5_MPORT_783_mask) begin
      pht_0_5[pht_0_5_MPORT_783_addr] <= pht_0_5_MPORT_783_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_785_en & pht_0_5_MPORT_785_mask) begin
      pht_0_5[pht_0_5_MPORT_785_addr] <= pht_0_5_MPORT_785_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_787_en & pht_0_5_MPORT_787_mask) begin
      pht_0_5[pht_0_5_MPORT_787_addr] <= pht_0_5_MPORT_787_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_789_en & pht_0_5_MPORT_789_mask) begin
      pht_0_5[pht_0_5_MPORT_789_addr] <= pht_0_5_MPORT_789_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_791_en & pht_0_5_MPORT_791_mask) begin
      pht_0_5[pht_0_5_MPORT_791_addr] <= pht_0_5_MPORT_791_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_793_en & pht_0_5_MPORT_793_mask) begin
      pht_0_5[pht_0_5_MPORT_793_addr] <= pht_0_5_MPORT_793_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_795_en & pht_0_5_MPORT_795_mask) begin
      pht_0_5[pht_0_5_MPORT_795_addr] <= pht_0_5_MPORT_795_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_797_en & pht_0_5_MPORT_797_mask) begin
      pht_0_5[pht_0_5_MPORT_797_addr] <= pht_0_5_MPORT_797_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_799_en & pht_0_5_MPORT_799_mask) begin
      pht_0_5[pht_0_5_MPORT_799_addr] <= pht_0_5_MPORT_799_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_801_en & pht_0_5_MPORT_801_mask) begin
      pht_0_5[pht_0_5_MPORT_801_addr] <= pht_0_5_MPORT_801_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_803_en & pht_0_5_MPORT_803_mask) begin
      pht_0_5[pht_0_5_MPORT_803_addr] <= pht_0_5_MPORT_803_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_805_en & pht_0_5_MPORT_805_mask) begin
      pht_0_5[pht_0_5_MPORT_805_addr] <= pht_0_5_MPORT_805_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_807_en & pht_0_5_MPORT_807_mask) begin
      pht_0_5[pht_0_5_MPORT_807_addr] <= pht_0_5_MPORT_807_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_809_en & pht_0_5_MPORT_809_mask) begin
      pht_0_5[pht_0_5_MPORT_809_addr] <= pht_0_5_MPORT_809_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_811_en & pht_0_5_MPORT_811_mask) begin
      pht_0_5[pht_0_5_MPORT_811_addr] <= pht_0_5_MPORT_811_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_813_en & pht_0_5_MPORT_813_mask) begin
      pht_0_5[pht_0_5_MPORT_813_addr] <= pht_0_5_MPORT_813_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_5_MPORT_815_en & pht_0_5_MPORT_815_mask) begin
      pht_0_5[pht_0_5_MPORT_815_addr] <= pht_0_5_MPORT_815_data; // @[PatternHistoryTable.scala 26:28]
    end
//     pht_0_5_MPORT_27_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_0_5_MPORT_27_addr_pipe_0 <= io_waddr;
    end
    if (pht_0_6_MPORT_45_en & pht_0_6_MPORT_45_mask) begin
      pht_0_6[pht_0_6_MPORT_45_addr] <= pht_0_6_MPORT_45_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_817_en & pht_0_6_MPORT_817_mask) begin
      pht_0_6[pht_0_6_MPORT_817_addr] <= pht_0_6_MPORT_817_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_819_en & pht_0_6_MPORT_819_mask) begin
      pht_0_6[pht_0_6_MPORT_819_addr] <= pht_0_6_MPORT_819_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_821_en & pht_0_6_MPORT_821_mask) begin
      pht_0_6[pht_0_6_MPORT_821_addr] <= pht_0_6_MPORT_821_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_823_en & pht_0_6_MPORT_823_mask) begin
      pht_0_6[pht_0_6_MPORT_823_addr] <= pht_0_6_MPORT_823_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_825_en & pht_0_6_MPORT_825_mask) begin
      pht_0_6[pht_0_6_MPORT_825_addr] <= pht_0_6_MPORT_825_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_827_en & pht_0_6_MPORT_827_mask) begin
      pht_0_6[pht_0_6_MPORT_827_addr] <= pht_0_6_MPORT_827_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_829_en & pht_0_6_MPORT_829_mask) begin
      pht_0_6[pht_0_6_MPORT_829_addr] <= pht_0_6_MPORT_829_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_831_en & pht_0_6_MPORT_831_mask) begin
      pht_0_6[pht_0_6_MPORT_831_addr] <= pht_0_6_MPORT_831_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_833_en & pht_0_6_MPORT_833_mask) begin
      pht_0_6[pht_0_6_MPORT_833_addr] <= pht_0_6_MPORT_833_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_835_en & pht_0_6_MPORT_835_mask) begin
      pht_0_6[pht_0_6_MPORT_835_addr] <= pht_0_6_MPORT_835_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_837_en & pht_0_6_MPORT_837_mask) begin
      pht_0_6[pht_0_6_MPORT_837_addr] <= pht_0_6_MPORT_837_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_839_en & pht_0_6_MPORT_839_mask) begin
      pht_0_6[pht_0_6_MPORT_839_addr] <= pht_0_6_MPORT_839_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_841_en & pht_0_6_MPORT_841_mask) begin
      pht_0_6[pht_0_6_MPORT_841_addr] <= pht_0_6_MPORT_841_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_843_en & pht_0_6_MPORT_843_mask) begin
      pht_0_6[pht_0_6_MPORT_843_addr] <= pht_0_6_MPORT_843_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_845_en & pht_0_6_MPORT_845_mask) begin
      pht_0_6[pht_0_6_MPORT_845_addr] <= pht_0_6_MPORT_845_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_847_en & pht_0_6_MPORT_847_mask) begin
      pht_0_6[pht_0_6_MPORT_847_addr] <= pht_0_6_MPORT_847_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_849_en & pht_0_6_MPORT_849_mask) begin
      pht_0_6[pht_0_6_MPORT_849_addr] <= pht_0_6_MPORT_849_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_851_en & pht_0_6_MPORT_851_mask) begin
      pht_0_6[pht_0_6_MPORT_851_addr] <= pht_0_6_MPORT_851_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_853_en & pht_0_6_MPORT_853_mask) begin
      pht_0_6[pht_0_6_MPORT_853_addr] <= pht_0_6_MPORT_853_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_855_en & pht_0_6_MPORT_855_mask) begin
      pht_0_6[pht_0_6_MPORT_855_addr] <= pht_0_6_MPORT_855_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_857_en & pht_0_6_MPORT_857_mask) begin
      pht_0_6[pht_0_6_MPORT_857_addr] <= pht_0_6_MPORT_857_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_859_en & pht_0_6_MPORT_859_mask) begin
      pht_0_6[pht_0_6_MPORT_859_addr] <= pht_0_6_MPORT_859_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_861_en & pht_0_6_MPORT_861_mask) begin
      pht_0_6[pht_0_6_MPORT_861_addr] <= pht_0_6_MPORT_861_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_863_en & pht_0_6_MPORT_863_mask) begin
      pht_0_6[pht_0_6_MPORT_863_addr] <= pht_0_6_MPORT_863_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_865_en & pht_0_6_MPORT_865_mask) begin
      pht_0_6[pht_0_6_MPORT_865_addr] <= pht_0_6_MPORT_865_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_867_en & pht_0_6_MPORT_867_mask) begin
      pht_0_6[pht_0_6_MPORT_867_addr] <= pht_0_6_MPORT_867_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_869_en & pht_0_6_MPORT_869_mask) begin
      pht_0_6[pht_0_6_MPORT_869_addr] <= pht_0_6_MPORT_869_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_871_en & pht_0_6_MPORT_871_mask) begin
      pht_0_6[pht_0_6_MPORT_871_addr] <= pht_0_6_MPORT_871_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_873_en & pht_0_6_MPORT_873_mask) begin
      pht_0_6[pht_0_6_MPORT_873_addr] <= pht_0_6_MPORT_873_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_875_en & pht_0_6_MPORT_875_mask) begin
      pht_0_6[pht_0_6_MPORT_875_addr] <= pht_0_6_MPORT_875_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_877_en & pht_0_6_MPORT_877_mask) begin
      pht_0_6[pht_0_6_MPORT_877_addr] <= pht_0_6_MPORT_877_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_879_en & pht_0_6_MPORT_879_mask) begin
      pht_0_6[pht_0_6_MPORT_879_addr] <= pht_0_6_MPORT_879_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_881_en & pht_0_6_MPORT_881_mask) begin
      pht_0_6[pht_0_6_MPORT_881_addr] <= pht_0_6_MPORT_881_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_883_en & pht_0_6_MPORT_883_mask) begin
      pht_0_6[pht_0_6_MPORT_883_addr] <= pht_0_6_MPORT_883_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_885_en & pht_0_6_MPORT_885_mask) begin
      pht_0_6[pht_0_6_MPORT_885_addr] <= pht_0_6_MPORT_885_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_887_en & pht_0_6_MPORT_887_mask) begin
      pht_0_6[pht_0_6_MPORT_887_addr] <= pht_0_6_MPORT_887_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_889_en & pht_0_6_MPORT_889_mask) begin
      pht_0_6[pht_0_6_MPORT_889_addr] <= pht_0_6_MPORT_889_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_891_en & pht_0_6_MPORT_891_mask) begin
      pht_0_6[pht_0_6_MPORT_891_addr] <= pht_0_6_MPORT_891_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_893_en & pht_0_6_MPORT_893_mask) begin
      pht_0_6[pht_0_6_MPORT_893_addr] <= pht_0_6_MPORT_893_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_895_en & pht_0_6_MPORT_895_mask) begin
      pht_0_6[pht_0_6_MPORT_895_addr] <= pht_0_6_MPORT_895_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_897_en & pht_0_6_MPORT_897_mask) begin
      pht_0_6[pht_0_6_MPORT_897_addr] <= pht_0_6_MPORT_897_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_899_en & pht_0_6_MPORT_899_mask) begin
      pht_0_6[pht_0_6_MPORT_899_addr] <= pht_0_6_MPORT_899_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_901_en & pht_0_6_MPORT_901_mask) begin
      pht_0_6[pht_0_6_MPORT_901_addr] <= pht_0_6_MPORT_901_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_903_en & pht_0_6_MPORT_903_mask) begin
      pht_0_6[pht_0_6_MPORT_903_addr] <= pht_0_6_MPORT_903_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_905_en & pht_0_6_MPORT_905_mask) begin
      pht_0_6[pht_0_6_MPORT_905_addr] <= pht_0_6_MPORT_905_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_907_en & pht_0_6_MPORT_907_mask) begin
      pht_0_6[pht_0_6_MPORT_907_addr] <= pht_0_6_MPORT_907_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_909_en & pht_0_6_MPORT_909_mask) begin
      pht_0_6[pht_0_6_MPORT_909_addr] <= pht_0_6_MPORT_909_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_911_en & pht_0_6_MPORT_911_mask) begin
      pht_0_6[pht_0_6_MPORT_911_addr] <= pht_0_6_MPORT_911_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_913_en & pht_0_6_MPORT_913_mask) begin
      pht_0_6[pht_0_6_MPORT_913_addr] <= pht_0_6_MPORT_913_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_915_en & pht_0_6_MPORT_915_mask) begin
      pht_0_6[pht_0_6_MPORT_915_addr] <= pht_0_6_MPORT_915_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_917_en & pht_0_6_MPORT_917_mask) begin
      pht_0_6[pht_0_6_MPORT_917_addr] <= pht_0_6_MPORT_917_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_919_en & pht_0_6_MPORT_919_mask) begin
      pht_0_6[pht_0_6_MPORT_919_addr] <= pht_0_6_MPORT_919_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_921_en & pht_0_6_MPORT_921_mask) begin
      pht_0_6[pht_0_6_MPORT_921_addr] <= pht_0_6_MPORT_921_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_923_en & pht_0_6_MPORT_923_mask) begin
      pht_0_6[pht_0_6_MPORT_923_addr] <= pht_0_6_MPORT_923_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_925_en & pht_0_6_MPORT_925_mask) begin
      pht_0_6[pht_0_6_MPORT_925_addr] <= pht_0_6_MPORT_925_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_927_en & pht_0_6_MPORT_927_mask) begin
      pht_0_6[pht_0_6_MPORT_927_addr] <= pht_0_6_MPORT_927_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_929_en & pht_0_6_MPORT_929_mask) begin
      pht_0_6[pht_0_6_MPORT_929_addr] <= pht_0_6_MPORT_929_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_931_en & pht_0_6_MPORT_931_mask) begin
      pht_0_6[pht_0_6_MPORT_931_addr] <= pht_0_6_MPORT_931_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_933_en & pht_0_6_MPORT_933_mask) begin
      pht_0_6[pht_0_6_MPORT_933_addr] <= pht_0_6_MPORT_933_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_935_en & pht_0_6_MPORT_935_mask) begin
      pht_0_6[pht_0_6_MPORT_935_addr] <= pht_0_6_MPORT_935_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_937_en & pht_0_6_MPORT_937_mask) begin
      pht_0_6[pht_0_6_MPORT_937_addr] <= pht_0_6_MPORT_937_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_939_en & pht_0_6_MPORT_939_mask) begin
      pht_0_6[pht_0_6_MPORT_939_addr] <= pht_0_6_MPORT_939_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_941_en & pht_0_6_MPORT_941_mask) begin
      pht_0_6[pht_0_6_MPORT_941_addr] <= pht_0_6_MPORT_941_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_6_MPORT_943_en & pht_0_6_MPORT_943_mask) begin
      pht_0_6[pht_0_6_MPORT_943_addr] <= pht_0_6_MPORT_943_data; // @[PatternHistoryTable.scala 26:28]
    end
//     pht_0_6_MPORT_29_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_0_6_MPORT_29_addr_pipe_0 <= io_waddr;
    end
    if (pht_0_7_MPORT_47_en & pht_0_7_MPORT_47_mask) begin
      pht_0_7[pht_0_7_MPORT_47_addr] <= pht_0_7_MPORT_47_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_945_en & pht_0_7_MPORT_945_mask) begin
      pht_0_7[pht_0_7_MPORT_945_addr] <= pht_0_7_MPORT_945_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_947_en & pht_0_7_MPORT_947_mask) begin
      pht_0_7[pht_0_7_MPORT_947_addr] <= pht_0_7_MPORT_947_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_949_en & pht_0_7_MPORT_949_mask) begin
      pht_0_7[pht_0_7_MPORT_949_addr] <= pht_0_7_MPORT_949_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_951_en & pht_0_7_MPORT_951_mask) begin
      pht_0_7[pht_0_7_MPORT_951_addr] <= pht_0_7_MPORT_951_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_953_en & pht_0_7_MPORT_953_mask) begin
      pht_0_7[pht_0_7_MPORT_953_addr] <= pht_0_7_MPORT_953_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_955_en & pht_0_7_MPORT_955_mask) begin
      pht_0_7[pht_0_7_MPORT_955_addr] <= pht_0_7_MPORT_955_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_957_en & pht_0_7_MPORT_957_mask) begin
      pht_0_7[pht_0_7_MPORT_957_addr] <= pht_0_7_MPORT_957_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_959_en & pht_0_7_MPORT_959_mask) begin
      pht_0_7[pht_0_7_MPORT_959_addr] <= pht_0_7_MPORT_959_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_961_en & pht_0_7_MPORT_961_mask) begin
      pht_0_7[pht_0_7_MPORT_961_addr] <= pht_0_7_MPORT_961_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_963_en & pht_0_7_MPORT_963_mask) begin
      pht_0_7[pht_0_7_MPORT_963_addr] <= pht_0_7_MPORT_963_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_965_en & pht_0_7_MPORT_965_mask) begin
      pht_0_7[pht_0_7_MPORT_965_addr] <= pht_0_7_MPORT_965_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_967_en & pht_0_7_MPORT_967_mask) begin
      pht_0_7[pht_0_7_MPORT_967_addr] <= pht_0_7_MPORT_967_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_969_en & pht_0_7_MPORT_969_mask) begin
      pht_0_7[pht_0_7_MPORT_969_addr] <= pht_0_7_MPORT_969_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_971_en & pht_0_7_MPORT_971_mask) begin
      pht_0_7[pht_0_7_MPORT_971_addr] <= pht_0_7_MPORT_971_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_973_en & pht_0_7_MPORT_973_mask) begin
      pht_0_7[pht_0_7_MPORT_973_addr] <= pht_0_7_MPORT_973_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_975_en & pht_0_7_MPORT_975_mask) begin
      pht_0_7[pht_0_7_MPORT_975_addr] <= pht_0_7_MPORT_975_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_977_en & pht_0_7_MPORT_977_mask) begin
      pht_0_7[pht_0_7_MPORT_977_addr] <= pht_0_7_MPORT_977_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_979_en & pht_0_7_MPORT_979_mask) begin
      pht_0_7[pht_0_7_MPORT_979_addr] <= pht_0_7_MPORT_979_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_981_en & pht_0_7_MPORT_981_mask) begin
      pht_0_7[pht_0_7_MPORT_981_addr] <= pht_0_7_MPORT_981_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_983_en & pht_0_7_MPORT_983_mask) begin
      pht_0_7[pht_0_7_MPORT_983_addr] <= pht_0_7_MPORT_983_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_985_en & pht_0_7_MPORT_985_mask) begin
      pht_0_7[pht_0_7_MPORT_985_addr] <= pht_0_7_MPORT_985_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_987_en & pht_0_7_MPORT_987_mask) begin
      pht_0_7[pht_0_7_MPORT_987_addr] <= pht_0_7_MPORT_987_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_989_en & pht_0_7_MPORT_989_mask) begin
      pht_0_7[pht_0_7_MPORT_989_addr] <= pht_0_7_MPORT_989_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_991_en & pht_0_7_MPORT_991_mask) begin
      pht_0_7[pht_0_7_MPORT_991_addr] <= pht_0_7_MPORT_991_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_993_en & pht_0_7_MPORT_993_mask) begin
      pht_0_7[pht_0_7_MPORT_993_addr] <= pht_0_7_MPORT_993_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_995_en & pht_0_7_MPORT_995_mask) begin
      pht_0_7[pht_0_7_MPORT_995_addr] <= pht_0_7_MPORT_995_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_997_en & pht_0_7_MPORT_997_mask) begin
      pht_0_7[pht_0_7_MPORT_997_addr] <= pht_0_7_MPORT_997_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_999_en & pht_0_7_MPORT_999_mask) begin
      pht_0_7[pht_0_7_MPORT_999_addr] <= pht_0_7_MPORT_999_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1001_en & pht_0_7_MPORT_1001_mask) begin
      pht_0_7[pht_0_7_MPORT_1001_addr] <= pht_0_7_MPORT_1001_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1003_en & pht_0_7_MPORT_1003_mask) begin
      pht_0_7[pht_0_7_MPORT_1003_addr] <= pht_0_7_MPORT_1003_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1005_en & pht_0_7_MPORT_1005_mask) begin
      pht_0_7[pht_0_7_MPORT_1005_addr] <= pht_0_7_MPORT_1005_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1007_en & pht_0_7_MPORT_1007_mask) begin
      pht_0_7[pht_0_7_MPORT_1007_addr] <= pht_0_7_MPORT_1007_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1009_en & pht_0_7_MPORT_1009_mask) begin
      pht_0_7[pht_0_7_MPORT_1009_addr] <= pht_0_7_MPORT_1009_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1011_en & pht_0_7_MPORT_1011_mask) begin
      pht_0_7[pht_0_7_MPORT_1011_addr] <= pht_0_7_MPORT_1011_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1013_en & pht_0_7_MPORT_1013_mask) begin
      pht_0_7[pht_0_7_MPORT_1013_addr] <= pht_0_7_MPORT_1013_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1015_en & pht_0_7_MPORT_1015_mask) begin
      pht_0_7[pht_0_7_MPORT_1015_addr] <= pht_0_7_MPORT_1015_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1017_en & pht_0_7_MPORT_1017_mask) begin
      pht_0_7[pht_0_7_MPORT_1017_addr] <= pht_0_7_MPORT_1017_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1019_en & pht_0_7_MPORT_1019_mask) begin
      pht_0_7[pht_0_7_MPORT_1019_addr] <= pht_0_7_MPORT_1019_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1021_en & pht_0_7_MPORT_1021_mask) begin
      pht_0_7[pht_0_7_MPORT_1021_addr] <= pht_0_7_MPORT_1021_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1023_en & pht_0_7_MPORT_1023_mask) begin
      pht_0_7[pht_0_7_MPORT_1023_addr] <= pht_0_7_MPORT_1023_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1025_en & pht_0_7_MPORT_1025_mask) begin
      pht_0_7[pht_0_7_MPORT_1025_addr] <= pht_0_7_MPORT_1025_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1027_en & pht_0_7_MPORT_1027_mask) begin
      pht_0_7[pht_0_7_MPORT_1027_addr] <= pht_0_7_MPORT_1027_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1029_en & pht_0_7_MPORT_1029_mask) begin
      pht_0_7[pht_0_7_MPORT_1029_addr] <= pht_0_7_MPORT_1029_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1031_en & pht_0_7_MPORT_1031_mask) begin
      pht_0_7[pht_0_7_MPORT_1031_addr] <= pht_0_7_MPORT_1031_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1033_en & pht_0_7_MPORT_1033_mask) begin
      pht_0_7[pht_0_7_MPORT_1033_addr] <= pht_0_7_MPORT_1033_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1035_en & pht_0_7_MPORT_1035_mask) begin
      pht_0_7[pht_0_7_MPORT_1035_addr] <= pht_0_7_MPORT_1035_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1037_en & pht_0_7_MPORT_1037_mask) begin
      pht_0_7[pht_0_7_MPORT_1037_addr] <= pht_0_7_MPORT_1037_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1039_en & pht_0_7_MPORT_1039_mask) begin
      pht_0_7[pht_0_7_MPORT_1039_addr] <= pht_0_7_MPORT_1039_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1041_en & pht_0_7_MPORT_1041_mask) begin
      pht_0_7[pht_0_7_MPORT_1041_addr] <= pht_0_7_MPORT_1041_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1043_en & pht_0_7_MPORT_1043_mask) begin
      pht_0_7[pht_0_7_MPORT_1043_addr] <= pht_0_7_MPORT_1043_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1045_en & pht_0_7_MPORT_1045_mask) begin
      pht_0_7[pht_0_7_MPORT_1045_addr] <= pht_0_7_MPORT_1045_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1047_en & pht_0_7_MPORT_1047_mask) begin
      pht_0_7[pht_0_7_MPORT_1047_addr] <= pht_0_7_MPORT_1047_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1049_en & pht_0_7_MPORT_1049_mask) begin
      pht_0_7[pht_0_7_MPORT_1049_addr] <= pht_0_7_MPORT_1049_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1051_en & pht_0_7_MPORT_1051_mask) begin
      pht_0_7[pht_0_7_MPORT_1051_addr] <= pht_0_7_MPORT_1051_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1053_en & pht_0_7_MPORT_1053_mask) begin
      pht_0_7[pht_0_7_MPORT_1053_addr] <= pht_0_7_MPORT_1053_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1055_en & pht_0_7_MPORT_1055_mask) begin
      pht_0_7[pht_0_7_MPORT_1055_addr] <= pht_0_7_MPORT_1055_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1057_en & pht_0_7_MPORT_1057_mask) begin
      pht_0_7[pht_0_7_MPORT_1057_addr] <= pht_0_7_MPORT_1057_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1059_en & pht_0_7_MPORT_1059_mask) begin
      pht_0_7[pht_0_7_MPORT_1059_addr] <= pht_0_7_MPORT_1059_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1061_en & pht_0_7_MPORT_1061_mask) begin
      pht_0_7[pht_0_7_MPORT_1061_addr] <= pht_0_7_MPORT_1061_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1063_en & pht_0_7_MPORT_1063_mask) begin
      pht_0_7[pht_0_7_MPORT_1063_addr] <= pht_0_7_MPORT_1063_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1065_en & pht_0_7_MPORT_1065_mask) begin
      pht_0_7[pht_0_7_MPORT_1065_addr] <= pht_0_7_MPORT_1065_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1067_en & pht_0_7_MPORT_1067_mask) begin
      pht_0_7[pht_0_7_MPORT_1067_addr] <= pht_0_7_MPORT_1067_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1069_en & pht_0_7_MPORT_1069_mask) begin
      pht_0_7[pht_0_7_MPORT_1069_addr] <= pht_0_7_MPORT_1069_data; // @[PatternHistoryTable.scala 26:28]
    end
    if (pht_0_7_MPORT_1071_en & pht_0_7_MPORT_1071_mask) begin
      pht_0_7[pht_0_7_MPORT_1071_addr] <= pht_0_7_MPORT_1071_data; // @[PatternHistoryTable.scala 26:28]
    end
//     pht_0_7_MPORT_31_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      pht_0_7_MPORT_31_addr_pipe_0 <= io_waddr;
    end
    REG <= io_rindex_0; // @[PatternHistoryTable.scala 42:20]
    REG_1 <= io_rindex_0; // @[PatternHistoryTable.scala 42:20]
    REG_2 <= io_rindex_0; // @[PatternHistoryTable.scala 42:20]
    REG_3 <= io_rindex_0; // @[PatternHistoryTable.scala 42:20]
    REG_4 <= io_rindex_0; // @[PatternHistoryTable.scala 42:20]
    REG_5 <= io_rindex_0; // @[PatternHistoryTable.scala 42:20]
    REG_6 <= io_rindex_0; // @[PatternHistoryTable.scala 42:20]
    REG_7 <= io_rindex_0; // @[PatternHistoryTable.scala 42:20]
    REG_8 <= io_rindex_1; // @[PatternHistoryTable.scala 42:20]
    REG_9 <= io_rindex_1; // @[PatternHistoryTable.scala 42:20]
    REG_10 <= io_rindex_1; // @[PatternHistoryTable.scala 42:20]
    REG_11 <= io_rindex_1; // @[PatternHistoryTable.scala 42:20]
    REG_12 <= io_rindex_1; // @[PatternHistoryTable.scala 42:20]
    REG_13 <= io_rindex_1; // @[PatternHistoryTable.scala 42:20]
    REG_14 <= io_rindex_1; // @[PatternHistoryTable.scala 42:20]
    REG_15 <= io_rindex_1; // @[PatternHistoryTable.scala 42:20]
    REG_16 <= io_wen; // @[PatternHistoryTable.scala 59:16]
    REG_17 <= io_windex; // @[PatternHistoryTable.scala 61:20]
    REG_18 <= io_windex; // @[PatternHistoryTable.scala 61:20]
    REG_19 <= io_windex; // @[PatternHistoryTable.scala 61:20]
    REG_20 <= io_windex; // @[PatternHistoryTable.scala 61:20]
    REG_21 <= io_windex; // @[PatternHistoryTable.scala 61:20]
    REG_22 <= io_windex; // @[PatternHistoryTable.scala 61:20]
    REG_23 <= io_windex; // @[PatternHistoryTable.scala 61:20]
    REG_24 <= io_windex; // @[PatternHistoryTable.scala 61:20]
    REG_25 <= io_wjmp; // @[PatternHistoryTable.scala 67:23]
    REG_26 <= io_wjmp; // @[PatternHistoryTable.scala 68:23]
    REG_27 <= io_wjmp; // @[PatternHistoryTable.scala 69:23]
    REG_28 <= io_wjmp; // @[PatternHistoryTable.scala 70:23]
    REG_29 <= io_wen; // @[PatternHistoryTable.scala 72:16]
    REG_30 <= io_windex == 3'h0; // @[PatternHistoryTable.scala 74:31]
    REG_31 <= io_waddr; // @[PatternHistoryTable.scala 75:31]
    REG_32 <= io_waddr; // @[PatternHistoryTable.scala 76:31]
    REG_33 <= io_windex == 3'h1; // @[PatternHistoryTable.scala 74:31]
    REG_34 <= io_waddr; // @[PatternHistoryTable.scala 75:31]
    REG_35 <= io_waddr; // @[PatternHistoryTable.scala 76:31]
    REG_36 <= io_windex == 3'h2; // @[PatternHistoryTable.scala 74:31]
    REG_37 <= io_waddr; // @[PatternHistoryTable.scala 75:31]
    REG_38 <= io_waddr; // @[PatternHistoryTable.scala 76:31]
    REG_39 <= io_windex == 3'h3; // @[PatternHistoryTable.scala 74:31]
    REG_40 <= io_waddr; // @[PatternHistoryTable.scala 75:31]
    REG_41 <= io_waddr; // @[PatternHistoryTable.scala 76:31]
    REG_42 <= io_windex == 3'h4; // @[PatternHistoryTable.scala 74:31]
    REG_43 <= io_waddr; // @[PatternHistoryTable.scala 75:31]
    REG_44 <= io_waddr; // @[PatternHistoryTable.scala 76:31]
    REG_45 <= io_windex == 3'h5; // @[PatternHistoryTable.scala 74:31]
    REG_46 <= io_waddr; // @[PatternHistoryTable.scala 75:31]
    REG_47 <= io_waddr; // @[PatternHistoryTable.scala 76:31]
    REG_48 <= io_windex == 3'h6; // @[PatternHistoryTable.scala 74:31]
    REG_49 <= io_waddr; // @[PatternHistoryTable.scala 75:31]
    REG_50 <= io_waddr; // @[PatternHistoryTable.scala 76:31]
    REG_51 <= io_windex == 3'h7; // @[PatternHistoryTable.scala 74:31]
    REG_52 <= io_waddr; // @[PatternHistoryTable.scala 75:31]
    REG_53 <= io_waddr; // @[PatternHistoryTable.scala 76:31]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_1_0[initvar] = _RAND_0[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_1_1[initvar] = _RAND_7[0:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_1_2[initvar] = _RAND_14[0:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_1_3[initvar] = _RAND_21[0:0];
  _RAND_28 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_1_4[initvar] = _RAND_28[0:0];
  _RAND_35 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_1_5[initvar] = _RAND_35[0:0];
  _RAND_42 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_1_6[initvar] = _RAND_42[0:0];
  _RAND_49 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_1_7[initvar] = _RAND_49[0:0];
  _RAND_56 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_0_0[initvar] = _RAND_56[0:0];
  _RAND_59 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_0_1[initvar] = _RAND_59[0:0];
  _RAND_62 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_0_2[initvar] = _RAND_62[0:0];
  _RAND_65 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_0_3[initvar] = _RAND_65[0:0];
  _RAND_68 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_0_4[initvar] = _RAND_68[0:0];
  _RAND_71 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_0_5[initvar] = _RAND_71[0:0];
  _RAND_74 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_0_6[initvar] = _RAND_74[0:0];
  _RAND_77 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    pht_0_7[initvar] = _RAND_77[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
//   pht_1_0_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  pht_1_0_MPORT_addr_pipe_0 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
//   pht_1_0_MPORT_8_en_pipe_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pht_1_0_MPORT_8_addr_pipe_0 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
//   pht_1_0_MPORT_16_en_pipe_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pht_1_0_MPORT_16_addr_pipe_0 = _RAND_6[5:0];
  _RAND_8 = {1{`RANDOM}};
//   pht_1_1_MPORT_1_en_pipe_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  pht_1_1_MPORT_1_addr_pipe_0 = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
//   pht_1_1_MPORT_9_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  pht_1_1_MPORT_9_addr_pipe_0 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
//   pht_1_1_MPORT_18_en_pipe_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  pht_1_1_MPORT_18_addr_pipe_0 = _RAND_13[5:0];
  _RAND_15 = {1{`RANDOM}};
//   pht_1_2_MPORT_2_en_pipe_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  pht_1_2_MPORT_2_addr_pipe_0 = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
//   pht_1_2_MPORT_10_en_pipe_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  pht_1_2_MPORT_10_addr_pipe_0 = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
//   pht_1_2_MPORT_20_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  pht_1_2_MPORT_20_addr_pipe_0 = _RAND_20[5:0];
  _RAND_22 = {1{`RANDOM}};
//   pht_1_3_MPORT_3_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  pht_1_3_MPORT_3_addr_pipe_0 = _RAND_23[5:0];
  _RAND_24 = {1{`RANDOM}};
//   pht_1_3_MPORT_11_en_pipe_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  pht_1_3_MPORT_11_addr_pipe_0 = _RAND_25[5:0];
  _RAND_26 = {1{`RANDOM}};
//   pht_1_3_MPORT_22_en_pipe_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  pht_1_3_MPORT_22_addr_pipe_0 = _RAND_27[5:0];
  _RAND_29 = {1{`RANDOM}};
//   pht_1_4_MPORT_4_en_pipe_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  pht_1_4_MPORT_4_addr_pipe_0 = _RAND_30[5:0];
  _RAND_31 = {1{`RANDOM}};
//   pht_1_4_MPORT_12_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  pht_1_4_MPORT_12_addr_pipe_0 = _RAND_32[5:0];
  _RAND_33 = {1{`RANDOM}};
//   pht_1_4_MPORT_24_en_pipe_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  pht_1_4_MPORT_24_addr_pipe_0 = _RAND_34[5:0];
  _RAND_36 = {1{`RANDOM}};
//   pht_1_5_MPORT_5_en_pipe_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  pht_1_5_MPORT_5_addr_pipe_0 = _RAND_37[5:0];
  _RAND_38 = {1{`RANDOM}};
//   pht_1_5_MPORT_13_en_pipe_0 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  pht_1_5_MPORT_13_addr_pipe_0 = _RAND_39[5:0];
  _RAND_40 = {1{`RANDOM}};
//   pht_1_5_MPORT_26_en_pipe_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  pht_1_5_MPORT_26_addr_pipe_0 = _RAND_41[5:0];
  _RAND_43 = {1{`RANDOM}};
//   pht_1_6_MPORT_6_en_pipe_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  pht_1_6_MPORT_6_addr_pipe_0 = _RAND_44[5:0];
  _RAND_45 = {1{`RANDOM}};
//   pht_1_6_MPORT_14_en_pipe_0 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  pht_1_6_MPORT_14_addr_pipe_0 = _RAND_46[5:0];
  _RAND_47 = {1{`RANDOM}};
//   pht_1_6_MPORT_28_en_pipe_0 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  pht_1_6_MPORT_28_addr_pipe_0 = _RAND_48[5:0];
  _RAND_50 = {1{`RANDOM}};
//   pht_1_7_MPORT_7_en_pipe_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  pht_1_7_MPORT_7_addr_pipe_0 = _RAND_51[5:0];
  _RAND_52 = {1{`RANDOM}};
//   pht_1_7_MPORT_15_en_pipe_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  pht_1_7_MPORT_15_addr_pipe_0 = _RAND_53[5:0];
  _RAND_54 = {1{`RANDOM}};
//   pht_1_7_MPORT_30_en_pipe_0 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  pht_1_7_MPORT_30_addr_pipe_0 = _RAND_55[5:0];
  _RAND_57 = {1{`RANDOM}};
//   pht_0_0_MPORT_17_en_pipe_0 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  pht_0_0_MPORT_17_addr_pipe_0 = _RAND_58[5:0];
  _RAND_60 = {1{`RANDOM}};
//   pht_0_1_MPORT_19_en_pipe_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  pht_0_1_MPORT_19_addr_pipe_0 = _RAND_61[5:0];
  _RAND_63 = {1{`RANDOM}};
//   pht_0_2_MPORT_21_en_pipe_0 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  pht_0_2_MPORT_21_addr_pipe_0 = _RAND_64[5:0];
  _RAND_66 = {1{`RANDOM}};
//   pht_0_3_MPORT_23_en_pipe_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  pht_0_3_MPORT_23_addr_pipe_0 = _RAND_67[5:0];
  _RAND_69 = {1{`RANDOM}};
//   pht_0_4_MPORT_25_en_pipe_0 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  pht_0_4_MPORT_25_addr_pipe_0 = _RAND_70[5:0];
  _RAND_72 = {1{`RANDOM}};
//   pht_0_5_MPORT_27_en_pipe_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  pht_0_5_MPORT_27_addr_pipe_0 = _RAND_73[5:0];
  _RAND_75 = {1{`RANDOM}};
//   pht_0_6_MPORT_29_en_pipe_0 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  pht_0_6_MPORT_29_addr_pipe_0 = _RAND_76[5:0];
  _RAND_78 = {1{`RANDOM}};
//   pht_0_7_MPORT_31_en_pipe_0 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  pht_0_7_MPORT_31_addr_pipe_0 = _RAND_79[5:0];
  _RAND_80 = {1{`RANDOM}};
  REG = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  REG_1 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  REG_2 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  REG_3 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  REG_4 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  REG_5 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  REG_6 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  REG_7 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  REG_8 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  REG_9 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  REG_10 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  REG_11 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  REG_12 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  REG_13 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  REG_14 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  REG_15 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  REG_16 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  REG_17 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  REG_18 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  REG_19 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  REG_20 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  REG_21 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  REG_22 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  REG_23 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  REG_24 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  REG_25 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  REG_26 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  REG_27 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  REG_28 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  REG_29 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  REG_30 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  REG_31 = _RAND_111[5:0];
  _RAND_112 = {1{`RANDOM}};
  REG_32 = _RAND_112[5:0];
  _RAND_113 = {1{`RANDOM}};
  REG_33 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  REG_34 = _RAND_114[5:0];
  _RAND_115 = {1{`RANDOM}};
  REG_35 = _RAND_115[5:0];
  _RAND_116 = {1{`RANDOM}};
  REG_36 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  REG_37 = _RAND_117[5:0];
  _RAND_118 = {1{`RANDOM}};
  REG_38 = _RAND_118[5:0];
  _RAND_119 = {1{`RANDOM}};
  REG_39 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  REG_40 = _RAND_120[5:0];
  _RAND_121 = {1{`RANDOM}};
  REG_41 = _RAND_121[5:0];
  _RAND_122 = {1{`RANDOM}};
  REG_42 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  REG_43 = _RAND_123[5:0];
  _RAND_124 = {1{`RANDOM}};
  REG_44 = _RAND_124[5:0];
  _RAND_125 = {1{`RANDOM}};
  REG_45 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  REG_46 = _RAND_126[5:0];
  _RAND_127 = {1{`RANDOM}};
  REG_47 = _RAND_127[5:0];
  _RAND_128 = {1{`RANDOM}};
  REG_48 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  REG_49 = _RAND_129[5:0];
  _RAND_130 = {1{`RANDOM}};
  REG_50 = _RAND_130[5:0];
  _RAND_131 = {1{`RANDOM}};
  REG_51 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  REG_52 = _RAND_132[5:0];
  _RAND_133 = {1{`RANDOM}};
  REG_53 = _RAND_133[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_BranchTargetBuffer4WayAssociative(
  input         clock,
  input         reset,
  input  [3:0]  io_raddr_0,
  input  [3:0]  io_raddr_1,
  input         io_ren_0,
  input         io_ren_1,
  input  [25:0] io_rtag_0,
  input  [25:0] io_rtag_1,
  output        io_rhit_0,
  output        io_rhit_1,
  output [31:0] io_rtarget_0,
  output [31:0] io_rtarget_1,
  input  [3:0]  io_waddr,
  input         io_wen,
  input  [25:0] io_wtag,
  input  [31:0] io_wtarget
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
`endif // RANDOMIZE_REG_INIT
  reg [25:0] btb_tag_0 [0:15]; // @[BranchTargetBuffer.scala 90:30]
//   wire  btb_tag_0_MPORT_en; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_addr; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_data; // @[BranchTargetBuffer.scala 90:30]
//   wire  btb_tag_0_MPORT_16_en; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_16_addr; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_16_data; // @[BranchTargetBuffer.scala 90:30]
//   wire  btb_tag_0_MPORT_32_en; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_32_addr; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_32_data; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_44_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_44_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_44_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_44_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_56_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_56_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_56_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_56_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_72_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_72_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_72_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_72_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_76_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_76_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_76_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_76_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_80_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_80_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_80_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_80_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_84_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_84_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_84_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_84_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_88_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_88_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_88_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_88_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_92_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_92_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_92_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_92_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_96_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_96_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_96_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_96_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_100_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_100_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_100_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_100_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_104_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_104_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_104_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_104_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_108_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_108_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_108_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_108_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_112_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_112_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_112_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_112_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_116_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_116_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_116_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_116_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_120_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_120_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_120_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_120_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_124_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_124_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_124_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_124_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_128_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_128_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_128_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_128_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_0_MPORT_132_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_0_MPORT_132_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_132_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_0_MPORT_132_en; // @[BranchTargetBuffer.scala 90:30]
//   reg  btb_tag_0_MPORT_en_pipe_0;
  reg [3:0] btb_tag_0_MPORT_addr_pipe_0;
//   reg  btb_tag_0_MPORT_16_en_pipe_0;
  reg [3:0] btb_tag_0_MPORT_16_addr_pipe_0;
//   reg  btb_tag_0_MPORT_32_en_pipe_0;
  reg [3:0] btb_tag_0_MPORT_32_addr_pipe_0;
  reg [25:0] btb_tag_1 [0:15]; // @[BranchTargetBuffer.scala 90:30]
//   wire  btb_tag_1_MPORT_4_en; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_4_addr; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_4_data; // @[BranchTargetBuffer.scala 90:30]
//   wire  btb_tag_1_MPORT_20_en; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_20_addr; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_20_data; // @[BranchTargetBuffer.scala 90:30]
//   wire  btb_tag_1_MPORT_35_en; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_35_addr; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_35_data; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_47_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_47_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_47_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_47_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_60_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_60_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_60_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_60_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_136_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_136_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_136_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_136_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_140_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_140_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_140_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_140_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_144_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_144_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_144_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_144_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_148_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_148_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_148_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_148_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_152_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_152_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_152_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_152_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_156_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_156_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_156_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_156_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_160_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_160_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_160_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_160_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_164_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_164_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_164_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_164_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_168_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_168_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_168_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_168_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_172_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_172_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_172_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_172_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_176_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_176_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_176_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_176_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_180_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_180_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_180_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_180_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_184_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_184_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_184_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_184_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_188_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_188_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_188_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_188_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_192_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_192_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_192_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_192_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_1_MPORT_196_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_1_MPORT_196_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_196_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_1_MPORT_196_en; // @[BranchTargetBuffer.scala 90:30]
//   reg  btb_tag_1_MPORT_4_en_pipe_0;
  reg [3:0] btb_tag_1_MPORT_4_addr_pipe_0;
//   reg  btb_tag_1_MPORT_20_en_pipe_0;
  reg [3:0] btb_tag_1_MPORT_20_addr_pipe_0;
//   reg  btb_tag_1_MPORT_35_en_pipe_0;
  reg [3:0] btb_tag_1_MPORT_35_addr_pipe_0;
  reg [25:0] btb_tag_2 [0:15]; // @[BranchTargetBuffer.scala 90:30]
//   wire  btb_tag_2_MPORT_8_en; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_8_addr; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_8_data; // @[BranchTargetBuffer.scala 90:30]
//   wire  btb_tag_2_MPORT_24_en; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_24_addr; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_24_data; // @[BranchTargetBuffer.scala 90:30]
//   wire  btb_tag_2_MPORT_38_en; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_38_addr; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_38_data; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_50_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_50_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_50_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_50_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_64_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_64_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_64_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_64_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_200_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_200_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_200_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_200_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_204_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_204_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_204_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_204_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_208_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_208_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_208_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_208_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_212_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_212_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_212_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_212_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_216_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_216_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_216_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_216_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_220_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_220_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_220_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_220_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_224_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_224_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_224_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_224_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_228_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_228_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_228_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_228_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_232_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_232_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_232_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_232_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_236_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_236_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_236_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_236_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_240_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_240_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_240_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_240_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_244_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_244_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_244_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_244_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_248_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_248_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_248_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_248_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_252_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_252_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_252_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_252_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_256_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_256_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_256_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_256_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_2_MPORT_260_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_2_MPORT_260_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_260_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_2_MPORT_260_en; // @[BranchTargetBuffer.scala 90:30]
//   reg  btb_tag_2_MPORT_8_en_pipe_0;
  reg [3:0] btb_tag_2_MPORT_8_addr_pipe_0;
//   reg  btb_tag_2_MPORT_24_en_pipe_0;
  reg [3:0] btb_tag_2_MPORT_24_addr_pipe_0;
//   reg  btb_tag_2_MPORT_38_en_pipe_0;
  reg [3:0] btb_tag_2_MPORT_38_addr_pipe_0;
  reg [25:0] btb_tag_3 [0:15]; // @[BranchTargetBuffer.scala 90:30]
//   wire  btb_tag_3_MPORT_12_en; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_12_addr; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_12_data; // @[BranchTargetBuffer.scala 90:30]
//   wire  btb_tag_3_MPORT_28_en; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_28_addr; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_28_data; // @[BranchTargetBuffer.scala 90:30]
//   wire  btb_tag_3_MPORT_41_en; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_41_addr; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_41_data; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_53_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_53_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_53_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_53_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_68_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_68_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_68_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_68_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_264_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_264_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_264_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_264_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_268_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_268_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_268_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_268_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_272_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_272_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_272_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_272_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_276_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_276_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_276_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_276_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_280_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_280_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_280_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_280_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_284_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_284_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_284_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_284_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_288_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_288_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_288_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_288_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_292_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_292_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_292_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_292_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_296_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_296_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_296_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_296_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_300_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_300_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_300_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_300_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_304_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_304_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_304_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_304_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_308_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_308_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_308_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_308_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_312_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_312_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_312_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_312_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_316_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_316_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_316_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_316_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_320_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_320_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_320_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_320_en; // @[BranchTargetBuffer.scala 90:30]
  wire [25:0] btb_tag_3_MPORT_324_data; // @[BranchTargetBuffer.scala 90:30]
  wire [3:0] btb_tag_3_MPORT_324_addr; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_324_mask; // @[BranchTargetBuffer.scala 90:30]
  wire  btb_tag_3_MPORT_324_en; // @[BranchTargetBuffer.scala 90:30]
//   reg  btb_tag_3_MPORT_12_en_pipe_0;
  reg [3:0] btb_tag_3_MPORT_12_addr_pipe_0;
//   reg  btb_tag_3_MPORT_28_en_pipe_0;
  reg [3:0] btb_tag_3_MPORT_28_addr_pipe_0;
//   reg  btb_tag_3_MPORT_41_en_pipe_0;
  reg [3:0] btb_tag_3_MPORT_41_addr_pipe_0;
  reg [31:0] btb_target_0 [0:15]; // @[BranchTargetBuffer.scala 94:33]
//   wire  btb_target_0_MPORT_1_en; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_1_addr; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_1_data; // @[BranchTargetBuffer.scala 94:33]
//   wire  btb_target_0_MPORT_17_en; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_17_addr; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_17_data; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_45_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_45_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_45_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_45_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_57_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_57_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_57_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_57_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_73_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_73_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_73_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_73_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_77_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_77_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_77_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_77_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_81_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_81_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_81_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_81_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_85_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_85_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_85_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_85_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_89_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_89_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_89_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_89_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_93_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_93_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_93_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_93_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_97_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_97_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_97_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_97_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_101_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_101_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_101_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_101_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_105_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_105_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_105_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_105_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_109_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_109_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_109_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_109_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_113_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_113_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_113_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_113_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_117_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_117_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_117_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_117_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_121_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_121_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_121_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_121_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_125_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_125_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_125_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_125_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_129_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_129_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_129_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_129_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_0_MPORT_133_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_0_MPORT_133_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_133_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_0_MPORT_133_en; // @[BranchTargetBuffer.scala 94:33]
//   reg  btb_target_0_MPORT_1_en_pipe_0;
  reg [3:0] btb_target_0_MPORT_1_addr_pipe_0;
//   reg  btb_target_0_MPORT_17_en_pipe_0;
  reg [3:0] btb_target_0_MPORT_17_addr_pipe_0;
  reg [31:0] btb_target_1 [0:15]; // @[BranchTargetBuffer.scala 94:33]
//   wire  btb_target_1_MPORT_5_en; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_5_addr; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_5_data; // @[BranchTargetBuffer.scala 94:33]
//   wire  btb_target_1_MPORT_21_en; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_21_addr; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_21_data; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_48_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_48_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_48_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_48_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_61_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_61_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_61_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_61_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_137_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_137_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_137_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_137_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_141_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_141_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_141_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_141_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_145_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_145_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_145_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_145_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_149_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_149_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_149_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_149_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_153_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_153_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_153_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_153_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_157_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_157_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_157_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_157_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_161_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_161_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_161_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_161_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_165_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_165_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_165_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_165_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_169_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_169_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_169_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_169_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_173_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_173_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_173_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_173_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_177_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_177_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_177_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_177_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_181_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_181_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_181_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_181_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_185_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_185_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_185_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_185_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_189_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_189_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_189_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_189_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_193_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_193_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_193_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_193_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_1_MPORT_197_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_1_MPORT_197_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_197_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_1_MPORT_197_en; // @[BranchTargetBuffer.scala 94:33]
//   reg  btb_target_1_MPORT_5_en_pipe_0;
  reg [3:0] btb_target_1_MPORT_5_addr_pipe_0;
//   reg  btb_target_1_MPORT_21_en_pipe_0;
  reg [3:0] btb_target_1_MPORT_21_addr_pipe_0;
  reg [31:0] btb_target_2 [0:15]; // @[BranchTargetBuffer.scala 94:33]
//   wire  btb_target_2_MPORT_9_en; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_9_addr; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_9_data; // @[BranchTargetBuffer.scala 94:33]
//   wire  btb_target_2_MPORT_25_en; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_25_addr; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_25_data; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_51_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_51_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_51_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_51_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_65_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_65_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_65_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_65_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_201_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_201_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_201_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_201_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_205_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_205_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_205_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_205_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_209_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_209_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_209_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_209_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_213_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_213_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_213_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_213_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_217_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_217_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_217_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_217_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_221_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_221_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_221_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_221_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_225_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_225_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_225_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_225_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_229_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_229_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_229_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_229_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_233_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_233_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_233_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_233_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_237_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_237_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_237_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_237_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_241_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_241_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_241_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_241_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_245_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_245_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_245_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_245_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_249_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_249_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_249_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_249_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_253_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_253_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_253_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_253_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_257_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_257_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_257_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_257_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_2_MPORT_261_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_2_MPORT_261_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_261_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_2_MPORT_261_en; // @[BranchTargetBuffer.scala 94:33]
//   reg  btb_target_2_MPORT_9_en_pipe_0;
  reg [3:0] btb_target_2_MPORT_9_addr_pipe_0;
//   reg  btb_target_2_MPORT_25_en_pipe_0;
  reg [3:0] btb_target_2_MPORT_25_addr_pipe_0;
  reg [31:0] btb_target_3 [0:15]; // @[BranchTargetBuffer.scala 94:33]
//   wire  btb_target_3_MPORT_13_en; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_13_addr; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_13_data; // @[BranchTargetBuffer.scala 94:33]
//   wire  btb_target_3_MPORT_29_en; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_29_addr; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_29_data; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_54_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_54_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_54_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_54_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_69_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_69_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_69_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_69_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_265_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_265_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_265_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_265_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_269_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_269_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_269_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_269_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_273_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_273_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_273_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_273_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_277_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_277_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_277_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_277_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_281_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_281_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_281_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_281_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_285_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_285_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_285_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_285_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_289_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_289_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_289_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_289_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_293_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_293_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_293_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_293_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_297_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_297_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_297_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_297_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_301_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_301_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_301_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_301_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_305_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_305_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_305_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_305_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_309_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_309_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_309_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_309_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_313_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_313_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_313_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_313_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_317_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_317_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_317_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_317_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_321_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_321_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_321_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_321_en; // @[BranchTargetBuffer.scala 94:33]
  wire [31:0] btb_target_3_MPORT_325_data; // @[BranchTargetBuffer.scala 94:33]
  wire [3:0] btb_target_3_MPORT_325_addr; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_325_mask; // @[BranchTargetBuffer.scala 94:33]
  wire  btb_target_3_MPORT_325_en; // @[BranchTargetBuffer.scala 94:33]
//   reg  btb_target_3_MPORT_13_en_pipe_0;
  reg [3:0] btb_target_3_MPORT_13_addr_pipe_0;
//   reg  btb_target_3_MPORT_29_en_pipe_0;
  reg [3:0] btb_target_3_MPORT_29_addr_pipe_0;
  reg  valid_0 [0:15]; // @[BranchTargetBuffer.scala 102:20]
//   wire  valid_0_MPORT_3_en; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_3_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_3_data; // @[BranchTargetBuffer.scala 102:20]
//   wire  valid_0_MPORT_19_en; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_19_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_19_data; // @[BranchTargetBuffer.scala 102:20]
//   wire  valid_0_MPORT_34_en; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_34_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_34_data; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_59_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_59_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_59_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_59_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_75_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_75_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_75_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_75_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_79_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_79_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_79_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_79_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_83_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_83_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_83_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_83_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_87_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_87_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_87_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_87_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_91_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_91_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_91_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_91_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_95_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_95_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_95_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_95_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_99_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_99_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_99_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_99_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_103_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_103_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_103_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_103_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_107_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_107_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_107_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_107_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_111_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_111_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_111_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_111_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_115_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_115_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_115_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_115_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_119_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_119_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_119_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_119_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_123_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_123_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_123_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_123_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_127_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_127_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_127_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_127_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_131_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_131_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_131_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_131_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_135_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_0_MPORT_135_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_135_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_0_MPORT_135_en; // @[BranchTargetBuffer.scala 102:20]
  reg  valid_1 [0:15]; // @[BranchTargetBuffer.scala 102:20]
//   wire  valid_1_MPORT_7_en; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_7_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_7_data; // @[BranchTargetBuffer.scala 102:20]
//   wire  valid_1_MPORT_23_en; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_23_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_23_data; // @[BranchTargetBuffer.scala 102:20]
//   wire  valid_1_MPORT_37_en; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_37_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_37_data; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_63_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_63_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_63_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_63_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_139_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_139_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_139_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_139_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_143_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_143_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_143_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_143_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_147_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_147_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_147_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_147_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_151_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_151_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_151_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_151_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_155_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_155_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_155_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_155_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_159_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_159_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_159_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_159_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_163_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_163_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_163_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_163_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_167_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_167_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_167_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_167_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_171_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_171_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_171_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_171_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_175_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_175_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_175_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_175_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_179_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_179_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_179_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_179_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_183_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_183_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_183_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_183_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_187_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_187_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_187_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_187_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_191_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_191_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_191_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_191_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_195_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_195_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_195_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_195_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_199_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_1_MPORT_199_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_199_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_1_MPORT_199_en; // @[BranchTargetBuffer.scala 102:20]
  reg  valid_2 [0:15]; // @[BranchTargetBuffer.scala 102:20]
//   wire  valid_2_MPORT_11_en; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_11_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_11_data; // @[BranchTargetBuffer.scala 102:20]
//   wire  valid_2_MPORT_27_en; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_27_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_27_data; // @[BranchTargetBuffer.scala 102:20]
//   wire  valid_2_MPORT_40_en; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_40_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_40_data; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_67_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_67_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_67_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_67_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_203_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_203_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_203_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_203_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_207_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_207_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_207_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_207_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_211_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_211_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_211_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_211_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_215_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_215_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_215_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_215_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_219_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_219_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_219_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_219_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_223_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_223_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_223_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_223_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_227_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_227_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_227_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_227_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_231_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_231_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_231_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_231_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_235_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_235_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_235_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_235_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_239_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_239_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_239_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_239_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_243_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_243_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_243_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_243_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_247_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_247_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_247_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_247_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_251_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_251_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_251_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_251_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_255_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_255_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_255_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_255_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_259_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_259_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_259_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_259_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_263_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_2_MPORT_263_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_263_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_2_MPORT_263_en; // @[BranchTargetBuffer.scala 102:20]
  reg  valid_3 [0:15]; // @[BranchTargetBuffer.scala 102:20]
//   wire  valid_3_MPORT_15_en; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_15_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_15_data; // @[BranchTargetBuffer.scala 102:20]
//   wire  valid_3_MPORT_31_en; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_31_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_31_data; // @[BranchTargetBuffer.scala 102:20]
//   wire  valid_3_MPORT_43_en; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_43_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_43_data; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_71_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_71_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_71_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_71_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_267_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_267_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_267_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_267_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_271_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_271_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_271_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_271_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_275_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_275_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_275_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_275_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_279_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_279_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_279_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_279_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_283_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_283_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_283_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_283_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_287_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_287_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_287_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_287_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_291_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_291_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_291_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_291_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_295_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_295_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_295_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_295_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_299_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_299_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_299_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_299_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_303_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_303_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_303_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_303_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_307_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_307_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_307_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_307_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_311_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_311_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_311_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_311_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_315_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_315_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_315_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_315_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_319_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_319_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_319_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_319_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_323_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_323_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_323_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_323_en; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_327_data; // @[BranchTargetBuffer.scala 102:20]
  wire [3:0] valid_3_MPORT_327_addr; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_327_mask; // @[BranchTargetBuffer.scala 102:20]
  wire  valid_3_MPORT_327_en; // @[BranchTargetBuffer.scala 102:20]
  reg  plru0_0; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_1; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_2; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_3; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_4; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_5; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_6; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_7; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_8; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_9; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_10; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_11; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_12; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_13; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_14; // @[BranchTargetBuffer.scala 107:22]
  reg  plru0_15; // @[BranchTargetBuffer.scala 107:22]
  reg  plru1_0; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_1; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_2; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_3; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_4; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_5; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_6; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_7; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_8; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_9; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_10; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_11; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_12; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_13; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_14; // @[BranchTargetBuffer.scala 109:22]
  reg  plru1_15; // @[BranchTargetBuffer.scala 109:22]
  reg  plru2_0; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_1; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_2; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_3; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_4; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_5; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_6; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_7; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_8; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_9; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_10; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_11; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_12; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_13; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_14; // @[BranchTargetBuffer.scala 111:22]
  reg  plru2_15; // @[BranchTargetBuffer.scala 111:22]
  reg  REG__0; // @[BranchTargetBuffer.scala 124:25]
  reg  REG__1; // @[BranchTargetBuffer.scala 124:25]
  reg  REG__2; // @[BranchTargetBuffer.scala 124:25]
  reg  REG__3; // @[BranchTargetBuffer.scala 124:25]
  reg [25:0] REG_1; // @[BranchTargetBuffer.scala 133:51]
  wire [25:0] _WIRE_8_0_tag = btb_tag_0_MPORT_data;
  reg  REG_2; // @[BranchTargetBuffer.scala 137:22]
  reg [3:0] REG_3; // @[BranchTargetBuffer.scala 138:33]
  wire  _GEN_2891 = 4'h0 == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_6 = 4'h0 == REG_3 | plru0_0; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2892 = 4'h1 == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_7 = 4'h1 == REG_3 | plru0_1; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2893 = 4'h2 == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_8 = 4'h2 == REG_3 | plru0_2; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2894 = 4'h3 == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_9 = 4'h3 == REG_3 | plru0_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2895 = 4'h4 == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_10 = 4'h4 == REG_3 | plru0_4; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2896 = 4'h5 == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_11 = 4'h5 == REG_3 | plru0_5; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2897 = 4'h6 == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_12 = 4'h6 == REG_3 | plru0_6; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2898 = 4'h7 == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_13 = 4'h7 == REG_3 | plru0_7; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2899 = 4'h8 == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_14 = 4'h8 == REG_3 | plru0_8; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2900 = 4'h9 == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_15 = 4'h9 == REG_3 | plru0_9; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2901 = 4'ha == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_16 = 4'ha == REG_3 | plru0_10; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2902 = 4'hb == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_17 = 4'hb == REG_3 | plru0_11; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2903 = 4'hc == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_18 = 4'hc == REG_3 | plru0_12; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2904 = 4'hd == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_19 = 4'hd == REG_3 | plru0_13; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2905 = 4'he == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_20 = 4'he == REG_3 | plru0_14; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_2906 = 4'hf == REG_3; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_21 = 4'hf == REG_3 | plru0_15; // @[BranchTargetBuffer.scala 114:{16,16} 107:22]
  wire  _GEN_22 = _GEN_2891 | plru1_0; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_23 = _GEN_2892 | plru1_1; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_24 = _GEN_2893 | plru1_2; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_25 = _GEN_2894 | plru1_3; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_26 = _GEN_2895 | plru1_4; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_27 = _GEN_2896 | plru1_5; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_28 = _GEN_2897 | plru1_6; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_29 = _GEN_2898 | plru1_7; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_30 = _GEN_2899 | plru1_8; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_31 = _GEN_2900 | plru1_9; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_32 = _GEN_2901 | plru1_10; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_33 = _GEN_2902 | plru1_11; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_34 = _GEN_2903 | plru1_12; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_35 = _GEN_2904 | plru1_13; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_36 = _GEN_2905 | plru1_14; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_37 = _GEN_2906 | plru1_15; // @[BranchTargetBuffer.scala 116:{18,18} 109:22]
  wire  _GEN_86 = REG_2 ? _GEN_6 : plru0_0; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_87 = REG_2 ? _GEN_7 : plru0_1; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_88 = REG_2 ? _GEN_8 : plru0_2; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_89 = REG_2 ? _GEN_9 : plru0_3; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_90 = REG_2 ? _GEN_10 : plru0_4; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_91 = REG_2 ? _GEN_11 : plru0_5; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_92 = REG_2 ? _GEN_12 : plru0_6; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_93 = REG_2 ? _GEN_13 : plru0_7; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_94 = REG_2 ? _GEN_14 : plru0_8; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_95 = REG_2 ? _GEN_15 : plru0_9; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_96 = REG_2 ? _GEN_16 : plru0_10; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_97 = REG_2 ? _GEN_17 : plru0_11; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_98 = REG_2 ? _GEN_18 : plru0_12; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_99 = REG_2 ? _GEN_19 : plru0_13; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_100 = REG_2 ? _GEN_20 : plru0_14; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_101 = REG_2 ? _GEN_21 : plru0_15; // @[BranchTargetBuffer.scala 107:22 137:35]
  wire  _GEN_102 = REG_2 ? _GEN_22 : plru1_0; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_103 = REG_2 ? _GEN_23 : plru1_1; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_104 = REG_2 ? _GEN_24 : plru1_2; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_105 = REG_2 ? _GEN_25 : plru1_3; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_106 = REG_2 ? _GEN_26 : plru1_4; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_107 = REG_2 ? _GEN_27 : plru1_5; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_108 = REG_2 ? _GEN_28 : plru1_6; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_109 = REG_2 ? _GEN_29 : plru1_7; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_110 = REG_2 ? _GEN_30 : plru1_8; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_111 = REG_2 ? _GEN_31 : plru1_9; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_112 = REG_2 ? _GEN_32 : plru1_10; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_113 = REG_2 ? _GEN_33 : plru1_11; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_114 = REG_2 ? _GEN_34 : plru1_12; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_115 = REG_2 ? _GEN_35 : plru1_13; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_116 = REG_2 ? _GEN_36 : plru1_14; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire  _GEN_117 = REG_2 ? _GEN_37 : plru1_15; // @[BranchTargetBuffer.scala 109:22 137:35]
  wire [31:0] _WIRE_8_0_target = btb_target_0_MPORT_1_data;
  wire [31:0] _GEN_135 = REG__0 & _WIRE_8_0_tag == REG_1 ? _WIRE_8_0_target : 32'h0; // @[BranchTargetBuffer.scala 126:19 133:66 135:23]
  wire  _GEN_137 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_86 : plru0_0; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_138 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_87 : plru0_1; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_139 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_88 : plru0_2; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_140 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_89 : plru0_3; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_141 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_90 : plru0_4; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_142 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_91 : plru0_5; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_143 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_92 : plru0_6; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_144 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_93 : plru0_7; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_145 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_94 : plru0_8; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_146 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_95 : plru0_9; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_147 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_96 : plru0_10; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_148 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_97 : plru0_11; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_149 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_98 : plru0_12; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_150 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_99 : plru0_13; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_151 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_100 : plru0_14; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_152 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_101 : plru0_15; // @[BranchTargetBuffer.scala 107:22 133:66]
  wire  _GEN_153 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_102 : plru1_0; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_154 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_103 : plru1_1; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_155 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_104 : plru1_2; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_156 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_105 : plru1_3; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_157 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_106 : plru1_4; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_158 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_107 : plru1_5; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_159 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_108 : plru1_6; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_160 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_109 : plru1_7; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_161 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_110 : plru1_8; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_162 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_111 : plru1_9; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_163 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_112 : plru1_10; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_164 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_113 : plru1_11; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_165 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_114 : plru1_12; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_166 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_115 : plru1_13; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_167 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_116 : plru1_14; // @[BranchTargetBuffer.scala 109:22 133:66]
  wire  _GEN_168 = REG__0 & _WIRE_8_0_tag == REG_1 ? _GEN_117 : plru1_15; // @[BranchTargetBuffer.scala 109:22 133:66]
  reg [25:0] REG_4; // @[BranchTargetBuffer.scala 133:51]
  wire [25:0] _WIRE_8_1_tag = btb_tag_1_MPORT_4_data;
  reg  REG_5; // @[BranchTargetBuffer.scala 137:22]
  reg [3:0] REG_6; // @[BranchTargetBuffer.scala 138:33]
  wire  _GEN_188 = 4'h0 == REG_6 | _GEN_137; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_189 = 4'h1 == REG_6 | _GEN_138; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_190 = 4'h2 == REG_6 | _GEN_139; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_191 = 4'h3 == REG_6 | _GEN_140; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_192 = 4'h4 == REG_6 | _GEN_141; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_193 = 4'h5 == REG_6 | _GEN_142; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_194 = 4'h6 == REG_6 | _GEN_143; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_195 = 4'h7 == REG_6 | _GEN_144; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_196 = 4'h8 == REG_6 | _GEN_145; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_197 = 4'h9 == REG_6 | _GEN_146; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_198 = 4'ha == REG_6 | _GEN_147; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_199 = 4'hb == REG_6 | _GEN_148; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_200 = 4'hc == REG_6 | _GEN_149; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_201 = 4'hd == REG_6 | _GEN_150; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_202 = 4'he == REG_6 | _GEN_151; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_203 = 4'hf == REG_6 | _GEN_152; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_204 = 4'h0 == REG_6 ? 1'h0 : _GEN_153; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_205 = 4'h1 == REG_6 ? 1'h0 : _GEN_154; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_206 = 4'h2 == REG_6 ? 1'h0 : _GEN_155; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_207 = 4'h3 == REG_6 ? 1'h0 : _GEN_156; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_208 = 4'h4 == REG_6 ? 1'h0 : _GEN_157; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_209 = 4'h5 == REG_6 ? 1'h0 : _GEN_158; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_210 = 4'h6 == REG_6 ? 1'h0 : _GEN_159; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_211 = 4'h7 == REG_6 ? 1'h0 : _GEN_160; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_212 = 4'h8 == REG_6 ? 1'h0 : _GEN_161; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_213 = 4'h9 == REG_6 ? 1'h0 : _GEN_162; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_214 = 4'ha == REG_6 ? 1'h0 : _GEN_163; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_215 = 4'hb == REG_6 ? 1'h0 : _GEN_164; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_216 = 4'hc == REG_6 ? 1'h0 : _GEN_165; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_217 = 4'hd == REG_6 ? 1'h0 : _GEN_166; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_218 = 4'he == REG_6 ? 1'h0 : _GEN_167; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_219 = 4'hf == REG_6 ? 1'h0 : _GEN_168; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_268 = REG_5 ? _GEN_188 : _GEN_137; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_269 = REG_5 ? _GEN_189 : _GEN_138; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_270 = REG_5 ? _GEN_190 : _GEN_139; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_271 = REG_5 ? _GEN_191 : _GEN_140; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_272 = REG_5 ? _GEN_192 : _GEN_141; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_273 = REG_5 ? _GEN_193 : _GEN_142; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_274 = REG_5 ? _GEN_194 : _GEN_143; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_275 = REG_5 ? _GEN_195 : _GEN_144; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_276 = REG_5 ? _GEN_196 : _GEN_145; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_277 = REG_5 ? _GEN_197 : _GEN_146; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_278 = REG_5 ? _GEN_198 : _GEN_147; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_279 = REG_5 ? _GEN_199 : _GEN_148; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_280 = REG_5 ? _GEN_200 : _GEN_149; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_281 = REG_5 ? _GEN_201 : _GEN_150; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_282 = REG_5 ? _GEN_202 : _GEN_151; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_283 = REG_5 ? _GEN_203 : _GEN_152; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_284 = REG_5 ? _GEN_204 : _GEN_153; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_285 = REG_5 ? _GEN_205 : _GEN_154; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_286 = REG_5 ? _GEN_206 : _GEN_155; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_287 = REG_5 ? _GEN_207 : _GEN_156; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_288 = REG_5 ? _GEN_208 : _GEN_157; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_289 = REG_5 ? _GEN_209 : _GEN_158; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_290 = REG_5 ? _GEN_210 : _GEN_159; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_291 = REG_5 ? _GEN_211 : _GEN_160; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_292 = REG_5 ? _GEN_212 : _GEN_161; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_293 = REG_5 ? _GEN_213 : _GEN_162; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_294 = REG_5 ? _GEN_214 : _GEN_163; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_295 = REG_5 ? _GEN_215 : _GEN_164; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_296 = REG_5 ? _GEN_216 : _GEN_165; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_297 = REG_5 ? _GEN_217 : _GEN_166; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_298 = REG_5 ? _GEN_218 : _GEN_167; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_299 = REG_5 ? _GEN_219 : _GEN_168; // @[BranchTargetBuffer.scala 137:35]
  wire [31:0] _WIRE_8_1_target = btb_target_1_MPORT_5_data;
  wire [31:0] _GEN_317 = REG__1 & _WIRE_8_1_tag == REG_4 ? _WIRE_8_1_target : _GEN_135; // @[BranchTargetBuffer.scala 133:66 135:23]
  wire  _GEN_319 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_268 : _GEN_137; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_320 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_269 : _GEN_138; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_321 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_270 : _GEN_139; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_322 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_271 : _GEN_140; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_323 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_272 : _GEN_141; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_324 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_273 : _GEN_142; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_325 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_274 : _GEN_143; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_326 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_275 : _GEN_144; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_327 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_276 : _GEN_145; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_328 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_277 : _GEN_146; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_329 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_278 : _GEN_147; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_330 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_279 : _GEN_148; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_331 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_280 : _GEN_149; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_332 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_281 : _GEN_150; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_333 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_282 : _GEN_151; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_334 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_283 : _GEN_152; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_335 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_284 : _GEN_153; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_336 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_285 : _GEN_154; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_337 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_286 : _GEN_155; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_338 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_287 : _GEN_156; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_339 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_288 : _GEN_157; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_340 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_289 : _GEN_158; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_341 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_290 : _GEN_159; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_342 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_291 : _GEN_160; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_343 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_292 : _GEN_161; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_344 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_293 : _GEN_162; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_345 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_294 : _GEN_163; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_346 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_295 : _GEN_164; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_347 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_296 : _GEN_165; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_348 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_297 : _GEN_166; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_349 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_298 : _GEN_167; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_350 = REG__1 & _WIRE_8_1_tag == REG_4 ? _GEN_299 : _GEN_168; // @[BranchTargetBuffer.scala 133:66]
  reg [25:0] REG_7; // @[BranchTargetBuffer.scala 133:51]
  wire [25:0] _WIRE_8_2_tag = btb_tag_2_MPORT_8_data;
  reg  REG_8; // @[BranchTargetBuffer.scala 137:22]
  reg [3:0] REG_9; // @[BranchTargetBuffer.scala 138:33]
  wire  _GEN_370 = 4'h0 == REG_9 ? 1'h0 : _GEN_319; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_371 = 4'h1 == REG_9 ? 1'h0 : _GEN_320; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_372 = 4'h2 == REG_9 ? 1'h0 : _GEN_321; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_373 = 4'h3 == REG_9 ? 1'h0 : _GEN_322; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_374 = 4'h4 == REG_9 ? 1'h0 : _GEN_323; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_375 = 4'h5 == REG_9 ? 1'h0 : _GEN_324; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_376 = 4'h6 == REG_9 ? 1'h0 : _GEN_325; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_377 = 4'h7 == REG_9 ? 1'h0 : _GEN_326; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_378 = 4'h8 == REG_9 ? 1'h0 : _GEN_327; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_379 = 4'h9 == REG_9 ? 1'h0 : _GEN_328; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_380 = 4'ha == REG_9 ? 1'h0 : _GEN_329; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_381 = 4'hb == REG_9 ? 1'h0 : _GEN_330; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_382 = 4'hc == REG_9 ? 1'h0 : _GEN_331; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_383 = 4'hd == REG_9 ? 1'h0 : _GEN_332; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_384 = 4'he == REG_9 ? 1'h0 : _GEN_333; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_385 = 4'hf == REG_9 ? 1'h0 : _GEN_334; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2955 = 4'h0 == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2956 = 4'h1 == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2957 = 4'h2 == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2958 = 4'h3 == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2959 = 4'h4 == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2960 = 4'h5 == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2961 = 4'h6 == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2962 = 4'h7 == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2963 = 4'h8 == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2964 = 4'h9 == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2965 = 4'ha == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2966 = 4'hb == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2967 = 4'hc == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2968 = 4'hd == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2969 = 4'he == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2970 = 4'hf == REG_9; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_402 = _GEN_2955 | plru2_0; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_403 = _GEN_2956 | plru2_1; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_404 = _GEN_2957 | plru2_2; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_405 = _GEN_2958 | plru2_3; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_406 = _GEN_2959 | plru2_4; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_407 = _GEN_2960 | plru2_5; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_408 = _GEN_2961 | plru2_6; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_409 = _GEN_2962 | plru2_7; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_410 = _GEN_2963 | plru2_8; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_411 = _GEN_2964 | plru2_9; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_412 = _GEN_2965 | plru2_10; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_413 = _GEN_2966 | plru2_11; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_414 = _GEN_2967 | plru2_12; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_415 = _GEN_2968 | plru2_13; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_416 = _GEN_2969 | plru2_14; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_417 = _GEN_2970 | plru2_15; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_450 = REG_8 ? _GEN_370 : _GEN_319; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_451 = REG_8 ? _GEN_371 : _GEN_320; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_452 = REG_8 ? _GEN_372 : _GEN_321; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_453 = REG_8 ? _GEN_373 : _GEN_322; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_454 = REG_8 ? _GEN_374 : _GEN_323; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_455 = REG_8 ? _GEN_375 : _GEN_324; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_456 = REG_8 ? _GEN_376 : _GEN_325; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_457 = REG_8 ? _GEN_377 : _GEN_326; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_458 = REG_8 ? _GEN_378 : _GEN_327; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_459 = REG_8 ? _GEN_379 : _GEN_328; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_460 = REG_8 ? _GEN_380 : _GEN_329; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_461 = REG_8 ? _GEN_381 : _GEN_330; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_462 = REG_8 ? _GEN_382 : _GEN_331; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_463 = REG_8 ? _GEN_383 : _GEN_332; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_464 = REG_8 ? _GEN_384 : _GEN_333; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_465 = REG_8 ? _GEN_385 : _GEN_334; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_482 = REG_8 ? _GEN_402 : plru2_0; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_483 = REG_8 ? _GEN_403 : plru2_1; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_484 = REG_8 ? _GEN_404 : plru2_2; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_485 = REG_8 ? _GEN_405 : plru2_3; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_486 = REG_8 ? _GEN_406 : plru2_4; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_487 = REG_8 ? _GEN_407 : plru2_5; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_488 = REG_8 ? _GEN_408 : plru2_6; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_489 = REG_8 ? _GEN_409 : plru2_7; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_490 = REG_8 ? _GEN_410 : plru2_8; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_491 = REG_8 ? _GEN_411 : plru2_9; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_492 = REG_8 ? _GEN_412 : plru2_10; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_493 = REG_8 ? _GEN_413 : plru2_11; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_494 = REG_8 ? _GEN_414 : plru2_12; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_495 = REG_8 ? _GEN_415 : plru2_13; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_496 = REG_8 ? _GEN_416 : plru2_14; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_497 = REG_8 ? _GEN_417 : plru2_15; // @[BranchTargetBuffer.scala 137:35]
  wire [31:0] _WIRE_8_2_target = btb_target_2_MPORT_9_data;
  wire [31:0] _GEN_499 = REG__2 & _WIRE_8_2_tag == REG_7 ? _WIRE_8_2_target : _GEN_317; // @[BranchTargetBuffer.scala 133:66 135:23]
  wire  _GEN_501 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_450 : _GEN_319; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_502 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_451 : _GEN_320; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_503 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_452 : _GEN_321; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_504 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_453 : _GEN_322; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_505 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_454 : _GEN_323; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_506 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_455 : _GEN_324; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_507 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_456 : _GEN_325; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_508 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_457 : _GEN_326; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_509 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_458 : _GEN_327; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_510 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_459 : _GEN_328; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_511 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_460 : _GEN_329; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_512 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_461 : _GEN_330; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_513 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_462 : _GEN_331; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_514 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_463 : _GEN_332; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_515 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_464 : _GEN_333; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_516 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_465 : _GEN_334; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_533 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_482 : plru2_0; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_534 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_483 : plru2_1; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_535 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_484 : plru2_2; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_536 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_485 : plru2_3; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_537 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_486 : plru2_4; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_538 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_487 : plru2_5; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_539 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_488 : plru2_6; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_540 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_489 : plru2_7; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_541 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_490 : plru2_8; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_542 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_491 : plru2_9; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_543 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_492 : plru2_10; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_544 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_493 : plru2_11; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_545 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_494 : plru2_12; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_546 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_495 : plru2_13; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_547 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_496 : plru2_14; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_548 = REG__2 & _WIRE_8_2_tag == REG_7 ? _GEN_497 : plru2_15; // @[BranchTargetBuffer.scala 133:66]
  reg [25:0] REG_10; // @[BranchTargetBuffer.scala 133:51]
  wire [25:0] _WIRE_8_3_tag = btb_tag_3_MPORT_12_data;
  reg  REG_11; // @[BranchTargetBuffer.scala 137:22]
  reg [3:0] REG_12; // @[BranchTargetBuffer.scala 138:33]
  wire  _GEN_552 = 4'h0 == REG_12 ? 1'h0 : _GEN_501; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_553 = 4'h1 == REG_12 ? 1'h0 : _GEN_502; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_554 = 4'h2 == REG_12 ? 1'h0 : _GEN_503; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_555 = 4'h3 == REG_12 ? 1'h0 : _GEN_504; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_556 = 4'h4 == REG_12 ? 1'h0 : _GEN_505; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_557 = 4'h5 == REG_12 ? 1'h0 : _GEN_506; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_558 = 4'h6 == REG_12 ? 1'h0 : _GEN_507; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_559 = 4'h7 == REG_12 ? 1'h0 : _GEN_508; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_560 = 4'h8 == REG_12 ? 1'h0 : _GEN_509; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_561 = 4'h9 == REG_12 ? 1'h0 : _GEN_510; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_562 = 4'ha == REG_12 ? 1'h0 : _GEN_511; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_563 = 4'hb == REG_12 ? 1'h0 : _GEN_512; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_564 = 4'hc == REG_12 ? 1'h0 : _GEN_513; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_565 = 4'hd == REG_12 ? 1'h0 : _GEN_514; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_566 = 4'he == REG_12 ? 1'h0 : _GEN_515; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_567 = 4'hf == REG_12 ? 1'h0 : _GEN_516; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_584 = 4'h0 == REG_12 ? 1'h0 : _GEN_533; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_585 = 4'h1 == REG_12 ? 1'h0 : _GEN_534; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_586 = 4'h2 == REG_12 ? 1'h0 : _GEN_535; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_587 = 4'h3 == REG_12 ? 1'h0 : _GEN_536; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_588 = 4'h4 == REG_12 ? 1'h0 : _GEN_537; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_589 = 4'h5 == REG_12 ? 1'h0 : _GEN_538; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_590 = 4'h6 == REG_12 ? 1'h0 : _GEN_539; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_591 = 4'h7 == REG_12 ? 1'h0 : _GEN_540; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_592 = 4'h8 == REG_12 ? 1'h0 : _GEN_541; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_593 = 4'h9 == REG_12 ? 1'h0 : _GEN_542; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_594 = 4'ha == REG_12 ? 1'h0 : _GEN_543; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_595 = 4'hb == REG_12 ? 1'h0 : _GEN_544; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_596 = 4'hc == REG_12 ? 1'h0 : _GEN_545; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_597 = 4'hd == REG_12 ? 1'h0 : _GEN_546; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_598 = 4'he == REG_12 ? 1'h0 : _GEN_547; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_599 = 4'hf == REG_12 ? 1'h0 : _GEN_548; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_632 = REG_11 ? _GEN_552 : _GEN_501; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_633 = REG_11 ? _GEN_553 : _GEN_502; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_634 = REG_11 ? _GEN_554 : _GEN_503; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_635 = REG_11 ? _GEN_555 : _GEN_504; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_636 = REG_11 ? _GEN_556 : _GEN_505; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_637 = REG_11 ? _GEN_557 : _GEN_506; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_638 = REG_11 ? _GEN_558 : _GEN_507; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_639 = REG_11 ? _GEN_559 : _GEN_508; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_640 = REG_11 ? _GEN_560 : _GEN_509; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_641 = REG_11 ? _GEN_561 : _GEN_510; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_642 = REG_11 ? _GEN_562 : _GEN_511; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_643 = REG_11 ? _GEN_563 : _GEN_512; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_644 = REG_11 ? _GEN_564 : _GEN_513; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_645 = REG_11 ? _GEN_565 : _GEN_514; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_646 = REG_11 ? _GEN_566 : _GEN_515; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_647 = REG_11 ? _GEN_567 : _GEN_516; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_664 = REG_11 ? _GEN_584 : _GEN_533; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_665 = REG_11 ? _GEN_585 : _GEN_534; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_666 = REG_11 ? _GEN_586 : _GEN_535; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_667 = REG_11 ? _GEN_587 : _GEN_536; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_668 = REG_11 ? _GEN_588 : _GEN_537; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_669 = REG_11 ? _GEN_589 : _GEN_538; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_670 = REG_11 ? _GEN_590 : _GEN_539; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_671 = REG_11 ? _GEN_591 : _GEN_540; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_672 = REG_11 ? _GEN_592 : _GEN_541; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_673 = REG_11 ? _GEN_593 : _GEN_542; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_674 = REG_11 ? _GEN_594 : _GEN_543; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_675 = REG_11 ? _GEN_595 : _GEN_544; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_676 = REG_11 ? _GEN_596 : _GEN_545; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_677 = REG_11 ? _GEN_597 : _GEN_546; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_678 = REG_11 ? _GEN_598 : _GEN_547; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_679 = REG_11 ? _GEN_599 : _GEN_548; // @[BranchTargetBuffer.scala 137:35]
  wire [31:0] _WIRE_8_3_target = btb_target_3_MPORT_13_data;
  wire  _GEN_683 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_632 : _GEN_501; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_684 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_633 : _GEN_502; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_685 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_634 : _GEN_503; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_686 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_635 : _GEN_504; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_687 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_636 : _GEN_505; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_688 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_637 : _GEN_506; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_689 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_638 : _GEN_507; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_690 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_639 : _GEN_508; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_691 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_640 : _GEN_509; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_692 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_641 : _GEN_510; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_693 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_642 : _GEN_511; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_694 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_643 : _GEN_512; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_695 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_644 : _GEN_513; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_696 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_645 : _GEN_514; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_697 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_646 : _GEN_515; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_698 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_647 : _GEN_516; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_715 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_664 : _GEN_533; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_716 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_665 : _GEN_534; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_717 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_666 : _GEN_535; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_718 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_667 : _GEN_536; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_719 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_668 : _GEN_537; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_720 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_669 : _GEN_538; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_721 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_670 : _GEN_539; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_722 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_671 : _GEN_540; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_723 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_672 : _GEN_541; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_724 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_673 : _GEN_542; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_725 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_674 : _GEN_543; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_726 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_675 : _GEN_544; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_727 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_676 : _GEN_545; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_728 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_677 : _GEN_546; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_729 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_678 : _GEN_547; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_730 = REG__3 & _WIRE_8_3_tag == REG_10 ? _GEN_679 : _GEN_548; // @[BranchTargetBuffer.scala 133:66]
  reg  REG_13_0; // @[BranchTargetBuffer.scala 124:25]
  reg  REG_13_1; // @[BranchTargetBuffer.scala 124:25]
  reg  REG_13_2; // @[BranchTargetBuffer.scala 124:25]
  reg  REG_13_3; // @[BranchTargetBuffer.scala 124:25]
  reg [25:0] REG_14; // @[BranchTargetBuffer.scala 133:51]
  wire [25:0] _WIRE_27_0_tag = btb_tag_0_MPORT_16_data;
  reg  REG_15; // @[BranchTargetBuffer.scala 137:22]
  reg [3:0] REG_16; // @[BranchTargetBuffer.scala 138:33]
  wire  _GEN_2987 = 4'h0 == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_735 = 4'h0 == REG_16 | _GEN_683; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2988 = 4'h1 == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_736 = 4'h1 == REG_16 | _GEN_684; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2989 = 4'h2 == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_737 = 4'h2 == REG_16 | _GEN_685; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2990 = 4'h3 == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_738 = 4'h3 == REG_16 | _GEN_686; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2991 = 4'h4 == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_739 = 4'h4 == REG_16 | _GEN_687; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2992 = 4'h5 == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_740 = 4'h5 == REG_16 | _GEN_688; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2993 = 4'h6 == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_741 = 4'h6 == REG_16 | _GEN_689; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2994 = 4'h7 == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_742 = 4'h7 == REG_16 | _GEN_690; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2995 = 4'h8 == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_743 = 4'h8 == REG_16 | _GEN_691; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2996 = 4'h9 == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_744 = 4'h9 == REG_16 | _GEN_692; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2997 = 4'ha == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_745 = 4'ha == REG_16 | _GEN_693; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2998 = 4'hb == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_746 = 4'hb == REG_16 | _GEN_694; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2999 = 4'hc == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_747 = 4'hc == REG_16 | _GEN_695; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3000 = 4'hd == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_748 = 4'hd == REG_16 | _GEN_696; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3001 = 4'he == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_749 = 4'he == REG_16 | _GEN_697; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3002 = 4'hf == REG_16; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_750 = 4'hf == REG_16 | _GEN_698; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_751 = _GEN_2987 | _GEN_335; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_752 = _GEN_2988 | _GEN_336; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_753 = _GEN_2989 | _GEN_337; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_754 = _GEN_2990 | _GEN_338; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_755 = _GEN_2991 | _GEN_339; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_756 = _GEN_2992 | _GEN_340; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_757 = _GEN_2993 | _GEN_341; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_758 = _GEN_2994 | _GEN_342; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_759 = _GEN_2995 | _GEN_343; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_760 = _GEN_2996 | _GEN_344; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_761 = _GEN_2997 | _GEN_345; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_762 = _GEN_2998 | _GEN_346; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_763 = _GEN_2999 | _GEN_347; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_764 = _GEN_3000 | _GEN_348; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_765 = _GEN_3001 | _GEN_349; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_766 = _GEN_3002 | _GEN_350; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_815 = REG_15 ? _GEN_735 : _GEN_683; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_816 = REG_15 ? _GEN_736 : _GEN_684; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_817 = REG_15 ? _GEN_737 : _GEN_685; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_818 = REG_15 ? _GEN_738 : _GEN_686; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_819 = REG_15 ? _GEN_739 : _GEN_687; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_820 = REG_15 ? _GEN_740 : _GEN_688; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_821 = REG_15 ? _GEN_741 : _GEN_689; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_822 = REG_15 ? _GEN_742 : _GEN_690; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_823 = REG_15 ? _GEN_743 : _GEN_691; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_824 = REG_15 ? _GEN_744 : _GEN_692; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_825 = REG_15 ? _GEN_745 : _GEN_693; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_826 = REG_15 ? _GEN_746 : _GEN_694; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_827 = REG_15 ? _GEN_747 : _GEN_695; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_828 = REG_15 ? _GEN_748 : _GEN_696; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_829 = REG_15 ? _GEN_749 : _GEN_697; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_830 = REG_15 ? _GEN_750 : _GEN_698; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_831 = REG_15 ? _GEN_751 : _GEN_335; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_832 = REG_15 ? _GEN_752 : _GEN_336; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_833 = REG_15 ? _GEN_753 : _GEN_337; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_834 = REG_15 ? _GEN_754 : _GEN_338; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_835 = REG_15 ? _GEN_755 : _GEN_339; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_836 = REG_15 ? _GEN_756 : _GEN_340; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_837 = REG_15 ? _GEN_757 : _GEN_341; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_838 = REG_15 ? _GEN_758 : _GEN_342; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_839 = REG_15 ? _GEN_759 : _GEN_343; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_840 = REG_15 ? _GEN_760 : _GEN_344; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_841 = REG_15 ? _GEN_761 : _GEN_345; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_842 = REG_15 ? _GEN_762 : _GEN_346; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_843 = REG_15 ? _GEN_763 : _GEN_347; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_844 = REG_15 ? _GEN_764 : _GEN_348; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_845 = REG_15 ? _GEN_765 : _GEN_349; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_846 = REG_15 ? _GEN_766 : _GEN_350; // @[BranchTargetBuffer.scala 137:35]
  wire [31:0] _WIRE_27_0_target = btb_target_0_MPORT_17_data;
  wire [31:0] _GEN_864 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _WIRE_27_0_target : 32'h0; // @[BranchTargetBuffer.scala 126:19 133:66 135:23]
  wire  _GEN_866 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_815 : _GEN_683; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_867 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_816 : _GEN_684; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_868 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_817 : _GEN_685; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_869 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_818 : _GEN_686; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_870 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_819 : _GEN_687; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_871 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_820 : _GEN_688; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_872 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_821 : _GEN_689; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_873 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_822 : _GEN_690; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_874 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_823 : _GEN_691; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_875 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_824 : _GEN_692; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_876 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_825 : _GEN_693; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_877 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_826 : _GEN_694; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_878 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_827 : _GEN_695; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_879 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_828 : _GEN_696; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_880 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_829 : _GEN_697; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_881 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_830 : _GEN_698; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_882 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_831 : _GEN_335; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_883 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_832 : _GEN_336; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_884 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_833 : _GEN_337; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_885 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_834 : _GEN_338; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_886 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_835 : _GEN_339; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_887 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_836 : _GEN_340; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_888 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_837 : _GEN_341; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_889 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_838 : _GEN_342; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_890 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_839 : _GEN_343; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_891 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_840 : _GEN_344; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_892 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_841 : _GEN_345; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_893 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_842 : _GEN_346; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_894 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_843 : _GEN_347; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_895 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_844 : _GEN_348; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_896 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_845 : _GEN_349; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_897 = REG_13_0 & _WIRE_27_0_tag == REG_14 ? _GEN_846 : _GEN_350; // @[BranchTargetBuffer.scala 133:66]
  reg [25:0] REG_17; // @[BranchTargetBuffer.scala 133:51]
  wire [25:0] _WIRE_27_1_tag = btb_tag_1_MPORT_20_data;
  reg  REG_18; // @[BranchTargetBuffer.scala 137:22]
  reg [3:0] REG_19; // @[BranchTargetBuffer.scala 138:33]
  wire  _GEN_917 = 4'h0 == REG_19 | _GEN_866; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_918 = 4'h1 == REG_19 | _GEN_867; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_919 = 4'h2 == REG_19 | _GEN_868; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_920 = 4'h3 == REG_19 | _GEN_869; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_921 = 4'h4 == REG_19 | _GEN_870; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_922 = 4'h5 == REG_19 | _GEN_871; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_923 = 4'h6 == REG_19 | _GEN_872; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_924 = 4'h7 == REG_19 | _GEN_873; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_925 = 4'h8 == REG_19 | _GEN_874; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_926 = 4'h9 == REG_19 | _GEN_875; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_927 = 4'ha == REG_19 | _GEN_876; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_928 = 4'hb == REG_19 | _GEN_877; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_929 = 4'hc == REG_19 | _GEN_878; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_930 = 4'hd == REG_19 | _GEN_879; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_931 = 4'he == REG_19 | _GEN_880; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_932 = 4'hf == REG_19 | _GEN_881; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_933 = 4'h0 == REG_19 ? 1'h0 : _GEN_882; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_934 = 4'h1 == REG_19 ? 1'h0 : _GEN_883; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_935 = 4'h2 == REG_19 ? 1'h0 : _GEN_884; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_936 = 4'h3 == REG_19 ? 1'h0 : _GEN_885; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_937 = 4'h4 == REG_19 ? 1'h0 : _GEN_886; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_938 = 4'h5 == REG_19 ? 1'h0 : _GEN_887; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_939 = 4'h6 == REG_19 ? 1'h0 : _GEN_888; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_940 = 4'h7 == REG_19 ? 1'h0 : _GEN_889; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_941 = 4'h8 == REG_19 ? 1'h0 : _GEN_890; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_942 = 4'h9 == REG_19 ? 1'h0 : _GEN_891; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_943 = 4'ha == REG_19 ? 1'h0 : _GEN_892; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_944 = 4'hb == REG_19 ? 1'h0 : _GEN_893; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_945 = 4'hc == REG_19 ? 1'h0 : _GEN_894; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_946 = 4'hd == REG_19 ? 1'h0 : _GEN_895; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_947 = 4'he == REG_19 ? 1'h0 : _GEN_896; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_948 = 4'hf == REG_19 ? 1'h0 : _GEN_897; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_997 = REG_18 ? _GEN_917 : _GEN_866; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_998 = REG_18 ? _GEN_918 : _GEN_867; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_999 = REG_18 ? _GEN_919 : _GEN_868; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1000 = REG_18 ? _GEN_920 : _GEN_869; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1001 = REG_18 ? _GEN_921 : _GEN_870; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1002 = REG_18 ? _GEN_922 : _GEN_871; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1003 = REG_18 ? _GEN_923 : _GEN_872; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1004 = REG_18 ? _GEN_924 : _GEN_873; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1005 = REG_18 ? _GEN_925 : _GEN_874; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1006 = REG_18 ? _GEN_926 : _GEN_875; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1007 = REG_18 ? _GEN_927 : _GEN_876; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1008 = REG_18 ? _GEN_928 : _GEN_877; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1009 = REG_18 ? _GEN_929 : _GEN_878; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1010 = REG_18 ? _GEN_930 : _GEN_879; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1011 = REG_18 ? _GEN_931 : _GEN_880; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1012 = REG_18 ? _GEN_932 : _GEN_881; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1013 = REG_18 ? _GEN_933 : _GEN_882; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1014 = REG_18 ? _GEN_934 : _GEN_883; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1015 = REG_18 ? _GEN_935 : _GEN_884; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1016 = REG_18 ? _GEN_936 : _GEN_885; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1017 = REG_18 ? _GEN_937 : _GEN_886; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1018 = REG_18 ? _GEN_938 : _GEN_887; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1019 = REG_18 ? _GEN_939 : _GEN_888; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1020 = REG_18 ? _GEN_940 : _GEN_889; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1021 = REG_18 ? _GEN_941 : _GEN_890; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1022 = REG_18 ? _GEN_942 : _GEN_891; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1023 = REG_18 ? _GEN_943 : _GEN_892; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1024 = REG_18 ? _GEN_944 : _GEN_893; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1025 = REG_18 ? _GEN_945 : _GEN_894; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1026 = REG_18 ? _GEN_946 : _GEN_895; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1027 = REG_18 ? _GEN_947 : _GEN_896; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1028 = REG_18 ? _GEN_948 : _GEN_897; // @[BranchTargetBuffer.scala 137:35]
  wire [31:0] _WIRE_27_1_target = btb_target_1_MPORT_21_data;
  wire [31:0] _GEN_1046 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _WIRE_27_1_target : _GEN_864; // @[BranchTargetBuffer.scala 133:66 135:23]
  wire  _GEN_1048 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_997 : _GEN_866; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1049 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_998 : _GEN_867; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1050 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_999 : _GEN_868; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1051 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1000 : _GEN_869; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1052 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1001 : _GEN_870; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1053 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1002 : _GEN_871; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1054 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1003 : _GEN_872; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1055 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1004 : _GEN_873; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1056 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1005 : _GEN_874; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1057 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1006 : _GEN_875; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1058 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1007 : _GEN_876; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1059 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1008 : _GEN_877; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1060 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1009 : _GEN_878; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1061 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1010 : _GEN_879; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1062 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1011 : _GEN_880; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1063 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1012 : _GEN_881; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1064 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1013 : _GEN_882; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1065 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1014 : _GEN_883; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1066 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1015 : _GEN_884; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1067 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1016 : _GEN_885; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1068 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1017 : _GEN_886; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1069 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1018 : _GEN_887; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1070 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1019 : _GEN_888; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1071 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1020 : _GEN_889; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1072 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1021 : _GEN_890; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1073 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1022 : _GEN_891; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1074 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1023 : _GEN_892; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1075 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1024 : _GEN_893; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1076 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1025 : _GEN_894; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1077 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1026 : _GEN_895; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1078 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1027 : _GEN_896; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1079 = REG_13_1 & _WIRE_27_1_tag == REG_17 ? _GEN_1028 : _GEN_897; // @[BranchTargetBuffer.scala 133:66]
  reg [25:0] REG_20; // @[BranchTargetBuffer.scala 133:51]
  wire [25:0] _WIRE_27_2_tag = btb_tag_2_MPORT_24_data;
  reg  REG_21; // @[BranchTargetBuffer.scala 137:22]
  reg [3:0] REG_22; // @[BranchTargetBuffer.scala 138:33]
  wire  _GEN_1099 = 4'h0 == REG_22 ? 1'h0 : _GEN_1048; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1100 = 4'h1 == REG_22 ? 1'h0 : _GEN_1049; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1101 = 4'h2 == REG_22 ? 1'h0 : _GEN_1050; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1102 = 4'h3 == REG_22 ? 1'h0 : _GEN_1051; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1103 = 4'h4 == REG_22 ? 1'h0 : _GEN_1052; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1104 = 4'h5 == REG_22 ? 1'h0 : _GEN_1053; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1105 = 4'h6 == REG_22 ? 1'h0 : _GEN_1054; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1106 = 4'h7 == REG_22 ? 1'h0 : _GEN_1055; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1107 = 4'h8 == REG_22 ? 1'h0 : _GEN_1056; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1108 = 4'h9 == REG_22 ? 1'h0 : _GEN_1057; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1109 = 4'ha == REG_22 ? 1'h0 : _GEN_1058; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1110 = 4'hb == REG_22 ? 1'h0 : _GEN_1059; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1111 = 4'hc == REG_22 ? 1'h0 : _GEN_1060; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1112 = 4'hd == REG_22 ? 1'h0 : _GEN_1061; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1113 = 4'he == REG_22 ? 1'h0 : _GEN_1062; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1114 = 4'hf == REG_22 ? 1'h0 : _GEN_1063; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3051 = 4'h0 == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3052 = 4'h1 == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3053 = 4'h2 == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3054 = 4'h3 == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3055 = 4'h4 == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3056 = 4'h5 == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3057 = 4'h6 == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3058 = 4'h7 == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3059 = 4'h8 == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3060 = 4'h9 == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3061 = 4'ha == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3062 = 4'hb == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3063 = 4'hc == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3064 = 4'hd == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3065 = 4'he == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3066 = 4'hf == REG_22; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1131 = _GEN_3051 | _GEN_715; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1132 = _GEN_3052 | _GEN_716; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1133 = _GEN_3053 | _GEN_717; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1134 = _GEN_3054 | _GEN_718; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1135 = _GEN_3055 | _GEN_719; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1136 = _GEN_3056 | _GEN_720; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1137 = _GEN_3057 | _GEN_721; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1138 = _GEN_3058 | _GEN_722; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1139 = _GEN_3059 | _GEN_723; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1140 = _GEN_3060 | _GEN_724; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1141 = _GEN_3061 | _GEN_725; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1142 = _GEN_3062 | _GEN_726; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1143 = _GEN_3063 | _GEN_727; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1144 = _GEN_3064 | _GEN_728; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1145 = _GEN_3065 | _GEN_729; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1146 = _GEN_3066 | _GEN_730; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1179 = REG_21 ? _GEN_1099 : _GEN_1048; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1180 = REG_21 ? _GEN_1100 : _GEN_1049; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1181 = REG_21 ? _GEN_1101 : _GEN_1050; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1182 = REG_21 ? _GEN_1102 : _GEN_1051; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1183 = REG_21 ? _GEN_1103 : _GEN_1052; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1184 = REG_21 ? _GEN_1104 : _GEN_1053; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1185 = REG_21 ? _GEN_1105 : _GEN_1054; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1186 = REG_21 ? _GEN_1106 : _GEN_1055; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1187 = REG_21 ? _GEN_1107 : _GEN_1056; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1188 = REG_21 ? _GEN_1108 : _GEN_1057; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1189 = REG_21 ? _GEN_1109 : _GEN_1058; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1190 = REG_21 ? _GEN_1110 : _GEN_1059; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1191 = REG_21 ? _GEN_1111 : _GEN_1060; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1192 = REG_21 ? _GEN_1112 : _GEN_1061; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1193 = REG_21 ? _GEN_1113 : _GEN_1062; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1194 = REG_21 ? _GEN_1114 : _GEN_1063; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1211 = REG_21 ? _GEN_1131 : _GEN_715; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1212 = REG_21 ? _GEN_1132 : _GEN_716; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1213 = REG_21 ? _GEN_1133 : _GEN_717; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1214 = REG_21 ? _GEN_1134 : _GEN_718; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1215 = REG_21 ? _GEN_1135 : _GEN_719; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1216 = REG_21 ? _GEN_1136 : _GEN_720; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1217 = REG_21 ? _GEN_1137 : _GEN_721; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1218 = REG_21 ? _GEN_1138 : _GEN_722; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1219 = REG_21 ? _GEN_1139 : _GEN_723; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1220 = REG_21 ? _GEN_1140 : _GEN_724; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1221 = REG_21 ? _GEN_1141 : _GEN_725; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1222 = REG_21 ? _GEN_1142 : _GEN_726; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1223 = REG_21 ? _GEN_1143 : _GEN_727; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1224 = REG_21 ? _GEN_1144 : _GEN_728; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1225 = REG_21 ? _GEN_1145 : _GEN_729; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1226 = REG_21 ? _GEN_1146 : _GEN_730; // @[BranchTargetBuffer.scala 137:35]
  wire [31:0] _WIRE_27_2_target = btb_target_2_MPORT_25_data;
  wire [31:0] _GEN_1228 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _WIRE_27_2_target : _GEN_1046; // @[BranchTargetBuffer.scala 133:66 135:23]
  wire  _GEN_1230 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1179 : _GEN_1048; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1231 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1180 : _GEN_1049; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1232 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1181 : _GEN_1050; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1233 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1182 : _GEN_1051; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1234 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1183 : _GEN_1052; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1235 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1184 : _GEN_1053; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1236 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1185 : _GEN_1054; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1237 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1186 : _GEN_1055; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1238 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1187 : _GEN_1056; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1239 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1188 : _GEN_1057; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1240 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1189 : _GEN_1058; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1241 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1190 : _GEN_1059; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1242 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1191 : _GEN_1060; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1243 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1192 : _GEN_1061; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1244 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1193 : _GEN_1062; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1245 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1194 : _GEN_1063; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1262 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1211 : _GEN_715; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1263 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1212 : _GEN_716; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1264 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1213 : _GEN_717; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1265 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1214 : _GEN_718; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1266 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1215 : _GEN_719; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1267 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1216 : _GEN_720; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1268 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1217 : _GEN_721; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1269 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1218 : _GEN_722; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1270 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1219 : _GEN_723; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1271 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1220 : _GEN_724; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1272 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1221 : _GEN_725; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1273 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1222 : _GEN_726; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1274 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1223 : _GEN_727; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1275 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1224 : _GEN_728; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1276 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1225 : _GEN_729; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1277 = REG_13_2 & _WIRE_27_2_tag == REG_20 ? _GEN_1226 : _GEN_730; // @[BranchTargetBuffer.scala 133:66]
  reg [25:0] REG_23; // @[BranchTargetBuffer.scala 133:51]
  wire [25:0] _WIRE_27_3_tag = btb_tag_3_MPORT_28_data;
  reg  REG_24; // @[BranchTargetBuffer.scala 137:22]
  reg [3:0] REG_25; // @[BranchTargetBuffer.scala 138:33]
  wire  _GEN_1281 = 4'h0 == REG_25 ? 1'h0 : _GEN_1230; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1282 = 4'h1 == REG_25 ? 1'h0 : _GEN_1231; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1283 = 4'h2 == REG_25 ? 1'h0 : _GEN_1232; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1284 = 4'h3 == REG_25 ? 1'h0 : _GEN_1233; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1285 = 4'h4 == REG_25 ? 1'h0 : _GEN_1234; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1286 = 4'h5 == REG_25 ? 1'h0 : _GEN_1235; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1287 = 4'h6 == REG_25 ? 1'h0 : _GEN_1236; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1288 = 4'h7 == REG_25 ? 1'h0 : _GEN_1237; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1289 = 4'h8 == REG_25 ? 1'h0 : _GEN_1238; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1290 = 4'h9 == REG_25 ? 1'h0 : _GEN_1239; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1291 = 4'ha == REG_25 ? 1'h0 : _GEN_1240; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1292 = 4'hb == REG_25 ? 1'h0 : _GEN_1241; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1293 = 4'hc == REG_25 ? 1'h0 : _GEN_1242; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1294 = 4'hd == REG_25 ? 1'h0 : _GEN_1243; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1295 = 4'he == REG_25 ? 1'h0 : _GEN_1244; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1296 = 4'hf == REG_25 ? 1'h0 : _GEN_1245; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1313 = 4'h0 == REG_25 ? 1'h0 : _GEN_1262; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1314 = 4'h1 == REG_25 ? 1'h0 : _GEN_1263; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1315 = 4'h2 == REG_25 ? 1'h0 : _GEN_1264; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1316 = 4'h3 == REG_25 ? 1'h0 : _GEN_1265; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1317 = 4'h4 == REG_25 ? 1'h0 : _GEN_1266; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1318 = 4'h5 == REG_25 ? 1'h0 : _GEN_1267; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1319 = 4'h6 == REG_25 ? 1'h0 : _GEN_1268; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1320 = 4'h7 == REG_25 ? 1'h0 : _GEN_1269; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1321 = 4'h8 == REG_25 ? 1'h0 : _GEN_1270; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1322 = 4'h9 == REG_25 ? 1'h0 : _GEN_1271; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1323 = 4'ha == REG_25 ? 1'h0 : _GEN_1272; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1324 = 4'hb == REG_25 ? 1'h0 : _GEN_1273; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1325 = 4'hc == REG_25 ? 1'h0 : _GEN_1274; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1326 = 4'hd == REG_25 ? 1'h0 : _GEN_1275; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1327 = 4'he == REG_25 ? 1'h0 : _GEN_1276; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1328 = 4'hf == REG_25 ? 1'h0 : _GEN_1277; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1361 = REG_24 ? _GEN_1281 : _GEN_1230; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1362 = REG_24 ? _GEN_1282 : _GEN_1231; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1363 = REG_24 ? _GEN_1283 : _GEN_1232; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1364 = REG_24 ? _GEN_1284 : _GEN_1233; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1365 = REG_24 ? _GEN_1285 : _GEN_1234; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1366 = REG_24 ? _GEN_1286 : _GEN_1235; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1367 = REG_24 ? _GEN_1287 : _GEN_1236; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1368 = REG_24 ? _GEN_1288 : _GEN_1237; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1369 = REG_24 ? _GEN_1289 : _GEN_1238; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1370 = REG_24 ? _GEN_1290 : _GEN_1239; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1371 = REG_24 ? _GEN_1291 : _GEN_1240; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1372 = REG_24 ? _GEN_1292 : _GEN_1241; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1373 = REG_24 ? _GEN_1293 : _GEN_1242; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1374 = REG_24 ? _GEN_1294 : _GEN_1243; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1375 = REG_24 ? _GEN_1295 : _GEN_1244; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1376 = REG_24 ? _GEN_1296 : _GEN_1245; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1393 = REG_24 ? _GEN_1313 : _GEN_1262; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1394 = REG_24 ? _GEN_1314 : _GEN_1263; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1395 = REG_24 ? _GEN_1315 : _GEN_1264; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1396 = REG_24 ? _GEN_1316 : _GEN_1265; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1397 = REG_24 ? _GEN_1317 : _GEN_1266; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1398 = REG_24 ? _GEN_1318 : _GEN_1267; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1399 = REG_24 ? _GEN_1319 : _GEN_1268; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1400 = REG_24 ? _GEN_1320 : _GEN_1269; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1401 = REG_24 ? _GEN_1321 : _GEN_1270; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1402 = REG_24 ? _GEN_1322 : _GEN_1271; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1403 = REG_24 ? _GEN_1323 : _GEN_1272; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1404 = REG_24 ? _GEN_1324 : _GEN_1273; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1405 = REG_24 ? _GEN_1325 : _GEN_1274; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1406 = REG_24 ? _GEN_1326 : _GEN_1275; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1407 = REG_24 ? _GEN_1327 : _GEN_1276; // @[BranchTargetBuffer.scala 137:35]
  wire  _GEN_1408 = REG_24 ? _GEN_1328 : _GEN_1277; // @[BranchTargetBuffer.scala 137:35]
  wire [31:0] _WIRE_27_3_target = btb_target_3_MPORT_29_data;
  wire  _GEN_1412 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1361 : _GEN_1230; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1413 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1362 : _GEN_1231; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1414 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1363 : _GEN_1232; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1415 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1364 : _GEN_1233; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1416 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1365 : _GEN_1234; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1417 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1366 : _GEN_1235; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1418 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1367 : _GEN_1236; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1419 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1368 : _GEN_1237; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1420 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1369 : _GEN_1238; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1421 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1370 : _GEN_1239; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1422 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1371 : _GEN_1240; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1423 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1372 : _GEN_1241; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1424 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1373 : _GEN_1242; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1425 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1374 : _GEN_1243; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1426 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1375 : _GEN_1244; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1427 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1376 : _GEN_1245; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1444 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1393 : _GEN_1262; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1445 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1394 : _GEN_1263; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1446 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1395 : _GEN_1264; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1447 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1396 : _GEN_1265; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1448 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1397 : _GEN_1266; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1449 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1398 : _GEN_1267; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1450 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1399 : _GEN_1268; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1451 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1400 : _GEN_1269; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1452 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1401 : _GEN_1270; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1453 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1402 : _GEN_1271; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1454 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1403 : _GEN_1272; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1455 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1404 : _GEN_1273; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1456 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1405 : _GEN_1274; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1457 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1406 : _GEN_1275; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1458 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1407 : _GEN_1276; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1459 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _GEN_1408 : _GEN_1277; // @[BranchTargetBuffer.scala 133:66]
  wire  _GEN_1461 = 4'h1 == io_waddr ? plru0_1 : plru0_0; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1462 = 4'h2 == io_waddr ? plru0_2 : _GEN_1461; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1463 = 4'h3 == io_waddr ? plru0_3 : _GEN_1462; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1464 = 4'h4 == io_waddr ? plru0_4 : _GEN_1463; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1465 = 4'h5 == io_waddr ? plru0_5 : _GEN_1464; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1466 = 4'h6 == io_waddr ? plru0_6 : _GEN_1465; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1467 = 4'h7 == io_waddr ? plru0_7 : _GEN_1466; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1468 = 4'h8 == io_waddr ? plru0_8 : _GEN_1467; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1469 = 4'h9 == io_waddr ? plru0_9 : _GEN_1468; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1470 = 4'ha == io_waddr ? plru0_10 : _GEN_1469; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1471 = 4'hb == io_waddr ? plru0_11 : _GEN_1470; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1472 = 4'hc == io_waddr ? plru0_12 : _GEN_1471; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1473 = 4'hd == io_waddr ? plru0_13 : _GEN_1472; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1474 = 4'he == io_waddr ? plru0_14 : _GEN_1473; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1475 = 4'hf == io_waddr ? plru0_15 : _GEN_1474; // @[BranchTargetBuffer.scala 154:{45,45}]
  wire  _GEN_1477 = 4'h1 == io_waddr ? plru1_1 : plru1_0; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1478 = 4'h2 == io_waddr ? plru1_2 : _GEN_1477; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1479 = 4'h3 == io_waddr ? plru1_3 : _GEN_1478; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1480 = 4'h4 == io_waddr ? plru1_4 : _GEN_1479; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1481 = 4'h5 == io_waddr ? plru1_5 : _GEN_1480; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1482 = 4'h6 == io_waddr ? plru1_6 : _GEN_1481; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1483 = 4'h7 == io_waddr ? plru1_7 : _GEN_1482; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1484 = 4'h8 == io_waddr ? plru1_8 : _GEN_1483; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1485 = 4'h9 == io_waddr ? plru1_9 : _GEN_1484; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1486 = 4'ha == io_waddr ? plru1_10 : _GEN_1485; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1487 = 4'hb == io_waddr ? plru1_11 : _GEN_1486; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1488 = 4'hc == io_waddr ? plru1_12 : _GEN_1487; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1489 = 4'hd == io_waddr ? plru1_13 : _GEN_1488; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1490 = 4'he == io_waddr ? plru1_14 : _GEN_1489; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1491 = 4'hf == io_waddr ? plru1_15 : _GEN_1490; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1493 = 4'h1 == io_waddr ? plru2_1 : plru2_0; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1494 = 4'h2 == io_waddr ? plru2_2 : _GEN_1493; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1495 = 4'h3 == io_waddr ? plru2_3 : _GEN_1494; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1496 = 4'h4 == io_waddr ? plru2_4 : _GEN_1495; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1497 = 4'h5 == io_waddr ? plru2_5 : _GEN_1496; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1498 = 4'h6 == io_waddr ? plru2_6 : _GEN_1497; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1499 = 4'h7 == io_waddr ? plru2_7 : _GEN_1498; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1500 = 4'h8 == io_waddr ? plru2_8 : _GEN_1499; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1501 = 4'h9 == io_waddr ? plru2_9 : _GEN_1500; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1502 = 4'ha == io_waddr ? plru2_10 : _GEN_1501; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1503 = 4'hb == io_waddr ? plru2_11 : _GEN_1502; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1504 = 4'hc == io_waddr ? plru2_12 : _GEN_1503; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1505 = 4'hd == io_waddr ? plru2_13 : _GEN_1504; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1506 = 4'he == io_waddr ? plru2_14 : _GEN_1505; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _GEN_1507 = 4'hf == io_waddr ? plru2_15 : _GEN_1506; // @[BranchTargetBuffer.scala 154:{28,28}]
  wire  _T_145 = ~_GEN_1475 ? _GEN_1491 : _GEN_1507; // @[BranchTargetBuffer.scala 154:28]
  wire [1:0] replace_way = {_GEN_1475,_T_145}; // @[Cat.scala 30:58]
  reg  w_rvalid_0; // @[BranchTargetBuffer.scala 157:25]
  reg  w_rvalid_1; // @[BranchTargetBuffer.scala 157:25]
  reg  w_rvalid_2; // @[BranchTargetBuffer.scala 157:25]
  reg  w_rvalid_3; // @[BranchTargetBuffer.scala 157:25]
  reg [25:0] REG_26; // @[BranchTargetBuffer.scala 166:53]
  wire [25:0] w_rdata_0_tag = btb_tag_0_MPORT_32_data;
  reg [25:0] REG_27; // @[BranchTargetBuffer.scala 166:53]
  wire [25:0] w_rdata_1_tag = btb_tag_1_MPORT_35_data;
  wire [1:0] _GEN_1516 = w_rvalid_1 & w_rdata_1_tag == REG_27 ? 2'h1 : 2'h0; // @[BranchTargetBuffer.scala 166:65 168:13]
  reg [25:0] REG_28; // @[BranchTargetBuffer.scala 166:53]
  wire [25:0] w_rdata_2_tag = btb_tag_2_MPORT_38_data;
  wire [1:0] _GEN_1520 = w_rvalid_2 & w_rdata_2_tag == REG_28 ? 2'h2 : _GEN_1516; // @[BranchTargetBuffer.scala 166:65 168:13]
  reg [25:0] REG_29; // @[BranchTargetBuffer.scala 166:53]
  wire [25:0] w_rdata_3_tag = btb_tag_3_MPORT_41_data;
  wire  w_hit = w_rvalid_3 & w_rdata_3_tag == REG_29 | (w_rvalid_2 & w_rdata_2_tag == REG_28 | (w_rvalid_1 &
    w_rdata_1_tag == REG_27 | w_rvalid_0 & w_rdata_0_tag == REG_26)); // @[BranchTargetBuffer.scala 166:65 167:13]
  wire [1:0] w_way = w_rvalid_3 & w_rdata_3_tag == REG_29 ? 2'h3 : _GEN_1520; // @[BranchTargetBuffer.scala 166:65 168:13]
  reg  REG_30; // @[BranchTargetBuffer.scala 172:16]
  wire  _T_170 = w_way == 2'h0; // @[BranchTargetBuffer.scala 175:21]
  reg [3:0] REG_31; // @[BranchTargetBuffer.scala 176:35]
  reg [25:0] REG_32; // @[BranchTargetBuffer.scala 176:54]
  reg [3:0] REG_33; // @[BranchTargetBuffer.scala 177:38]
  reg [31:0] REG_34; // @[BranchTargetBuffer.scala 177:57]
  reg [3:0] REG_37; // @[BranchTargetBuffer.scala 179:33]
  wire  _GEN_3083 = 4'h0 == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1525 = 4'h0 == REG_37 | _GEN_1412; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3084 = 4'h1 == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1526 = 4'h1 == REG_37 | _GEN_1413; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3085 = 4'h2 == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1527 = 4'h2 == REG_37 | _GEN_1414; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3086 = 4'h3 == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1528 = 4'h3 == REG_37 | _GEN_1415; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3087 = 4'h4 == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1529 = 4'h4 == REG_37 | _GEN_1416; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3088 = 4'h5 == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1530 = 4'h5 == REG_37 | _GEN_1417; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3089 = 4'h6 == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1531 = 4'h6 == REG_37 | _GEN_1418; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3090 = 4'h7 == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1532 = 4'h7 == REG_37 | _GEN_1419; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3091 = 4'h8 == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1533 = 4'h8 == REG_37 | _GEN_1420; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3092 = 4'h9 == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1534 = 4'h9 == REG_37 | _GEN_1421; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3093 = 4'ha == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1535 = 4'ha == REG_37 | _GEN_1422; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3094 = 4'hb == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1536 = 4'hb == REG_37 | _GEN_1423; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3095 = 4'hc == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1537 = 4'hc == REG_37 | _GEN_1424; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3096 = 4'hd == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1538 = 4'hd == REG_37 | _GEN_1425; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3097 = 4'he == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1539 = 4'he == REG_37 | _GEN_1426; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3098 = 4'hf == REG_37; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1540 = 4'hf == REG_37 | _GEN_1427; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1541 = _GEN_3083 | _GEN_1064; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1542 = _GEN_3084 | _GEN_1065; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1543 = _GEN_3085 | _GEN_1066; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1544 = _GEN_3086 | _GEN_1067; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1545 = _GEN_3087 | _GEN_1068; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1546 = _GEN_3088 | _GEN_1069; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1547 = _GEN_3089 | _GEN_1070; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1548 = _GEN_3090 | _GEN_1071; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1549 = _GEN_3091 | _GEN_1072; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1550 = _GEN_3092 | _GEN_1073; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1551 = _GEN_3093 | _GEN_1074; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1552 = _GEN_3094 | _GEN_1075; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1553 = _GEN_3095 | _GEN_1076; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1554 = _GEN_3096 | _GEN_1077; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1555 = _GEN_3097 | _GEN_1078; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1556 = _GEN_3098 | _GEN_1079; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1614 = w_way == 2'h0 ? _GEN_1525 : _GEN_1412; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1615 = w_way == 2'h0 ? _GEN_1526 : _GEN_1413; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1616 = w_way == 2'h0 ? _GEN_1527 : _GEN_1414; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1617 = w_way == 2'h0 ? _GEN_1528 : _GEN_1415; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1618 = w_way == 2'h0 ? _GEN_1529 : _GEN_1416; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1619 = w_way == 2'h0 ? _GEN_1530 : _GEN_1417; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1620 = w_way == 2'h0 ? _GEN_1531 : _GEN_1418; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1621 = w_way == 2'h0 ? _GEN_1532 : _GEN_1419; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1622 = w_way == 2'h0 ? _GEN_1533 : _GEN_1420; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1623 = w_way == 2'h0 ? _GEN_1534 : _GEN_1421; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1624 = w_way == 2'h0 ? _GEN_1535 : _GEN_1422; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1625 = w_way == 2'h0 ? _GEN_1536 : _GEN_1423; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1626 = w_way == 2'h0 ? _GEN_1537 : _GEN_1424; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1627 = w_way == 2'h0 ? _GEN_1538 : _GEN_1425; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1628 = w_way == 2'h0 ? _GEN_1539 : _GEN_1426; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1629 = w_way == 2'h0 ? _GEN_1540 : _GEN_1427; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1630 = w_way == 2'h0 ? _GEN_1541 : _GEN_1064; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1631 = w_way == 2'h0 ? _GEN_1542 : _GEN_1065; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1632 = w_way == 2'h0 ? _GEN_1543 : _GEN_1066; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1633 = w_way == 2'h0 ? _GEN_1544 : _GEN_1067; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1634 = w_way == 2'h0 ? _GEN_1545 : _GEN_1068; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1635 = w_way == 2'h0 ? _GEN_1546 : _GEN_1069; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1636 = w_way == 2'h0 ? _GEN_1547 : _GEN_1070; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1637 = w_way == 2'h0 ? _GEN_1548 : _GEN_1071; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1638 = w_way == 2'h0 ? _GEN_1549 : _GEN_1072; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1639 = w_way == 2'h0 ? _GEN_1550 : _GEN_1073; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1640 = w_way == 2'h0 ? _GEN_1551 : _GEN_1074; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1641 = w_way == 2'h0 ? _GEN_1552 : _GEN_1075; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1642 = w_way == 2'h0 ? _GEN_1553 : _GEN_1076; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1643 = w_way == 2'h0 ? _GEN_1554 : _GEN_1077; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1644 = w_way == 2'h0 ? _GEN_1555 : _GEN_1078; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1645 = w_way == 2'h0 ? _GEN_1556 : _GEN_1079; // @[BranchTargetBuffer.scala 175:30]
  wire  _T_187 = w_way == 2'h1; // @[BranchTargetBuffer.scala 175:21]
  reg [3:0] REG_38; // @[BranchTargetBuffer.scala 176:35]
  reg [25:0] REG_39; // @[BranchTargetBuffer.scala 176:54]
  reg [3:0] REG_40; // @[BranchTargetBuffer.scala 177:38]
  reg [31:0] REG_41; // @[BranchTargetBuffer.scala 177:57]
  reg [3:0] REG_44; // @[BranchTargetBuffer.scala 179:33]
  wire  _GEN_1662 = 4'h0 == REG_44 | _GEN_1614; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1663 = 4'h1 == REG_44 | _GEN_1615; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1664 = 4'h2 == REG_44 | _GEN_1616; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1665 = 4'h3 == REG_44 | _GEN_1617; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1666 = 4'h4 == REG_44 | _GEN_1618; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1667 = 4'h5 == REG_44 | _GEN_1619; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1668 = 4'h6 == REG_44 | _GEN_1620; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1669 = 4'h7 == REG_44 | _GEN_1621; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1670 = 4'h8 == REG_44 | _GEN_1622; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1671 = 4'h9 == REG_44 | _GEN_1623; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1672 = 4'ha == REG_44 | _GEN_1624; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1673 = 4'hb == REG_44 | _GEN_1625; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1674 = 4'hc == REG_44 | _GEN_1626; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1675 = 4'hd == REG_44 | _GEN_1627; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1676 = 4'he == REG_44 | _GEN_1628; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1677 = 4'hf == REG_44 | _GEN_1629; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1678 = 4'h0 == REG_44 ? 1'h0 : _GEN_1630; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1679 = 4'h1 == REG_44 ? 1'h0 : _GEN_1631; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1680 = 4'h2 == REG_44 ? 1'h0 : _GEN_1632; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1681 = 4'h3 == REG_44 ? 1'h0 : _GEN_1633; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1682 = 4'h4 == REG_44 ? 1'h0 : _GEN_1634; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1683 = 4'h5 == REG_44 ? 1'h0 : _GEN_1635; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1684 = 4'h6 == REG_44 ? 1'h0 : _GEN_1636; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1685 = 4'h7 == REG_44 ? 1'h0 : _GEN_1637; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1686 = 4'h8 == REG_44 ? 1'h0 : _GEN_1638; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1687 = 4'h9 == REG_44 ? 1'h0 : _GEN_1639; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1688 = 4'ha == REG_44 ? 1'h0 : _GEN_1640; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1689 = 4'hb == REG_44 ? 1'h0 : _GEN_1641; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1690 = 4'hc == REG_44 ? 1'h0 : _GEN_1642; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1691 = 4'hd == REG_44 ? 1'h0 : _GEN_1643; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1692 = 4'he == REG_44 ? 1'h0 : _GEN_1644; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1693 = 4'hf == REG_44 ? 1'h0 : _GEN_1645; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1751 = w_way == 2'h1 ? _GEN_1662 : _GEN_1614; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1752 = w_way == 2'h1 ? _GEN_1663 : _GEN_1615; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1753 = w_way == 2'h1 ? _GEN_1664 : _GEN_1616; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1754 = w_way == 2'h1 ? _GEN_1665 : _GEN_1617; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1755 = w_way == 2'h1 ? _GEN_1666 : _GEN_1618; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1756 = w_way == 2'h1 ? _GEN_1667 : _GEN_1619; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1757 = w_way == 2'h1 ? _GEN_1668 : _GEN_1620; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1758 = w_way == 2'h1 ? _GEN_1669 : _GEN_1621; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1759 = w_way == 2'h1 ? _GEN_1670 : _GEN_1622; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1760 = w_way == 2'h1 ? _GEN_1671 : _GEN_1623; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1761 = w_way == 2'h1 ? _GEN_1672 : _GEN_1624; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1762 = w_way == 2'h1 ? _GEN_1673 : _GEN_1625; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1763 = w_way == 2'h1 ? _GEN_1674 : _GEN_1626; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1764 = w_way == 2'h1 ? _GEN_1675 : _GEN_1627; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1765 = w_way == 2'h1 ? _GEN_1676 : _GEN_1628; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1766 = w_way == 2'h1 ? _GEN_1677 : _GEN_1629; // @[BranchTargetBuffer.scala 175:30]
  wire  _T_204 = w_way == 2'h2; // @[BranchTargetBuffer.scala 175:21]
  reg [3:0] REG_45; // @[BranchTargetBuffer.scala 176:35]
  reg [25:0] REG_46; // @[BranchTargetBuffer.scala 176:54]
  reg [3:0] REG_47; // @[BranchTargetBuffer.scala 177:38]
  reg [31:0] REG_48; // @[BranchTargetBuffer.scala 177:57]
  reg [3:0] REG_51; // @[BranchTargetBuffer.scala 179:33]
  wire  _GEN_1799 = 4'h0 == REG_51 ? 1'h0 : _GEN_1751; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1800 = 4'h1 == REG_51 ? 1'h0 : _GEN_1752; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1801 = 4'h2 == REG_51 ? 1'h0 : _GEN_1753; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1802 = 4'h3 == REG_51 ? 1'h0 : _GEN_1754; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1803 = 4'h4 == REG_51 ? 1'h0 : _GEN_1755; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1804 = 4'h5 == REG_51 ? 1'h0 : _GEN_1756; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1805 = 4'h6 == REG_51 ? 1'h0 : _GEN_1757; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1806 = 4'h7 == REG_51 ? 1'h0 : _GEN_1758; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1807 = 4'h8 == REG_51 ? 1'h0 : _GEN_1759; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1808 = 4'h9 == REG_51 ? 1'h0 : _GEN_1760; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1809 = 4'ha == REG_51 ? 1'h0 : _GEN_1761; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1810 = 4'hb == REG_51 ? 1'h0 : _GEN_1762; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1811 = 4'hc == REG_51 ? 1'h0 : _GEN_1763; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1812 = 4'hd == REG_51 ? 1'h0 : _GEN_1764; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1813 = 4'he == REG_51 ? 1'h0 : _GEN_1765; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1814 = 4'hf == REG_51 ? 1'h0 : _GEN_1766; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3147 = 4'h0 == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3148 = 4'h1 == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3149 = 4'h2 == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3150 = 4'h3 == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3151 = 4'h4 == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3152 = 4'h5 == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3153 = 4'h6 == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3154 = 4'h7 == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3155 = 4'h8 == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3156 = 4'h9 == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3157 = 4'ha == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3158 = 4'hb == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3159 = 4'hc == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3160 = 4'hd == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3161 = 4'he == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3162 = 4'hf == REG_51; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_1831 = _GEN_3147 | _GEN_1444; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1832 = _GEN_3148 | _GEN_1445; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1833 = _GEN_3149 | _GEN_1446; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1834 = _GEN_3150 | _GEN_1447; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1835 = _GEN_3151 | _GEN_1448; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1836 = _GEN_3152 | _GEN_1449; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1837 = _GEN_3153 | _GEN_1450; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1838 = _GEN_3154 | _GEN_1451; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1839 = _GEN_3155 | _GEN_1452; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1840 = _GEN_3156 | _GEN_1453; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1841 = _GEN_3157 | _GEN_1454; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1842 = _GEN_3158 | _GEN_1455; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1843 = _GEN_3159 | _GEN_1456; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1844 = _GEN_3160 | _GEN_1457; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1845 = _GEN_3161 | _GEN_1458; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1846 = _GEN_3162 | _GEN_1459; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1888 = w_way == 2'h2 ? _GEN_1799 : _GEN_1751; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1889 = w_way == 2'h2 ? _GEN_1800 : _GEN_1752; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1890 = w_way == 2'h2 ? _GEN_1801 : _GEN_1753; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1891 = w_way == 2'h2 ? _GEN_1802 : _GEN_1754; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1892 = w_way == 2'h2 ? _GEN_1803 : _GEN_1755; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1893 = w_way == 2'h2 ? _GEN_1804 : _GEN_1756; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1894 = w_way == 2'h2 ? _GEN_1805 : _GEN_1757; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1895 = w_way == 2'h2 ? _GEN_1806 : _GEN_1758; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1896 = w_way == 2'h2 ? _GEN_1807 : _GEN_1759; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1897 = w_way == 2'h2 ? _GEN_1808 : _GEN_1760; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1898 = w_way == 2'h2 ? _GEN_1809 : _GEN_1761; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1899 = w_way == 2'h2 ? _GEN_1810 : _GEN_1762; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1900 = w_way == 2'h2 ? _GEN_1811 : _GEN_1763; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1901 = w_way == 2'h2 ? _GEN_1812 : _GEN_1764; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1902 = w_way == 2'h2 ? _GEN_1813 : _GEN_1765; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1903 = w_way == 2'h2 ? _GEN_1814 : _GEN_1766; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1920 = w_way == 2'h2 ? _GEN_1831 : _GEN_1444; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1921 = w_way == 2'h2 ? _GEN_1832 : _GEN_1445; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1922 = w_way == 2'h2 ? _GEN_1833 : _GEN_1446; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1923 = w_way == 2'h2 ? _GEN_1834 : _GEN_1447; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1924 = w_way == 2'h2 ? _GEN_1835 : _GEN_1448; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1925 = w_way == 2'h2 ? _GEN_1836 : _GEN_1449; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1926 = w_way == 2'h2 ? _GEN_1837 : _GEN_1450; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1927 = w_way == 2'h2 ? _GEN_1838 : _GEN_1451; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1928 = w_way == 2'h2 ? _GEN_1839 : _GEN_1452; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1929 = w_way == 2'h2 ? _GEN_1840 : _GEN_1453; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1930 = w_way == 2'h2 ? _GEN_1841 : _GEN_1454; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1931 = w_way == 2'h2 ? _GEN_1842 : _GEN_1455; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1932 = w_way == 2'h2 ? _GEN_1843 : _GEN_1456; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1933 = w_way == 2'h2 ? _GEN_1844 : _GEN_1457; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1934 = w_way == 2'h2 ? _GEN_1845 : _GEN_1458; // @[BranchTargetBuffer.scala 175:30]
  wire  _GEN_1935 = w_way == 2'h2 ? _GEN_1846 : _GEN_1459; // @[BranchTargetBuffer.scala 175:30]
  wire  _T_221 = w_way == 2'h3; // @[BranchTargetBuffer.scala 175:21]
  reg [3:0] REG_52; // @[BranchTargetBuffer.scala 176:35]
  reg [25:0] REG_53; // @[BranchTargetBuffer.scala 176:54]
  reg [3:0] REG_54; // @[BranchTargetBuffer.scala 177:38]
  reg [31:0] REG_55; // @[BranchTargetBuffer.scala 177:57]
  reg [3:0] REG_58; // @[BranchTargetBuffer.scala 179:33]
  wire  _GEN_1936 = 4'h0 == REG_58 ? 1'h0 : _GEN_1888; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1937 = 4'h1 == REG_58 ? 1'h0 : _GEN_1889; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1938 = 4'h2 == REG_58 ? 1'h0 : _GEN_1890; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1939 = 4'h3 == REG_58 ? 1'h0 : _GEN_1891; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1940 = 4'h4 == REG_58 ? 1'h0 : _GEN_1892; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1941 = 4'h5 == REG_58 ? 1'h0 : _GEN_1893; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1942 = 4'h6 == REG_58 ? 1'h0 : _GEN_1894; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1943 = 4'h7 == REG_58 ? 1'h0 : _GEN_1895; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1944 = 4'h8 == REG_58 ? 1'h0 : _GEN_1896; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1945 = 4'h9 == REG_58 ? 1'h0 : _GEN_1897; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1946 = 4'ha == REG_58 ? 1'h0 : _GEN_1898; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1947 = 4'hb == REG_58 ? 1'h0 : _GEN_1899; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1948 = 4'hc == REG_58 ? 1'h0 : _GEN_1900; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1949 = 4'hd == REG_58 ? 1'h0 : _GEN_1901; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1950 = 4'he == REG_58 ? 1'h0 : _GEN_1902; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1951 = 4'hf == REG_58 ? 1'h0 : _GEN_1903; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_1968 = 4'h0 == REG_58 ? 1'h0 : _GEN_1920; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1969 = 4'h1 == REG_58 ? 1'h0 : _GEN_1921; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1970 = 4'h2 == REG_58 ? 1'h0 : _GEN_1922; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1971 = 4'h3 == REG_58 ? 1'h0 : _GEN_1923; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1972 = 4'h4 == REG_58 ? 1'h0 : _GEN_1924; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1973 = 4'h5 == REG_58 ? 1'h0 : _GEN_1925; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1974 = 4'h6 == REG_58 ? 1'h0 : _GEN_1926; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1975 = 4'h7 == REG_58 ? 1'h0 : _GEN_1927; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1976 = 4'h8 == REG_58 ? 1'h0 : _GEN_1928; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1977 = 4'h9 == REG_58 ? 1'h0 : _GEN_1929; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1978 = 4'ha == REG_58 ? 1'h0 : _GEN_1930; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1979 = 4'hb == REG_58 ? 1'h0 : _GEN_1931; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1980 = 4'hc == REG_58 ? 1'h0 : _GEN_1932; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1981 = 4'hd == REG_58 ? 1'h0 : _GEN_1933; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1982 = 4'he == REG_58 ? 1'h0 : _GEN_1934; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_1983 = 4'hf == REG_58 ? 1'h0 : _GEN_1935; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _T_238 = replace_way == 2'h0; // @[BranchTargetBuffer.scala 187:27]
  reg [3:0] REG_59; // @[BranchTargetBuffer.scala 188:35]
  reg [25:0] REG_60; // @[BranchTargetBuffer.scala 188:54]
  reg [3:0] REG_61; // @[BranchTargetBuffer.scala 189:38]
  reg [31:0] REG_62; // @[BranchTargetBuffer.scala 189:57]
  reg [3:0] REG_65; // @[BranchTargetBuffer.scala 191:27]
  reg [3:0] REG_66; // @[BranchTargetBuffer.scala 192:33]
  wire  _GEN_3179 = 4'h0 == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2073 = 4'h0 == REG_66 | _GEN_1412; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3180 = 4'h1 == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2074 = 4'h1 == REG_66 | _GEN_1413; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3181 = 4'h2 == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2075 = 4'h2 == REG_66 | _GEN_1414; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3182 = 4'h3 == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2076 = 4'h3 == REG_66 | _GEN_1415; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3183 = 4'h4 == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2077 = 4'h4 == REG_66 | _GEN_1416; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3184 = 4'h5 == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2078 = 4'h5 == REG_66 | _GEN_1417; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3185 = 4'h6 == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2079 = 4'h6 == REG_66 | _GEN_1418; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3186 = 4'h7 == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2080 = 4'h7 == REG_66 | _GEN_1419; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3187 = 4'h8 == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2081 = 4'h8 == REG_66 | _GEN_1420; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3188 = 4'h9 == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2082 = 4'h9 == REG_66 | _GEN_1421; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3189 = 4'ha == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2083 = 4'ha == REG_66 | _GEN_1422; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3190 = 4'hb == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2084 = 4'hb == REG_66 | _GEN_1423; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3191 = 4'hc == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2085 = 4'hc == REG_66 | _GEN_1424; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3192 = 4'hd == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2086 = 4'hd == REG_66 | _GEN_1425; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3193 = 4'he == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2087 = 4'he == REG_66 | _GEN_1426; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3194 = 4'hf == REG_66; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2088 = 4'hf == REG_66 | _GEN_1427; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2089 = _GEN_3179 | _GEN_1064; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2090 = _GEN_3180 | _GEN_1065; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2091 = _GEN_3181 | _GEN_1066; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2092 = _GEN_3182 | _GEN_1067; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2093 = _GEN_3183 | _GEN_1068; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2094 = _GEN_3184 | _GEN_1069; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2095 = _GEN_3185 | _GEN_1070; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2096 = _GEN_3186 | _GEN_1071; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2097 = _GEN_3187 | _GEN_1072; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2098 = _GEN_3188 | _GEN_1073; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2099 = _GEN_3189 | _GEN_1074; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2100 = _GEN_3190 | _GEN_1075; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2101 = _GEN_3191 | _GEN_1076; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2102 = _GEN_3192 | _GEN_1077; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2103 = _GEN_3193 | _GEN_1078; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2104 = _GEN_3194 | _GEN_1079; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2163 = replace_way == 2'h0 ? _GEN_2073 : _GEN_1412; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2164 = replace_way == 2'h0 ? _GEN_2074 : _GEN_1413; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2165 = replace_way == 2'h0 ? _GEN_2075 : _GEN_1414; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2166 = replace_way == 2'h0 ? _GEN_2076 : _GEN_1415; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2167 = replace_way == 2'h0 ? _GEN_2077 : _GEN_1416; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2168 = replace_way == 2'h0 ? _GEN_2078 : _GEN_1417; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2169 = replace_way == 2'h0 ? _GEN_2079 : _GEN_1418; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2170 = replace_way == 2'h0 ? _GEN_2080 : _GEN_1419; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2171 = replace_way == 2'h0 ? _GEN_2081 : _GEN_1420; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2172 = replace_way == 2'h0 ? _GEN_2082 : _GEN_1421; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2173 = replace_way == 2'h0 ? _GEN_2083 : _GEN_1422; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2174 = replace_way == 2'h0 ? _GEN_2084 : _GEN_1423; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2175 = replace_way == 2'h0 ? _GEN_2085 : _GEN_1424; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2176 = replace_way == 2'h0 ? _GEN_2086 : _GEN_1425; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2177 = replace_way == 2'h0 ? _GEN_2087 : _GEN_1426; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2178 = replace_way == 2'h0 ? _GEN_2088 : _GEN_1427; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2179 = replace_way == 2'h0 ? _GEN_2089 : _GEN_1064; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2180 = replace_way == 2'h0 ? _GEN_2090 : _GEN_1065; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2181 = replace_way == 2'h0 ? _GEN_2091 : _GEN_1066; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2182 = replace_way == 2'h0 ? _GEN_2092 : _GEN_1067; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2183 = replace_way == 2'h0 ? _GEN_2093 : _GEN_1068; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2184 = replace_way == 2'h0 ? _GEN_2094 : _GEN_1069; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2185 = replace_way == 2'h0 ? _GEN_2095 : _GEN_1070; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2186 = replace_way == 2'h0 ? _GEN_2096 : _GEN_1071; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2187 = replace_way == 2'h0 ? _GEN_2097 : _GEN_1072; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2188 = replace_way == 2'h0 ? _GEN_2098 : _GEN_1073; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2189 = replace_way == 2'h0 ? _GEN_2099 : _GEN_1074; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2190 = replace_way == 2'h0 ? _GEN_2100 : _GEN_1075; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2191 = replace_way == 2'h0 ? _GEN_2101 : _GEN_1076; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2192 = replace_way == 2'h0 ? _GEN_2102 : _GEN_1077; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2193 = replace_way == 2'h0 ? _GEN_2103 : _GEN_1078; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2194 = replace_way == 2'h0 ? _GEN_2104 : _GEN_1079; // @[BranchTargetBuffer.scala 187:36]
  wire  _T_257 = replace_way == 2'h1; // @[BranchTargetBuffer.scala 187:27]
  reg [3:0] REG_67; // @[BranchTargetBuffer.scala 188:35]
  reg [25:0] REG_68; // @[BranchTargetBuffer.scala 188:54]
  reg [3:0] REG_69; // @[BranchTargetBuffer.scala 189:38]
  reg [31:0] REG_70; // @[BranchTargetBuffer.scala 189:57]
  reg [3:0] REG_73; // @[BranchTargetBuffer.scala 191:27]
  reg [3:0] REG_74; // @[BranchTargetBuffer.scala 192:33]
  wire  _GEN_2211 = 4'h0 == REG_74 | _GEN_2163; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2212 = 4'h1 == REG_74 | _GEN_2164; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2213 = 4'h2 == REG_74 | _GEN_2165; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2214 = 4'h3 == REG_74 | _GEN_2166; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2215 = 4'h4 == REG_74 | _GEN_2167; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2216 = 4'h5 == REG_74 | _GEN_2168; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2217 = 4'h6 == REG_74 | _GEN_2169; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2218 = 4'h7 == REG_74 | _GEN_2170; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2219 = 4'h8 == REG_74 | _GEN_2171; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2220 = 4'h9 == REG_74 | _GEN_2172; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2221 = 4'ha == REG_74 | _GEN_2173; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2222 = 4'hb == REG_74 | _GEN_2174; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2223 = 4'hc == REG_74 | _GEN_2175; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2224 = 4'hd == REG_74 | _GEN_2176; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2225 = 4'he == REG_74 | _GEN_2177; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2226 = 4'hf == REG_74 | _GEN_2178; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2227 = 4'h0 == REG_74 ? 1'h0 : _GEN_2179; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2228 = 4'h1 == REG_74 ? 1'h0 : _GEN_2180; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2229 = 4'h2 == REG_74 ? 1'h0 : _GEN_2181; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2230 = 4'h3 == REG_74 ? 1'h0 : _GEN_2182; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2231 = 4'h4 == REG_74 ? 1'h0 : _GEN_2183; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2232 = 4'h5 == REG_74 ? 1'h0 : _GEN_2184; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2233 = 4'h6 == REG_74 ? 1'h0 : _GEN_2185; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2234 = 4'h7 == REG_74 ? 1'h0 : _GEN_2186; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2235 = 4'h8 == REG_74 ? 1'h0 : _GEN_2187; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2236 = 4'h9 == REG_74 ? 1'h0 : _GEN_2188; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2237 = 4'ha == REG_74 ? 1'h0 : _GEN_2189; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2238 = 4'hb == REG_74 ? 1'h0 : _GEN_2190; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2239 = 4'hc == REG_74 ? 1'h0 : _GEN_2191; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2240 = 4'hd == REG_74 ? 1'h0 : _GEN_2192; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2241 = 4'he == REG_74 ? 1'h0 : _GEN_2193; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2242 = 4'hf == REG_74 ? 1'h0 : _GEN_2194; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2301 = replace_way == 2'h1 ? _GEN_2211 : _GEN_2163; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2302 = replace_way == 2'h1 ? _GEN_2212 : _GEN_2164; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2303 = replace_way == 2'h1 ? _GEN_2213 : _GEN_2165; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2304 = replace_way == 2'h1 ? _GEN_2214 : _GEN_2166; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2305 = replace_way == 2'h1 ? _GEN_2215 : _GEN_2167; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2306 = replace_way == 2'h1 ? _GEN_2216 : _GEN_2168; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2307 = replace_way == 2'h1 ? _GEN_2217 : _GEN_2169; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2308 = replace_way == 2'h1 ? _GEN_2218 : _GEN_2170; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2309 = replace_way == 2'h1 ? _GEN_2219 : _GEN_2171; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2310 = replace_way == 2'h1 ? _GEN_2220 : _GEN_2172; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2311 = replace_way == 2'h1 ? _GEN_2221 : _GEN_2173; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2312 = replace_way == 2'h1 ? _GEN_2222 : _GEN_2174; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2313 = replace_way == 2'h1 ? _GEN_2223 : _GEN_2175; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2314 = replace_way == 2'h1 ? _GEN_2224 : _GEN_2176; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2315 = replace_way == 2'h1 ? _GEN_2225 : _GEN_2177; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2316 = replace_way == 2'h1 ? _GEN_2226 : _GEN_2178; // @[BranchTargetBuffer.scala 187:36]
  wire  _T_276 = replace_way == 2'h2; // @[BranchTargetBuffer.scala 187:27]
  reg [3:0] REG_75; // @[BranchTargetBuffer.scala 188:35]
  reg [25:0] REG_76; // @[BranchTargetBuffer.scala 188:54]
  reg [3:0] REG_77; // @[BranchTargetBuffer.scala 189:38]
  reg [31:0] REG_78; // @[BranchTargetBuffer.scala 189:57]
  reg [3:0] REG_81; // @[BranchTargetBuffer.scala 191:27]
  reg [3:0] REG_82; // @[BranchTargetBuffer.scala 192:33]
  wire  _GEN_2349 = 4'h0 == REG_82 ? 1'h0 : _GEN_2301; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2350 = 4'h1 == REG_82 ? 1'h0 : _GEN_2302; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2351 = 4'h2 == REG_82 ? 1'h0 : _GEN_2303; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2352 = 4'h3 == REG_82 ? 1'h0 : _GEN_2304; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2353 = 4'h4 == REG_82 ? 1'h0 : _GEN_2305; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2354 = 4'h5 == REG_82 ? 1'h0 : _GEN_2306; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2355 = 4'h6 == REG_82 ? 1'h0 : _GEN_2307; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2356 = 4'h7 == REG_82 ? 1'h0 : _GEN_2308; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2357 = 4'h8 == REG_82 ? 1'h0 : _GEN_2309; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2358 = 4'h9 == REG_82 ? 1'h0 : _GEN_2310; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2359 = 4'ha == REG_82 ? 1'h0 : _GEN_2311; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2360 = 4'hb == REG_82 ? 1'h0 : _GEN_2312; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2361 = 4'hc == REG_82 ? 1'h0 : _GEN_2313; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2362 = 4'hd == REG_82 ? 1'h0 : _GEN_2314; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2363 = 4'he == REG_82 ? 1'h0 : _GEN_2315; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2364 = 4'hf == REG_82 ? 1'h0 : _GEN_2316; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_3243 = 4'h0 == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3244 = 4'h1 == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3245 = 4'h2 == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3246 = 4'h3 == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3247 = 4'h4 == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3248 = 4'h5 == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3249 = 4'h6 == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3250 = 4'h7 == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3251 = 4'h8 == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3252 = 4'h9 == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3253 = 4'ha == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3254 = 4'hb == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3255 = 4'hc == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3256 = 4'hd == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3257 = 4'he == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_3258 = 4'hf == REG_82; // @[BranchTargetBuffer.scala 116:{18,18}]
  wire  _GEN_2381 = _GEN_3243 | _GEN_1444; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2382 = _GEN_3244 | _GEN_1445; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2383 = _GEN_3245 | _GEN_1446; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2384 = _GEN_3246 | _GEN_1447; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2385 = _GEN_3247 | _GEN_1448; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2386 = _GEN_3248 | _GEN_1449; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2387 = _GEN_3249 | _GEN_1450; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2388 = _GEN_3250 | _GEN_1451; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2389 = _GEN_3251 | _GEN_1452; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2390 = _GEN_3252 | _GEN_1453; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2391 = _GEN_3253 | _GEN_1454; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2392 = _GEN_3254 | _GEN_1455; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2393 = _GEN_3255 | _GEN_1456; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2394 = _GEN_3256 | _GEN_1457; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2395 = _GEN_3257 | _GEN_1458; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2396 = _GEN_3258 | _GEN_1459; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2439 = replace_way == 2'h2 ? _GEN_2349 : _GEN_2301; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2440 = replace_way == 2'h2 ? _GEN_2350 : _GEN_2302; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2441 = replace_way == 2'h2 ? _GEN_2351 : _GEN_2303; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2442 = replace_way == 2'h2 ? _GEN_2352 : _GEN_2304; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2443 = replace_way == 2'h2 ? _GEN_2353 : _GEN_2305; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2444 = replace_way == 2'h2 ? _GEN_2354 : _GEN_2306; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2445 = replace_way == 2'h2 ? _GEN_2355 : _GEN_2307; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2446 = replace_way == 2'h2 ? _GEN_2356 : _GEN_2308; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2447 = replace_way == 2'h2 ? _GEN_2357 : _GEN_2309; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2448 = replace_way == 2'h2 ? _GEN_2358 : _GEN_2310; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2449 = replace_way == 2'h2 ? _GEN_2359 : _GEN_2311; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2450 = replace_way == 2'h2 ? _GEN_2360 : _GEN_2312; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2451 = replace_way == 2'h2 ? _GEN_2361 : _GEN_2313; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2452 = replace_way == 2'h2 ? _GEN_2362 : _GEN_2314; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2453 = replace_way == 2'h2 ? _GEN_2363 : _GEN_2315; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2454 = replace_way == 2'h2 ? _GEN_2364 : _GEN_2316; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2471 = replace_way == 2'h2 ? _GEN_2381 : _GEN_1444; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2472 = replace_way == 2'h2 ? _GEN_2382 : _GEN_1445; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2473 = replace_way == 2'h2 ? _GEN_2383 : _GEN_1446; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2474 = replace_way == 2'h2 ? _GEN_2384 : _GEN_1447; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2475 = replace_way == 2'h2 ? _GEN_2385 : _GEN_1448; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2476 = replace_way == 2'h2 ? _GEN_2386 : _GEN_1449; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2477 = replace_way == 2'h2 ? _GEN_2387 : _GEN_1450; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2478 = replace_way == 2'h2 ? _GEN_2388 : _GEN_1451; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2479 = replace_way == 2'h2 ? _GEN_2389 : _GEN_1452; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2480 = replace_way == 2'h2 ? _GEN_2390 : _GEN_1453; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2481 = replace_way == 2'h2 ? _GEN_2391 : _GEN_1454; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2482 = replace_way == 2'h2 ? _GEN_2392 : _GEN_1455; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2483 = replace_way == 2'h2 ? _GEN_2393 : _GEN_1456; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2484 = replace_way == 2'h2 ? _GEN_2394 : _GEN_1457; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2485 = replace_way == 2'h2 ? _GEN_2395 : _GEN_1458; // @[BranchTargetBuffer.scala 187:36]
  wire  _GEN_2486 = replace_way == 2'h2 ? _GEN_2396 : _GEN_1459; // @[BranchTargetBuffer.scala 187:36]
  wire  _T_295 = replace_way == 2'h3; // @[BranchTargetBuffer.scala 187:27]
  reg [3:0] REG_83; // @[BranchTargetBuffer.scala 188:35]
  reg [25:0] REG_84; // @[BranchTargetBuffer.scala 188:54]
  reg [3:0] REG_85; // @[BranchTargetBuffer.scala 189:38]
  reg [31:0] REG_86; // @[BranchTargetBuffer.scala 189:57]
  reg [3:0] REG_89; // @[BranchTargetBuffer.scala 191:27]
  reg [3:0] REG_90; // @[BranchTargetBuffer.scala 192:33]
  wire  _GEN_2487 = 4'h0 == REG_90 ? 1'h0 : _GEN_2439; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2488 = 4'h1 == REG_90 ? 1'h0 : _GEN_2440; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2489 = 4'h2 == REG_90 ? 1'h0 : _GEN_2441; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2490 = 4'h3 == REG_90 ? 1'h0 : _GEN_2442; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2491 = 4'h4 == REG_90 ? 1'h0 : _GEN_2443; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2492 = 4'h5 == REG_90 ? 1'h0 : _GEN_2444; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2493 = 4'h6 == REG_90 ? 1'h0 : _GEN_2445; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2494 = 4'h7 == REG_90 ? 1'h0 : _GEN_2446; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2495 = 4'h8 == REG_90 ? 1'h0 : _GEN_2447; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2496 = 4'h9 == REG_90 ? 1'h0 : _GEN_2448; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2497 = 4'ha == REG_90 ? 1'h0 : _GEN_2449; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2498 = 4'hb == REG_90 ? 1'h0 : _GEN_2450; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2499 = 4'hc == REG_90 ? 1'h0 : _GEN_2451; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2500 = 4'hd == REG_90 ? 1'h0 : _GEN_2452; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2501 = 4'he == REG_90 ? 1'h0 : _GEN_2453; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2502 = 4'hf == REG_90 ? 1'h0 : _GEN_2454; // @[BranchTargetBuffer.scala 114:{16,16}]
  wire  _GEN_2519 = 4'h0 == REG_90 ? 1'h0 : _GEN_2471; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2520 = 4'h1 == REG_90 ? 1'h0 : _GEN_2472; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2521 = 4'h2 == REG_90 ? 1'h0 : _GEN_2473; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2522 = 4'h3 == REG_90 ? 1'h0 : _GEN_2474; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2523 = 4'h4 == REG_90 ? 1'h0 : _GEN_2475; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2524 = 4'h5 == REG_90 ? 1'h0 : _GEN_2476; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2525 = 4'h6 == REG_90 ? 1'h0 : _GEN_2477; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2526 = 4'h7 == REG_90 ? 1'h0 : _GEN_2478; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2527 = 4'h8 == REG_90 ? 1'h0 : _GEN_2479; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2528 = 4'h9 == REG_90 ? 1'h0 : _GEN_2480; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2529 = 4'ha == REG_90 ? 1'h0 : _GEN_2481; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2530 = 4'hb == REG_90 ? 1'h0 : _GEN_2482; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2531 = 4'hc == REG_90 ? 1'h0 : _GEN_2483; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2532 = 4'hd == REG_90 ? 1'h0 : _GEN_2484; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2533 = 4'he == REG_90 ? 1'h0 : _GEN_2485; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2534 = 4'hf == REG_90 ? 1'h0 : _GEN_2486; // @[BranchTargetBuffer.scala 118:{18,18}]
  wire  _GEN_2627 = w_hit & _T_170; // @[BranchTargetBuffer.scala 173:18 90:30]
  wire  _GEN_2684 = w_hit & _T_187; // @[BranchTargetBuffer.scala 173:18 90:30]
  wire  _GEN_2693 = w_hit & _T_204; // @[BranchTargetBuffer.scala 173:18 90:30]
  wire  _GEN_2702 = w_hit & _T_221; // @[BranchTargetBuffer.scala 173:18 90:30]
  wire  _GEN_2711 = w_hit ? 1'h0 : _T_238; // @[BranchTargetBuffer.scala 173:18 90:30]
  wire  _GEN_2721 = w_hit ? 1'h0 : _T_257; // @[BranchTargetBuffer.scala 173:18 90:30]
  wire  _GEN_2731 = w_hit ? 1'h0 : _T_276; // @[BranchTargetBuffer.scala 173:18 90:30]
  wire  _GEN_2741 = w_hit ? 1'h0 : _T_295; // @[BranchTargetBuffer.scala 173:18 90:30]
//   assign btb_tag_0_MPORT_en = btb_tag_0_MPORT_en_pipe_0;
  assign btb_tag_0_MPORT_addr = btb_tag_0_MPORT_addr_pipe_0;
  assign btb_tag_0_MPORT_data = btb_tag_0[btb_tag_0_MPORT_addr]; // @[BranchTargetBuffer.scala 90:30]
//   assign btb_tag_0_MPORT_16_en = btb_tag_0_MPORT_16_en_pipe_0;
  assign btb_tag_0_MPORT_16_addr = btb_tag_0_MPORT_16_addr_pipe_0;
  assign btb_tag_0_MPORT_16_data = btb_tag_0[btb_tag_0_MPORT_16_addr]; // @[BranchTargetBuffer.scala 90:30]
//   assign btb_tag_0_MPORT_32_en = btb_tag_0_MPORT_32_en_pipe_0;
  assign btb_tag_0_MPORT_32_addr = btb_tag_0_MPORT_32_addr_pipe_0;
  assign btb_tag_0_MPORT_32_data = btb_tag_0[btb_tag_0_MPORT_32_addr]; // @[BranchTargetBuffer.scala 90:30]
  assign btb_tag_0_MPORT_44_data = REG_32;
  assign btb_tag_0_MPORT_44_addr = REG_31;
  assign btb_tag_0_MPORT_44_mask = 1'h1;
  assign btb_tag_0_MPORT_44_en = REG_30 & _GEN_2627;
  assign btb_tag_0_MPORT_56_data = REG_60;
  assign btb_tag_0_MPORT_56_addr = REG_59;
  assign btb_tag_0_MPORT_56_mask = 1'h1;
  assign btb_tag_0_MPORT_56_en = REG_30 & _GEN_2711;
  assign btb_tag_0_MPORT_72_data = 26'h0;
  assign btb_tag_0_MPORT_72_addr = 4'h0;
  assign btb_tag_0_MPORT_72_mask = 1'h1;
  assign btb_tag_0_MPORT_72_en = reset;
  assign btb_tag_0_MPORT_76_data = 26'h0;
  assign btb_tag_0_MPORT_76_addr = 4'h1;
  assign btb_tag_0_MPORT_76_mask = 1'h1;
  assign btb_tag_0_MPORT_76_en = reset;
  assign btb_tag_0_MPORT_80_data = 26'h0;
  assign btb_tag_0_MPORT_80_addr = 4'h2;
  assign btb_tag_0_MPORT_80_mask = 1'h1;
  assign btb_tag_0_MPORT_80_en = reset;
  assign btb_tag_0_MPORT_84_data = 26'h0;
  assign btb_tag_0_MPORT_84_addr = 4'h3;
  assign btb_tag_0_MPORT_84_mask = 1'h1;
  assign btb_tag_0_MPORT_84_en = reset;
  assign btb_tag_0_MPORT_88_data = 26'h0;
  assign btb_tag_0_MPORT_88_addr = 4'h4;
  assign btb_tag_0_MPORT_88_mask = 1'h1;
  assign btb_tag_0_MPORT_88_en = reset;
  assign btb_tag_0_MPORT_92_data = 26'h0;
  assign btb_tag_0_MPORT_92_addr = 4'h5;
  assign btb_tag_0_MPORT_92_mask = 1'h1;
  assign btb_tag_0_MPORT_92_en = reset;
  assign btb_tag_0_MPORT_96_data = 26'h0;
  assign btb_tag_0_MPORT_96_addr = 4'h6;
  assign btb_tag_0_MPORT_96_mask = 1'h1;
  assign btb_tag_0_MPORT_96_en = reset;
  assign btb_tag_0_MPORT_100_data = 26'h0;
  assign btb_tag_0_MPORT_100_addr = 4'h7;
  assign btb_tag_0_MPORT_100_mask = 1'h1;
  assign btb_tag_0_MPORT_100_en = reset;
  assign btb_tag_0_MPORT_104_data = 26'h0;
  assign btb_tag_0_MPORT_104_addr = 4'h8;
  assign btb_tag_0_MPORT_104_mask = 1'h1;
  assign btb_tag_0_MPORT_104_en = reset;
  assign btb_tag_0_MPORT_108_data = 26'h0;
  assign btb_tag_0_MPORT_108_addr = 4'h9;
  assign btb_tag_0_MPORT_108_mask = 1'h1;
  assign btb_tag_0_MPORT_108_en = reset;
  assign btb_tag_0_MPORT_112_data = 26'h0;
  assign btb_tag_0_MPORT_112_addr = 4'ha;
  assign btb_tag_0_MPORT_112_mask = 1'h1;
  assign btb_tag_0_MPORT_112_en = reset;
  assign btb_tag_0_MPORT_116_data = 26'h0;
  assign btb_tag_0_MPORT_116_addr = 4'hb;
  assign btb_tag_0_MPORT_116_mask = 1'h1;
  assign btb_tag_0_MPORT_116_en = reset;
  assign btb_tag_0_MPORT_120_data = 26'h0;
  assign btb_tag_0_MPORT_120_addr = 4'hc;
  assign btb_tag_0_MPORT_120_mask = 1'h1;
  assign btb_tag_0_MPORT_120_en = reset;
  assign btb_tag_0_MPORT_124_data = 26'h0;
  assign btb_tag_0_MPORT_124_addr = 4'hd;
  assign btb_tag_0_MPORT_124_mask = 1'h1;
  assign btb_tag_0_MPORT_124_en = reset;
  assign btb_tag_0_MPORT_128_data = 26'h0;
  assign btb_tag_0_MPORT_128_addr = 4'he;
  assign btb_tag_0_MPORT_128_mask = 1'h1;
  assign btb_tag_0_MPORT_128_en = reset;
  assign btb_tag_0_MPORT_132_data = 26'h0;
  assign btb_tag_0_MPORT_132_addr = 4'hf;
  assign btb_tag_0_MPORT_132_mask = 1'h1;
  assign btb_tag_0_MPORT_132_en = reset;
//   assign btb_tag_1_MPORT_4_en = btb_tag_1_MPORT_4_en_pipe_0;
  assign btb_tag_1_MPORT_4_addr = btb_tag_1_MPORT_4_addr_pipe_0;
  assign btb_tag_1_MPORT_4_data = btb_tag_1[btb_tag_1_MPORT_4_addr]; // @[BranchTargetBuffer.scala 90:30]
//   assign btb_tag_1_MPORT_20_en = btb_tag_1_MPORT_20_en_pipe_0;
  assign btb_tag_1_MPORT_20_addr = btb_tag_1_MPORT_20_addr_pipe_0;
  assign btb_tag_1_MPORT_20_data = btb_tag_1[btb_tag_1_MPORT_20_addr]; // @[BranchTargetBuffer.scala 90:30]
//   assign btb_tag_1_MPORT_35_en = btb_tag_1_MPORT_35_en_pipe_0;
  assign btb_tag_1_MPORT_35_addr = btb_tag_1_MPORT_35_addr_pipe_0;
  assign btb_tag_1_MPORT_35_data = btb_tag_1[btb_tag_1_MPORT_35_addr]; // @[BranchTargetBuffer.scala 90:30]
  assign btb_tag_1_MPORT_47_data = REG_39;
  assign btb_tag_1_MPORT_47_addr = REG_38;
  assign btb_tag_1_MPORT_47_mask = 1'h1;
  assign btb_tag_1_MPORT_47_en = REG_30 & _GEN_2684;
  assign btb_tag_1_MPORT_60_data = REG_68;
  assign btb_tag_1_MPORT_60_addr = REG_67;
  assign btb_tag_1_MPORT_60_mask = 1'h1;
  assign btb_tag_1_MPORT_60_en = REG_30 & _GEN_2721;
  assign btb_tag_1_MPORT_136_data = 26'h0;
  assign btb_tag_1_MPORT_136_addr = 4'h0;
  assign btb_tag_1_MPORT_136_mask = 1'h1;
  assign btb_tag_1_MPORT_136_en = reset;
  assign btb_tag_1_MPORT_140_data = 26'h0;
  assign btb_tag_1_MPORT_140_addr = 4'h1;
  assign btb_tag_1_MPORT_140_mask = 1'h1;
  assign btb_tag_1_MPORT_140_en = reset;
  assign btb_tag_1_MPORT_144_data = 26'h0;
  assign btb_tag_1_MPORT_144_addr = 4'h2;
  assign btb_tag_1_MPORT_144_mask = 1'h1;
  assign btb_tag_1_MPORT_144_en = reset;
  assign btb_tag_1_MPORT_148_data = 26'h0;
  assign btb_tag_1_MPORT_148_addr = 4'h3;
  assign btb_tag_1_MPORT_148_mask = 1'h1;
  assign btb_tag_1_MPORT_148_en = reset;
  assign btb_tag_1_MPORT_152_data = 26'h0;
  assign btb_tag_1_MPORT_152_addr = 4'h4;
  assign btb_tag_1_MPORT_152_mask = 1'h1;
  assign btb_tag_1_MPORT_152_en = reset;
  assign btb_tag_1_MPORT_156_data = 26'h0;
  assign btb_tag_1_MPORT_156_addr = 4'h5;
  assign btb_tag_1_MPORT_156_mask = 1'h1;
  assign btb_tag_1_MPORT_156_en = reset;
  assign btb_tag_1_MPORT_160_data = 26'h0;
  assign btb_tag_1_MPORT_160_addr = 4'h6;
  assign btb_tag_1_MPORT_160_mask = 1'h1;
  assign btb_tag_1_MPORT_160_en = reset;
  assign btb_tag_1_MPORT_164_data = 26'h0;
  assign btb_tag_1_MPORT_164_addr = 4'h7;
  assign btb_tag_1_MPORT_164_mask = 1'h1;
  assign btb_tag_1_MPORT_164_en = reset;
  assign btb_tag_1_MPORT_168_data = 26'h0;
  assign btb_tag_1_MPORT_168_addr = 4'h8;
  assign btb_tag_1_MPORT_168_mask = 1'h1;
  assign btb_tag_1_MPORT_168_en = reset;
  assign btb_tag_1_MPORT_172_data = 26'h0;
  assign btb_tag_1_MPORT_172_addr = 4'h9;
  assign btb_tag_1_MPORT_172_mask = 1'h1;
  assign btb_tag_1_MPORT_172_en = reset;
  assign btb_tag_1_MPORT_176_data = 26'h0;
  assign btb_tag_1_MPORT_176_addr = 4'ha;
  assign btb_tag_1_MPORT_176_mask = 1'h1;
  assign btb_tag_1_MPORT_176_en = reset;
  assign btb_tag_1_MPORT_180_data = 26'h0;
  assign btb_tag_1_MPORT_180_addr = 4'hb;
  assign btb_tag_1_MPORT_180_mask = 1'h1;
  assign btb_tag_1_MPORT_180_en = reset;
  assign btb_tag_1_MPORT_184_data = 26'h0;
  assign btb_tag_1_MPORT_184_addr = 4'hc;
  assign btb_tag_1_MPORT_184_mask = 1'h1;
  assign btb_tag_1_MPORT_184_en = reset;
  assign btb_tag_1_MPORT_188_data = 26'h0;
  assign btb_tag_1_MPORT_188_addr = 4'hd;
  assign btb_tag_1_MPORT_188_mask = 1'h1;
  assign btb_tag_1_MPORT_188_en = reset;
  assign btb_tag_1_MPORT_192_data = 26'h0;
  assign btb_tag_1_MPORT_192_addr = 4'he;
  assign btb_tag_1_MPORT_192_mask = 1'h1;
  assign btb_tag_1_MPORT_192_en = reset;
  assign btb_tag_1_MPORT_196_data = 26'h0;
  assign btb_tag_1_MPORT_196_addr = 4'hf;
  assign btb_tag_1_MPORT_196_mask = 1'h1;
  assign btb_tag_1_MPORT_196_en = reset;
//   assign btb_tag_2_MPORT_8_en = btb_tag_2_MPORT_8_en_pipe_0;
  assign btb_tag_2_MPORT_8_addr = btb_tag_2_MPORT_8_addr_pipe_0;
  assign btb_tag_2_MPORT_8_data = btb_tag_2[btb_tag_2_MPORT_8_addr]; // @[BranchTargetBuffer.scala 90:30]
//   assign btb_tag_2_MPORT_24_en = btb_tag_2_MPORT_24_en_pipe_0;
  assign btb_tag_2_MPORT_24_addr = btb_tag_2_MPORT_24_addr_pipe_0;
  assign btb_tag_2_MPORT_24_data = btb_tag_2[btb_tag_2_MPORT_24_addr]; // @[BranchTargetBuffer.scala 90:30]
//   assign btb_tag_2_MPORT_38_en = btb_tag_2_MPORT_38_en_pipe_0;
  assign btb_tag_2_MPORT_38_addr = btb_tag_2_MPORT_38_addr_pipe_0;
  assign btb_tag_2_MPORT_38_data = btb_tag_2[btb_tag_2_MPORT_38_addr]; // @[BranchTargetBuffer.scala 90:30]
  assign btb_tag_2_MPORT_50_data = REG_46;
  assign btb_tag_2_MPORT_50_addr = REG_45;
  assign btb_tag_2_MPORT_50_mask = 1'h1;
  assign btb_tag_2_MPORT_50_en = REG_30 & _GEN_2693;
  assign btb_tag_2_MPORT_64_data = REG_76;
  assign btb_tag_2_MPORT_64_addr = REG_75;
  assign btb_tag_2_MPORT_64_mask = 1'h1;
  assign btb_tag_2_MPORT_64_en = REG_30 & _GEN_2731;
  assign btb_tag_2_MPORT_200_data = 26'h0;
  assign btb_tag_2_MPORT_200_addr = 4'h0;
  assign btb_tag_2_MPORT_200_mask = 1'h1;
  assign btb_tag_2_MPORT_200_en = reset;
  assign btb_tag_2_MPORT_204_data = 26'h0;
  assign btb_tag_2_MPORT_204_addr = 4'h1;
  assign btb_tag_2_MPORT_204_mask = 1'h1;
  assign btb_tag_2_MPORT_204_en = reset;
  assign btb_tag_2_MPORT_208_data = 26'h0;
  assign btb_tag_2_MPORT_208_addr = 4'h2;
  assign btb_tag_2_MPORT_208_mask = 1'h1;
  assign btb_tag_2_MPORT_208_en = reset;
  assign btb_tag_2_MPORT_212_data = 26'h0;
  assign btb_tag_2_MPORT_212_addr = 4'h3;
  assign btb_tag_2_MPORT_212_mask = 1'h1;
  assign btb_tag_2_MPORT_212_en = reset;
  assign btb_tag_2_MPORT_216_data = 26'h0;
  assign btb_tag_2_MPORT_216_addr = 4'h4;
  assign btb_tag_2_MPORT_216_mask = 1'h1;
  assign btb_tag_2_MPORT_216_en = reset;
  assign btb_tag_2_MPORT_220_data = 26'h0;
  assign btb_tag_2_MPORT_220_addr = 4'h5;
  assign btb_tag_2_MPORT_220_mask = 1'h1;
  assign btb_tag_2_MPORT_220_en = reset;
  assign btb_tag_2_MPORT_224_data = 26'h0;
  assign btb_tag_2_MPORT_224_addr = 4'h6;
  assign btb_tag_2_MPORT_224_mask = 1'h1;
  assign btb_tag_2_MPORT_224_en = reset;
  assign btb_tag_2_MPORT_228_data = 26'h0;
  assign btb_tag_2_MPORT_228_addr = 4'h7;
  assign btb_tag_2_MPORT_228_mask = 1'h1;
  assign btb_tag_2_MPORT_228_en = reset;
  assign btb_tag_2_MPORT_232_data = 26'h0;
  assign btb_tag_2_MPORT_232_addr = 4'h8;
  assign btb_tag_2_MPORT_232_mask = 1'h1;
  assign btb_tag_2_MPORT_232_en = reset;
  assign btb_tag_2_MPORT_236_data = 26'h0;
  assign btb_tag_2_MPORT_236_addr = 4'h9;
  assign btb_tag_2_MPORT_236_mask = 1'h1;
  assign btb_tag_2_MPORT_236_en = reset;
  assign btb_tag_2_MPORT_240_data = 26'h0;
  assign btb_tag_2_MPORT_240_addr = 4'ha;
  assign btb_tag_2_MPORT_240_mask = 1'h1;
  assign btb_tag_2_MPORT_240_en = reset;
  assign btb_tag_2_MPORT_244_data = 26'h0;
  assign btb_tag_2_MPORT_244_addr = 4'hb;
  assign btb_tag_2_MPORT_244_mask = 1'h1;
  assign btb_tag_2_MPORT_244_en = reset;
  assign btb_tag_2_MPORT_248_data = 26'h0;
  assign btb_tag_2_MPORT_248_addr = 4'hc;
  assign btb_tag_2_MPORT_248_mask = 1'h1;
  assign btb_tag_2_MPORT_248_en = reset;
  assign btb_tag_2_MPORT_252_data = 26'h0;
  assign btb_tag_2_MPORT_252_addr = 4'hd;
  assign btb_tag_2_MPORT_252_mask = 1'h1;
  assign btb_tag_2_MPORT_252_en = reset;
  assign btb_tag_2_MPORT_256_data = 26'h0;
  assign btb_tag_2_MPORT_256_addr = 4'he;
  assign btb_tag_2_MPORT_256_mask = 1'h1;
  assign btb_tag_2_MPORT_256_en = reset;
  assign btb_tag_2_MPORT_260_data = 26'h0;
  assign btb_tag_2_MPORT_260_addr = 4'hf;
  assign btb_tag_2_MPORT_260_mask = 1'h1;
  assign btb_tag_2_MPORT_260_en = reset;
//   assign btb_tag_3_MPORT_12_en = btb_tag_3_MPORT_12_en_pipe_0;
  assign btb_tag_3_MPORT_12_addr = btb_tag_3_MPORT_12_addr_pipe_0;
  assign btb_tag_3_MPORT_12_data = btb_tag_3[btb_tag_3_MPORT_12_addr]; // @[BranchTargetBuffer.scala 90:30]
//   assign btb_tag_3_MPORT_28_en = btb_tag_3_MPORT_28_en_pipe_0;
  assign btb_tag_3_MPORT_28_addr = btb_tag_3_MPORT_28_addr_pipe_0;
  assign btb_tag_3_MPORT_28_data = btb_tag_3[btb_tag_3_MPORT_28_addr]; // @[BranchTargetBuffer.scala 90:30]
//   assign btb_tag_3_MPORT_41_en = btb_tag_3_MPORT_41_en_pipe_0;
  assign btb_tag_3_MPORT_41_addr = btb_tag_3_MPORT_41_addr_pipe_0;
  assign btb_tag_3_MPORT_41_data = btb_tag_3[btb_tag_3_MPORT_41_addr]; // @[BranchTargetBuffer.scala 90:30]
  assign btb_tag_3_MPORT_53_data = REG_53;
  assign btb_tag_3_MPORT_53_addr = REG_52;
  assign btb_tag_3_MPORT_53_mask = 1'h1;
  assign btb_tag_3_MPORT_53_en = REG_30 & _GEN_2702;
  assign btb_tag_3_MPORT_68_data = REG_84;
  assign btb_tag_3_MPORT_68_addr = REG_83;
  assign btb_tag_3_MPORT_68_mask = 1'h1;
  assign btb_tag_3_MPORT_68_en = REG_30 & _GEN_2741;
  assign btb_tag_3_MPORT_264_data = 26'h0;
  assign btb_tag_3_MPORT_264_addr = 4'h0;
  assign btb_tag_3_MPORT_264_mask = 1'h1;
  assign btb_tag_3_MPORT_264_en = reset;
  assign btb_tag_3_MPORT_268_data = 26'h0;
  assign btb_tag_3_MPORT_268_addr = 4'h1;
  assign btb_tag_3_MPORT_268_mask = 1'h1;
  assign btb_tag_3_MPORT_268_en = reset;
  assign btb_tag_3_MPORT_272_data = 26'h0;
  assign btb_tag_3_MPORT_272_addr = 4'h2;
  assign btb_tag_3_MPORT_272_mask = 1'h1;
  assign btb_tag_3_MPORT_272_en = reset;
  assign btb_tag_3_MPORT_276_data = 26'h0;
  assign btb_tag_3_MPORT_276_addr = 4'h3;
  assign btb_tag_3_MPORT_276_mask = 1'h1;
  assign btb_tag_3_MPORT_276_en = reset;
  assign btb_tag_3_MPORT_280_data = 26'h0;
  assign btb_tag_3_MPORT_280_addr = 4'h4;
  assign btb_tag_3_MPORT_280_mask = 1'h1;
  assign btb_tag_3_MPORT_280_en = reset;
  assign btb_tag_3_MPORT_284_data = 26'h0;
  assign btb_tag_3_MPORT_284_addr = 4'h5;
  assign btb_tag_3_MPORT_284_mask = 1'h1;
  assign btb_tag_3_MPORT_284_en = reset;
  assign btb_tag_3_MPORT_288_data = 26'h0;
  assign btb_tag_3_MPORT_288_addr = 4'h6;
  assign btb_tag_3_MPORT_288_mask = 1'h1;
  assign btb_tag_3_MPORT_288_en = reset;
  assign btb_tag_3_MPORT_292_data = 26'h0;
  assign btb_tag_3_MPORT_292_addr = 4'h7;
  assign btb_tag_3_MPORT_292_mask = 1'h1;
  assign btb_tag_3_MPORT_292_en = reset;
  assign btb_tag_3_MPORT_296_data = 26'h0;
  assign btb_tag_3_MPORT_296_addr = 4'h8;
  assign btb_tag_3_MPORT_296_mask = 1'h1;
  assign btb_tag_3_MPORT_296_en = reset;
  assign btb_tag_3_MPORT_300_data = 26'h0;
  assign btb_tag_3_MPORT_300_addr = 4'h9;
  assign btb_tag_3_MPORT_300_mask = 1'h1;
  assign btb_tag_3_MPORT_300_en = reset;
  assign btb_tag_3_MPORT_304_data = 26'h0;
  assign btb_tag_3_MPORT_304_addr = 4'ha;
  assign btb_tag_3_MPORT_304_mask = 1'h1;
  assign btb_tag_3_MPORT_304_en = reset;
  assign btb_tag_3_MPORT_308_data = 26'h0;
  assign btb_tag_3_MPORT_308_addr = 4'hb;
  assign btb_tag_3_MPORT_308_mask = 1'h1;
  assign btb_tag_3_MPORT_308_en = reset;
  assign btb_tag_3_MPORT_312_data = 26'h0;
  assign btb_tag_3_MPORT_312_addr = 4'hc;
  assign btb_tag_3_MPORT_312_mask = 1'h1;
  assign btb_tag_3_MPORT_312_en = reset;
  assign btb_tag_3_MPORT_316_data = 26'h0;
  assign btb_tag_3_MPORT_316_addr = 4'hd;
  assign btb_tag_3_MPORT_316_mask = 1'h1;
  assign btb_tag_3_MPORT_316_en = reset;
  assign btb_tag_3_MPORT_320_data = 26'h0;
  assign btb_tag_3_MPORT_320_addr = 4'he;
  assign btb_tag_3_MPORT_320_mask = 1'h1;
  assign btb_tag_3_MPORT_320_en = reset;
  assign btb_tag_3_MPORT_324_data = 26'h0;
  assign btb_tag_3_MPORT_324_addr = 4'hf;
  assign btb_tag_3_MPORT_324_mask = 1'h1;
  assign btb_tag_3_MPORT_324_en = reset;
//   assign btb_target_0_MPORT_1_en = btb_target_0_MPORT_1_en_pipe_0;
  assign btb_target_0_MPORT_1_addr = btb_target_0_MPORT_1_addr_pipe_0;
  assign btb_target_0_MPORT_1_data = btb_target_0[btb_target_0_MPORT_1_addr]; // @[BranchTargetBuffer.scala 94:33]
//   assign btb_target_0_MPORT_17_en = btb_target_0_MPORT_17_en_pipe_0;
  assign btb_target_0_MPORT_17_addr = btb_target_0_MPORT_17_addr_pipe_0;
  assign btb_target_0_MPORT_17_data = btb_target_0[btb_target_0_MPORT_17_addr]; // @[BranchTargetBuffer.scala 94:33]
  assign btb_target_0_MPORT_45_data = REG_34;
  assign btb_target_0_MPORT_45_addr = REG_33;
  assign btb_target_0_MPORT_45_mask = 1'h1;
  assign btb_target_0_MPORT_45_en = REG_30 & _GEN_2627;
  assign btb_target_0_MPORT_57_data = REG_62;
  assign btb_target_0_MPORT_57_addr = REG_61;
  assign btb_target_0_MPORT_57_mask = 1'h1;
  assign btb_target_0_MPORT_57_en = REG_30 & _GEN_2711;
  assign btb_target_0_MPORT_73_data = 32'h0;
  assign btb_target_0_MPORT_73_addr = 4'h0;
  assign btb_target_0_MPORT_73_mask = 1'h1;
  assign btb_target_0_MPORT_73_en = reset;
  assign btb_target_0_MPORT_77_data = 32'h0;
  assign btb_target_0_MPORT_77_addr = 4'h1;
  assign btb_target_0_MPORT_77_mask = 1'h1;
  assign btb_target_0_MPORT_77_en = reset;
  assign btb_target_0_MPORT_81_data = 32'h0;
  assign btb_target_0_MPORT_81_addr = 4'h2;
  assign btb_target_0_MPORT_81_mask = 1'h1;
  assign btb_target_0_MPORT_81_en = reset;
  assign btb_target_0_MPORT_85_data = 32'h0;
  assign btb_target_0_MPORT_85_addr = 4'h3;
  assign btb_target_0_MPORT_85_mask = 1'h1;
  assign btb_target_0_MPORT_85_en = reset;
  assign btb_target_0_MPORT_89_data = 32'h0;
  assign btb_target_0_MPORT_89_addr = 4'h4;
  assign btb_target_0_MPORT_89_mask = 1'h1;
  assign btb_target_0_MPORT_89_en = reset;
  assign btb_target_0_MPORT_93_data = 32'h0;
  assign btb_target_0_MPORT_93_addr = 4'h5;
  assign btb_target_0_MPORT_93_mask = 1'h1;
  assign btb_target_0_MPORT_93_en = reset;
  assign btb_target_0_MPORT_97_data = 32'h0;
  assign btb_target_0_MPORT_97_addr = 4'h6;
  assign btb_target_0_MPORT_97_mask = 1'h1;
  assign btb_target_0_MPORT_97_en = reset;
  assign btb_target_0_MPORT_101_data = 32'h0;
  assign btb_target_0_MPORT_101_addr = 4'h7;
  assign btb_target_0_MPORT_101_mask = 1'h1;
  assign btb_target_0_MPORT_101_en = reset;
  assign btb_target_0_MPORT_105_data = 32'h0;
  assign btb_target_0_MPORT_105_addr = 4'h8;
  assign btb_target_0_MPORT_105_mask = 1'h1;
  assign btb_target_0_MPORT_105_en = reset;
  assign btb_target_0_MPORT_109_data = 32'h0;
  assign btb_target_0_MPORT_109_addr = 4'h9;
  assign btb_target_0_MPORT_109_mask = 1'h1;
  assign btb_target_0_MPORT_109_en = reset;
  assign btb_target_0_MPORT_113_data = 32'h0;
  assign btb_target_0_MPORT_113_addr = 4'ha;
  assign btb_target_0_MPORT_113_mask = 1'h1;
  assign btb_target_0_MPORT_113_en = reset;
  assign btb_target_0_MPORT_117_data = 32'h0;
  assign btb_target_0_MPORT_117_addr = 4'hb;
  assign btb_target_0_MPORT_117_mask = 1'h1;
  assign btb_target_0_MPORT_117_en = reset;
  assign btb_target_0_MPORT_121_data = 32'h0;
  assign btb_target_0_MPORT_121_addr = 4'hc;
  assign btb_target_0_MPORT_121_mask = 1'h1;
  assign btb_target_0_MPORT_121_en = reset;
  assign btb_target_0_MPORT_125_data = 32'h0;
  assign btb_target_0_MPORT_125_addr = 4'hd;
  assign btb_target_0_MPORT_125_mask = 1'h1;
  assign btb_target_0_MPORT_125_en = reset;
  assign btb_target_0_MPORT_129_data = 32'h0;
  assign btb_target_0_MPORT_129_addr = 4'he;
  assign btb_target_0_MPORT_129_mask = 1'h1;
  assign btb_target_0_MPORT_129_en = reset;
  assign btb_target_0_MPORT_133_data = 32'h0;
  assign btb_target_0_MPORT_133_addr = 4'hf;
  assign btb_target_0_MPORT_133_mask = 1'h1;
  assign btb_target_0_MPORT_133_en = reset;
//   assign btb_target_1_MPORT_5_en = btb_target_1_MPORT_5_en_pipe_0;
  assign btb_target_1_MPORT_5_addr = btb_target_1_MPORT_5_addr_pipe_0;
  assign btb_target_1_MPORT_5_data = btb_target_1[btb_target_1_MPORT_5_addr]; // @[BranchTargetBuffer.scala 94:33]
//   assign btb_target_1_MPORT_21_en = btb_target_1_MPORT_21_en_pipe_0;
  assign btb_target_1_MPORT_21_addr = btb_target_1_MPORT_21_addr_pipe_0;
  assign btb_target_1_MPORT_21_data = btb_target_1[btb_target_1_MPORT_21_addr]; // @[BranchTargetBuffer.scala 94:33]
  assign btb_target_1_MPORT_48_data = REG_41;
  assign btb_target_1_MPORT_48_addr = REG_40;
  assign btb_target_1_MPORT_48_mask = 1'h1;
  assign btb_target_1_MPORT_48_en = REG_30 & _GEN_2684;
  assign btb_target_1_MPORT_61_data = REG_70;
  assign btb_target_1_MPORT_61_addr = REG_69;
  assign btb_target_1_MPORT_61_mask = 1'h1;
  assign btb_target_1_MPORT_61_en = REG_30 & _GEN_2721;
  assign btb_target_1_MPORT_137_data = 32'h0;
  assign btb_target_1_MPORT_137_addr = 4'h0;
  assign btb_target_1_MPORT_137_mask = 1'h1;
  assign btb_target_1_MPORT_137_en = reset;
  assign btb_target_1_MPORT_141_data = 32'h0;
  assign btb_target_1_MPORT_141_addr = 4'h1;
  assign btb_target_1_MPORT_141_mask = 1'h1;
  assign btb_target_1_MPORT_141_en = reset;
  assign btb_target_1_MPORT_145_data = 32'h0;
  assign btb_target_1_MPORT_145_addr = 4'h2;
  assign btb_target_1_MPORT_145_mask = 1'h1;
  assign btb_target_1_MPORT_145_en = reset;
  assign btb_target_1_MPORT_149_data = 32'h0;
  assign btb_target_1_MPORT_149_addr = 4'h3;
  assign btb_target_1_MPORT_149_mask = 1'h1;
  assign btb_target_1_MPORT_149_en = reset;
  assign btb_target_1_MPORT_153_data = 32'h0;
  assign btb_target_1_MPORT_153_addr = 4'h4;
  assign btb_target_1_MPORT_153_mask = 1'h1;
  assign btb_target_1_MPORT_153_en = reset;
  assign btb_target_1_MPORT_157_data = 32'h0;
  assign btb_target_1_MPORT_157_addr = 4'h5;
  assign btb_target_1_MPORT_157_mask = 1'h1;
  assign btb_target_1_MPORT_157_en = reset;
  assign btb_target_1_MPORT_161_data = 32'h0;
  assign btb_target_1_MPORT_161_addr = 4'h6;
  assign btb_target_1_MPORT_161_mask = 1'h1;
  assign btb_target_1_MPORT_161_en = reset;
  assign btb_target_1_MPORT_165_data = 32'h0;
  assign btb_target_1_MPORT_165_addr = 4'h7;
  assign btb_target_1_MPORT_165_mask = 1'h1;
  assign btb_target_1_MPORT_165_en = reset;
  assign btb_target_1_MPORT_169_data = 32'h0;
  assign btb_target_1_MPORT_169_addr = 4'h8;
  assign btb_target_1_MPORT_169_mask = 1'h1;
  assign btb_target_1_MPORT_169_en = reset;
  assign btb_target_1_MPORT_173_data = 32'h0;
  assign btb_target_1_MPORT_173_addr = 4'h9;
  assign btb_target_1_MPORT_173_mask = 1'h1;
  assign btb_target_1_MPORT_173_en = reset;
  assign btb_target_1_MPORT_177_data = 32'h0;
  assign btb_target_1_MPORT_177_addr = 4'ha;
  assign btb_target_1_MPORT_177_mask = 1'h1;
  assign btb_target_1_MPORT_177_en = reset;
  assign btb_target_1_MPORT_181_data = 32'h0;
  assign btb_target_1_MPORT_181_addr = 4'hb;
  assign btb_target_1_MPORT_181_mask = 1'h1;
  assign btb_target_1_MPORT_181_en = reset;
  assign btb_target_1_MPORT_185_data = 32'h0;
  assign btb_target_1_MPORT_185_addr = 4'hc;
  assign btb_target_1_MPORT_185_mask = 1'h1;
  assign btb_target_1_MPORT_185_en = reset;
  assign btb_target_1_MPORT_189_data = 32'h0;
  assign btb_target_1_MPORT_189_addr = 4'hd;
  assign btb_target_1_MPORT_189_mask = 1'h1;
  assign btb_target_1_MPORT_189_en = reset;
  assign btb_target_1_MPORT_193_data = 32'h0;
  assign btb_target_1_MPORT_193_addr = 4'he;
  assign btb_target_1_MPORT_193_mask = 1'h1;
  assign btb_target_1_MPORT_193_en = reset;
  assign btb_target_1_MPORT_197_data = 32'h0;
  assign btb_target_1_MPORT_197_addr = 4'hf;
  assign btb_target_1_MPORT_197_mask = 1'h1;
  assign btb_target_1_MPORT_197_en = reset;
//   assign btb_target_2_MPORT_9_en = btb_target_2_MPORT_9_en_pipe_0;
  assign btb_target_2_MPORT_9_addr = btb_target_2_MPORT_9_addr_pipe_0;
  assign btb_target_2_MPORT_9_data = btb_target_2[btb_target_2_MPORT_9_addr]; // @[BranchTargetBuffer.scala 94:33]
//   assign btb_target_2_MPORT_25_en = btb_target_2_MPORT_25_en_pipe_0;
  assign btb_target_2_MPORT_25_addr = btb_target_2_MPORT_25_addr_pipe_0;
  assign btb_target_2_MPORT_25_data = btb_target_2[btb_target_2_MPORT_25_addr]; // @[BranchTargetBuffer.scala 94:33]
  assign btb_target_2_MPORT_51_data = REG_48;
  assign btb_target_2_MPORT_51_addr = REG_47;
  assign btb_target_2_MPORT_51_mask = 1'h1;
  assign btb_target_2_MPORT_51_en = REG_30 & _GEN_2693;
  assign btb_target_2_MPORT_65_data = REG_78;
  assign btb_target_2_MPORT_65_addr = REG_77;
  assign btb_target_2_MPORT_65_mask = 1'h1;
  assign btb_target_2_MPORT_65_en = REG_30 & _GEN_2731;
  assign btb_target_2_MPORT_201_data = 32'h0;
  assign btb_target_2_MPORT_201_addr = 4'h0;
  assign btb_target_2_MPORT_201_mask = 1'h1;
  assign btb_target_2_MPORT_201_en = reset;
  assign btb_target_2_MPORT_205_data = 32'h0;
  assign btb_target_2_MPORT_205_addr = 4'h1;
  assign btb_target_2_MPORT_205_mask = 1'h1;
  assign btb_target_2_MPORT_205_en = reset;
  assign btb_target_2_MPORT_209_data = 32'h0;
  assign btb_target_2_MPORT_209_addr = 4'h2;
  assign btb_target_2_MPORT_209_mask = 1'h1;
  assign btb_target_2_MPORT_209_en = reset;
  assign btb_target_2_MPORT_213_data = 32'h0;
  assign btb_target_2_MPORT_213_addr = 4'h3;
  assign btb_target_2_MPORT_213_mask = 1'h1;
  assign btb_target_2_MPORT_213_en = reset;
  assign btb_target_2_MPORT_217_data = 32'h0;
  assign btb_target_2_MPORT_217_addr = 4'h4;
  assign btb_target_2_MPORT_217_mask = 1'h1;
  assign btb_target_2_MPORT_217_en = reset;
  assign btb_target_2_MPORT_221_data = 32'h0;
  assign btb_target_2_MPORT_221_addr = 4'h5;
  assign btb_target_2_MPORT_221_mask = 1'h1;
  assign btb_target_2_MPORT_221_en = reset;
  assign btb_target_2_MPORT_225_data = 32'h0;
  assign btb_target_2_MPORT_225_addr = 4'h6;
  assign btb_target_2_MPORT_225_mask = 1'h1;
  assign btb_target_2_MPORT_225_en = reset;
  assign btb_target_2_MPORT_229_data = 32'h0;
  assign btb_target_2_MPORT_229_addr = 4'h7;
  assign btb_target_2_MPORT_229_mask = 1'h1;
  assign btb_target_2_MPORT_229_en = reset;
  assign btb_target_2_MPORT_233_data = 32'h0;
  assign btb_target_2_MPORT_233_addr = 4'h8;
  assign btb_target_2_MPORT_233_mask = 1'h1;
  assign btb_target_2_MPORT_233_en = reset;
  assign btb_target_2_MPORT_237_data = 32'h0;
  assign btb_target_2_MPORT_237_addr = 4'h9;
  assign btb_target_2_MPORT_237_mask = 1'h1;
  assign btb_target_2_MPORT_237_en = reset;
  assign btb_target_2_MPORT_241_data = 32'h0;
  assign btb_target_2_MPORT_241_addr = 4'ha;
  assign btb_target_2_MPORT_241_mask = 1'h1;
  assign btb_target_2_MPORT_241_en = reset;
  assign btb_target_2_MPORT_245_data = 32'h0;
  assign btb_target_2_MPORT_245_addr = 4'hb;
  assign btb_target_2_MPORT_245_mask = 1'h1;
  assign btb_target_2_MPORT_245_en = reset;
  assign btb_target_2_MPORT_249_data = 32'h0;
  assign btb_target_2_MPORT_249_addr = 4'hc;
  assign btb_target_2_MPORT_249_mask = 1'h1;
  assign btb_target_2_MPORT_249_en = reset;
  assign btb_target_2_MPORT_253_data = 32'h0;
  assign btb_target_2_MPORT_253_addr = 4'hd;
  assign btb_target_2_MPORT_253_mask = 1'h1;
  assign btb_target_2_MPORT_253_en = reset;
  assign btb_target_2_MPORT_257_data = 32'h0;
  assign btb_target_2_MPORT_257_addr = 4'he;
  assign btb_target_2_MPORT_257_mask = 1'h1;
  assign btb_target_2_MPORT_257_en = reset;
  assign btb_target_2_MPORT_261_data = 32'h0;
  assign btb_target_2_MPORT_261_addr = 4'hf;
  assign btb_target_2_MPORT_261_mask = 1'h1;
  assign btb_target_2_MPORT_261_en = reset;
//   assign btb_target_3_MPORT_13_en = btb_target_3_MPORT_13_en_pipe_0;
  assign btb_target_3_MPORT_13_addr = btb_target_3_MPORT_13_addr_pipe_0;
  assign btb_target_3_MPORT_13_data = btb_target_3[btb_target_3_MPORT_13_addr]; // @[BranchTargetBuffer.scala 94:33]
//   assign btb_target_3_MPORT_29_en = btb_target_3_MPORT_29_en_pipe_0;
  assign btb_target_3_MPORT_29_addr = btb_target_3_MPORT_29_addr_pipe_0;
  assign btb_target_3_MPORT_29_data = btb_target_3[btb_target_3_MPORT_29_addr]; // @[BranchTargetBuffer.scala 94:33]
  assign btb_target_3_MPORT_54_data = REG_55;
  assign btb_target_3_MPORT_54_addr = REG_54;
  assign btb_target_3_MPORT_54_mask = 1'h1;
  assign btb_target_3_MPORT_54_en = REG_30 & _GEN_2702;
  assign btb_target_3_MPORT_69_data = REG_86;
  assign btb_target_3_MPORT_69_addr = REG_85;
  assign btb_target_3_MPORT_69_mask = 1'h1;
  assign btb_target_3_MPORT_69_en = REG_30 & _GEN_2741;
  assign btb_target_3_MPORT_265_data = 32'h0;
  assign btb_target_3_MPORT_265_addr = 4'h0;
  assign btb_target_3_MPORT_265_mask = 1'h1;
  assign btb_target_3_MPORT_265_en = reset;
  assign btb_target_3_MPORT_269_data = 32'h0;
  assign btb_target_3_MPORT_269_addr = 4'h1;
  assign btb_target_3_MPORT_269_mask = 1'h1;
  assign btb_target_3_MPORT_269_en = reset;
  assign btb_target_3_MPORT_273_data = 32'h0;
  assign btb_target_3_MPORT_273_addr = 4'h2;
  assign btb_target_3_MPORT_273_mask = 1'h1;
  assign btb_target_3_MPORT_273_en = reset;
  assign btb_target_3_MPORT_277_data = 32'h0;
  assign btb_target_3_MPORT_277_addr = 4'h3;
  assign btb_target_3_MPORT_277_mask = 1'h1;
  assign btb_target_3_MPORT_277_en = reset;
  assign btb_target_3_MPORT_281_data = 32'h0;
  assign btb_target_3_MPORT_281_addr = 4'h4;
  assign btb_target_3_MPORT_281_mask = 1'h1;
  assign btb_target_3_MPORT_281_en = reset;
  assign btb_target_3_MPORT_285_data = 32'h0;
  assign btb_target_3_MPORT_285_addr = 4'h5;
  assign btb_target_3_MPORT_285_mask = 1'h1;
  assign btb_target_3_MPORT_285_en = reset;
  assign btb_target_3_MPORT_289_data = 32'h0;
  assign btb_target_3_MPORT_289_addr = 4'h6;
  assign btb_target_3_MPORT_289_mask = 1'h1;
  assign btb_target_3_MPORT_289_en = reset;
  assign btb_target_3_MPORT_293_data = 32'h0;
  assign btb_target_3_MPORT_293_addr = 4'h7;
  assign btb_target_3_MPORT_293_mask = 1'h1;
  assign btb_target_3_MPORT_293_en = reset;
  assign btb_target_3_MPORT_297_data = 32'h0;
  assign btb_target_3_MPORT_297_addr = 4'h8;
  assign btb_target_3_MPORT_297_mask = 1'h1;
  assign btb_target_3_MPORT_297_en = reset;
  assign btb_target_3_MPORT_301_data = 32'h0;
  assign btb_target_3_MPORT_301_addr = 4'h9;
  assign btb_target_3_MPORT_301_mask = 1'h1;
  assign btb_target_3_MPORT_301_en = reset;
  assign btb_target_3_MPORT_305_data = 32'h0;
  assign btb_target_3_MPORT_305_addr = 4'ha;
  assign btb_target_3_MPORT_305_mask = 1'h1;
  assign btb_target_3_MPORT_305_en = reset;
  assign btb_target_3_MPORT_309_data = 32'h0;
  assign btb_target_3_MPORT_309_addr = 4'hb;
  assign btb_target_3_MPORT_309_mask = 1'h1;
  assign btb_target_3_MPORT_309_en = reset;
  assign btb_target_3_MPORT_313_data = 32'h0;
  assign btb_target_3_MPORT_313_addr = 4'hc;
  assign btb_target_3_MPORT_313_mask = 1'h1;
  assign btb_target_3_MPORT_313_en = reset;
  assign btb_target_3_MPORT_317_data = 32'h0;
  assign btb_target_3_MPORT_317_addr = 4'hd;
  assign btb_target_3_MPORT_317_mask = 1'h1;
  assign btb_target_3_MPORT_317_en = reset;
  assign btb_target_3_MPORT_321_data = 32'h0;
  assign btb_target_3_MPORT_321_addr = 4'he;
  assign btb_target_3_MPORT_321_mask = 1'h1;
  assign btb_target_3_MPORT_321_en = reset;
  assign btb_target_3_MPORT_325_data = 32'h0;
  assign btb_target_3_MPORT_325_addr = 4'hf;
  assign btb_target_3_MPORT_325_mask = 1'h1;
  assign btb_target_3_MPORT_325_en = reset;
//   assign valid_0_MPORT_3_en = 1'h1;
  assign valid_0_MPORT_3_addr = io_raddr_0;
  assign valid_0_MPORT_3_data = valid_0[valid_0_MPORT_3_addr]; // @[BranchTargetBuffer.scala 102:20]
//   assign valid_0_MPORT_19_en = 1'h1;
  assign valid_0_MPORT_19_addr = io_raddr_1;
  assign valid_0_MPORT_19_data = valid_0[valid_0_MPORT_19_addr]; // @[BranchTargetBuffer.scala 102:20]
//   assign valid_0_MPORT_34_en = 1'h1;
  assign valid_0_MPORT_34_addr = io_waddr;
  assign valid_0_MPORT_34_data = valid_0[valid_0_MPORT_34_addr]; // @[BranchTargetBuffer.scala 102:20]
  assign valid_0_MPORT_59_data = 1'h1;
  assign valid_0_MPORT_59_addr = REG_65;
  assign valid_0_MPORT_59_mask = 1'h1;
  assign valid_0_MPORT_59_en = REG_30 & _GEN_2711;
  assign valid_0_MPORT_75_data = 1'h0;
  assign valid_0_MPORT_75_addr = 4'h0;
  assign valid_0_MPORT_75_mask = 1'h1;
  assign valid_0_MPORT_75_en = reset;
  assign valid_0_MPORT_79_data = 1'h0;
  assign valid_0_MPORT_79_addr = 4'h1;
  assign valid_0_MPORT_79_mask = 1'h1;
  assign valid_0_MPORT_79_en = reset;
  assign valid_0_MPORT_83_data = 1'h0;
  assign valid_0_MPORT_83_addr = 4'h2;
  assign valid_0_MPORT_83_mask = 1'h1;
  assign valid_0_MPORT_83_en = reset;
  assign valid_0_MPORT_87_data = 1'h0;
  assign valid_0_MPORT_87_addr = 4'h3;
  assign valid_0_MPORT_87_mask = 1'h1;
  assign valid_0_MPORT_87_en = reset;
  assign valid_0_MPORT_91_data = 1'h0;
  assign valid_0_MPORT_91_addr = 4'h4;
  assign valid_0_MPORT_91_mask = 1'h1;
  assign valid_0_MPORT_91_en = reset;
  assign valid_0_MPORT_95_data = 1'h0;
  assign valid_0_MPORT_95_addr = 4'h5;
  assign valid_0_MPORT_95_mask = 1'h1;
  assign valid_0_MPORT_95_en = reset;
  assign valid_0_MPORT_99_data = 1'h0;
  assign valid_0_MPORT_99_addr = 4'h6;
  assign valid_0_MPORT_99_mask = 1'h1;
  assign valid_0_MPORT_99_en = reset;
  assign valid_0_MPORT_103_data = 1'h0;
  assign valid_0_MPORT_103_addr = 4'h7;
  assign valid_0_MPORT_103_mask = 1'h1;
  assign valid_0_MPORT_103_en = reset;
  assign valid_0_MPORT_107_data = 1'h0;
  assign valid_0_MPORT_107_addr = 4'h8;
  assign valid_0_MPORT_107_mask = 1'h1;
  assign valid_0_MPORT_107_en = reset;
  assign valid_0_MPORT_111_data = 1'h0;
  assign valid_0_MPORT_111_addr = 4'h9;
  assign valid_0_MPORT_111_mask = 1'h1;
  assign valid_0_MPORT_111_en = reset;
  assign valid_0_MPORT_115_data = 1'h0;
  assign valid_0_MPORT_115_addr = 4'ha;
  assign valid_0_MPORT_115_mask = 1'h1;
  assign valid_0_MPORT_115_en = reset;
  assign valid_0_MPORT_119_data = 1'h0;
  assign valid_0_MPORT_119_addr = 4'hb;
  assign valid_0_MPORT_119_mask = 1'h1;
  assign valid_0_MPORT_119_en = reset;
  assign valid_0_MPORT_123_data = 1'h0;
  assign valid_0_MPORT_123_addr = 4'hc;
  assign valid_0_MPORT_123_mask = 1'h1;
  assign valid_0_MPORT_123_en = reset;
  assign valid_0_MPORT_127_data = 1'h0;
  assign valid_0_MPORT_127_addr = 4'hd;
  assign valid_0_MPORT_127_mask = 1'h1;
  assign valid_0_MPORT_127_en = reset;
  assign valid_0_MPORT_131_data = 1'h0;
  assign valid_0_MPORT_131_addr = 4'he;
  assign valid_0_MPORT_131_mask = 1'h1;
  assign valid_0_MPORT_131_en = reset;
  assign valid_0_MPORT_135_data = 1'h0;
  assign valid_0_MPORT_135_addr = 4'hf;
  assign valid_0_MPORT_135_mask = 1'h1;
  assign valid_0_MPORT_135_en = reset;
//   assign valid_1_MPORT_7_en = 1'h1;
  assign valid_1_MPORT_7_addr = io_raddr_0;
  assign valid_1_MPORT_7_data = valid_1[valid_1_MPORT_7_addr]; // @[BranchTargetBuffer.scala 102:20]
//   assign valid_1_MPORT_23_en = 1'h1;
  assign valid_1_MPORT_23_addr = io_raddr_1;
  assign valid_1_MPORT_23_data = valid_1[valid_1_MPORT_23_addr]; // @[BranchTargetBuffer.scala 102:20]
//   assign valid_1_MPORT_37_en = 1'h1;
  assign valid_1_MPORT_37_addr = io_waddr;
  assign valid_1_MPORT_37_data = valid_1[valid_1_MPORT_37_addr]; // @[BranchTargetBuffer.scala 102:20]
  assign valid_1_MPORT_63_data = 1'h1;
  assign valid_1_MPORT_63_addr = REG_73;
  assign valid_1_MPORT_63_mask = 1'h1;
  assign valid_1_MPORT_63_en = REG_30 & _GEN_2721;
  assign valid_1_MPORT_139_data = 1'h0;
  assign valid_1_MPORT_139_addr = 4'h0;
  assign valid_1_MPORT_139_mask = 1'h1;
  assign valid_1_MPORT_139_en = reset;
  assign valid_1_MPORT_143_data = 1'h0;
  assign valid_1_MPORT_143_addr = 4'h1;
  assign valid_1_MPORT_143_mask = 1'h1;
  assign valid_1_MPORT_143_en = reset;
  assign valid_1_MPORT_147_data = 1'h0;
  assign valid_1_MPORT_147_addr = 4'h2;
  assign valid_1_MPORT_147_mask = 1'h1;
  assign valid_1_MPORT_147_en = reset;
  assign valid_1_MPORT_151_data = 1'h0;
  assign valid_1_MPORT_151_addr = 4'h3;
  assign valid_1_MPORT_151_mask = 1'h1;
  assign valid_1_MPORT_151_en = reset;
  assign valid_1_MPORT_155_data = 1'h0;
  assign valid_1_MPORT_155_addr = 4'h4;
  assign valid_1_MPORT_155_mask = 1'h1;
  assign valid_1_MPORT_155_en = reset;
  assign valid_1_MPORT_159_data = 1'h0;
  assign valid_1_MPORT_159_addr = 4'h5;
  assign valid_1_MPORT_159_mask = 1'h1;
  assign valid_1_MPORT_159_en = reset;
  assign valid_1_MPORT_163_data = 1'h0;
  assign valid_1_MPORT_163_addr = 4'h6;
  assign valid_1_MPORT_163_mask = 1'h1;
  assign valid_1_MPORT_163_en = reset;
  assign valid_1_MPORT_167_data = 1'h0;
  assign valid_1_MPORT_167_addr = 4'h7;
  assign valid_1_MPORT_167_mask = 1'h1;
  assign valid_1_MPORT_167_en = reset;
  assign valid_1_MPORT_171_data = 1'h0;
  assign valid_1_MPORT_171_addr = 4'h8;
  assign valid_1_MPORT_171_mask = 1'h1;
  assign valid_1_MPORT_171_en = reset;
  assign valid_1_MPORT_175_data = 1'h0;
  assign valid_1_MPORT_175_addr = 4'h9;
  assign valid_1_MPORT_175_mask = 1'h1;
  assign valid_1_MPORT_175_en = reset;
  assign valid_1_MPORT_179_data = 1'h0;
  assign valid_1_MPORT_179_addr = 4'ha;
  assign valid_1_MPORT_179_mask = 1'h1;
  assign valid_1_MPORT_179_en = reset;
  assign valid_1_MPORT_183_data = 1'h0;
  assign valid_1_MPORT_183_addr = 4'hb;
  assign valid_1_MPORT_183_mask = 1'h1;
  assign valid_1_MPORT_183_en = reset;
  assign valid_1_MPORT_187_data = 1'h0;
  assign valid_1_MPORT_187_addr = 4'hc;
  assign valid_1_MPORT_187_mask = 1'h1;
  assign valid_1_MPORT_187_en = reset;
  assign valid_1_MPORT_191_data = 1'h0;
  assign valid_1_MPORT_191_addr = 4'hd;
  assign valid_1_MPORT_191_mask = 1'h1;
  assign valid_1_MPORT_191_en = reset;
  assign valid_1_MPORT_195_data = 1'h0;
  assign valid_1_MPORT_195_addr = 4'he;
  assign valid_1_MPORT_195_mask = 1'h1;
  assign valid_1_MPORT_195_en = reset;
  assign valid_1_MPORT_199_data = 1'h0;
  assign valid_1_MPORT_199_addr = 4'hf;
  assign valid_1_MPORT_199_mask = 1'h1;
  assign valid_1_MPORT_199_en = reset;
//   assign valid_2_MPORT_11_en = 1'h1;
  assign valid_2_MPORT_11_addr = io_raddr_0;
  assign valid_2_MPORT_11_data = valid_2[valid_2_MPORT_11_addr]; // @[BranchTargetBuffer.scala 102:20]
//   assign valid_2_MPORT_27_en = 1'h1;
  assign valid_2_MPORT_27_addr = io_raddr_1;
  assign valid_2_MPORT_27_data = valid_2[valid_2_MPORT_27_addr]; // @[BranchTargetBuffer.scala 102:20]
//   assign valid_2_MPORT_40_en = 1'h1;
  assign valid_2_MPORT_40_addr = io_waddr;
  assign valid_2_MPORT_40_data = valid_2[valid_2_MPORT_40_addr]; // @[BranchTargetBuffer.scala 102:20]
  assign valid_2_MPORT_67_data = 1'h1;
  assign valid_2_MPORT_67_addr = REG_81;
  assign valid_2_MPORT_67_mask = 1'h1;
  assign valid_2_MPORT_67_en = REG_30 & _GEN_2731;
  assign valid_2_MPORT_203_data = 1'h0;
  assign valid_2_MPORT_203_addr = 4'h0;
  assign valid_2_MPORT_203_mask = 1'h1;
  assign valid_2_MPORT_203_en = reset;
  assign valid_2_MPORT_207_data = 1'h0;
  assign valid_2_MPORT_207_addr = 4'h1;
  assign valid_2_MPORT_207_mask = 1'h1;
  assign valid_2_MPORT_207_en = reset;
  assign valid_2_MPORT_211_data = 1'h0;
  assign valid_2_MPORT_211_addr = 4'h2;
  assign valid_2_MPORT_211_mask = 1'h1;
  assign valid_2_MPORT_211_en = reset;
  assign valid_2_MPORT_215_data = 1'h0;
  assign valid_2_MPORT_215_addr = 4'h3;
  assign valid_2_MPORT_215_mask = 1'h1;
  assign valid_2_MPORT_215_en = reset;
  assign valid_2_MPORT_219_data = 1'h0;
  assign valid_2_MPORT_219_addr = 4'h4;
  assign valid_2_MPORT_219_mask = 1'h1;
  assign valid_2_MPORT_219_en = reset;
  assign valid_2_MPORT_223_data = 1'h0;
  assign valid_2_MPORT_223_addr = 4'h5;
  assign valid_2_MPORT_223_mask = 1'h1;
  assign valid_2_MPORT_223_en = reset;
  assign valid_2_MPORT_227_data = 1'h0;
  assign valid_2_MPORT_227_addr = 4'h6;
  assign valid_2_MPORT_227_mask = 1'h1;
  assign valid_2_MPORT_227_en = reset;
  assign valid_2_MPORT_231_data = 1'h0;
  assign valid_2_MPORT_231_addr = 4'h7;
  assign valid_2_MPORT_231_mask = 1'h1;
  assign valid_2_MPORT_231_en = reset;
  assign valid_2_MPORT_235_data = 1'h0;
  assign valid_2_MPORT_235_addr = 4'h8;
  assign valid_2_MPORT_235_mask = 1'h1;
  assign valid_2_MPORT_235_en = reset;
  assign valid_2_MPORT_239_data = 1'h0;
  assign valid_2_MPORT_239_addr = 4'h9;
  assign valid_2_MPORT_239_mask = 1'h1;
  assign valid_2_MPORT_239_en = reset;
  assign valid_2_MPORT_243_data = 1'h0;
  assign valid_2_MPORT_243_addr = 4'ha;
  assign valid_2_MPORT_243_mask = 1'h1;
  assign valid_2_MPORT_243_en = reset;
  assign valid_2_MPORT_247_data = 1'h0;
  assign valid_2_MPORT_247_addr = 4'hb;
  assign valid_2_MPORT_247_mask = 1'h1;
  assign valid_2_MPORT_247_en = reset;
  assign valid_2_MPORT_251_data = 1'h0;
  assign valid_2_MPORT_251_addr = 4'hc;
  assign valid_2_MPORT_251_mask = 1'h1;
  assign valid_2_MPORT_251_en = reset;
  assign valid_2_MPORT_255_data = 1'h0;
  assign valid_2_MPORT_255_addr = 4'hd;
  assign valid_2_MPORT_255_mask = 1'h1;
  assign valid_2_MPORT_255_en = reset;
  assign valid_2_MPORT_259_data = 1'h0;
  assign valid_2_MPORT_259_addr = 4'he;
  assign valid_2_MPORT_259_mask = 1'h1;
  assign valid_2_MPORT_259_en = reset;
  assign valid_2_MPORT_263_data = 1'h0;
  assign valid_2_MPORT_263_addr = 4'hf;
  assign valid_2_MPORT_263_mask = 1'h1;
  assign valid_2_MPORT_263_en = reset;
//   assign valid_3_MPORT_15_en = 1'h1;
  assign valid_3_MPORT_15_addr = io_raddr_0;
  assign valid_3_MPORT_15_data = valid_3[valid_3_MPORT_15_addr]; // @[BranchTargetBuffer.scala 102:20]
//   assign valid_3_MPORT_31_en = 1'h1;
  assign valid_3_MPORT_31_addr = io_raddr_1;
  assign valid_3_MPORT_31_data = valid_3[valid_3_MPORT_31_addr]; // @[BranchTargetBuffer.scala 102:20]
//   assign valid_3_MPORT_43_en = 1'h1;
  assign valid_3_MPORT_43_addr = io_waddr;
  assign valid_3_MPORT_43_data = valid_3[valid_3_MPORT_43_addr]; // @[BranchTargetBuffer.scala 102:20]
  assign valid_3_MPORT_71_data = 1'h1;
  assign valid_3_MPORT_71_addr = REG_89;
  assign valid_3_MPORT_71_mask = 1'h1;
  assign valid_3_MPORT_71_en = REG_30 & _GEN_2741;
  assign valid_3_MPORT_267_data = 1'h0;
  assign valid_3_MPORT_267_addr = 4'h0;
  assign valid_3_MPORT_267_mask = 1'h1;
  assign valid_3_MPORT_267_en = reset;
  assign valid_3_MPORT_271_data = 1'h0;
  assign valid_3_MPORT_271_addr = 4'h1;
  assign valid_3_MPORT_271_mask = 1'h1;
  assign valid_3_MPORT_271_en = reset;
  assign valid_3_MPORT_275_data = 1'h0;
  assign valid_3_MPORT_275_addr = 4'h2;
  assign valid_3_MPORT_275_mask = 1'h1;
  assign valid_3_MPORT_275_en = reset;
  assign valid_3_MPORT_279_data = 1'h0;
  assign valid_3_MPORT_279_addr = 4'h3;
  assign valid_3_MPORT_279_mask = 1'h1;
  assign valid_3_MPORT_279_en = reset;
  assign valid_3_MPORT_283_data = 1'h0;
  assign valid_3_MPORT_283_addr = 4'h4;
  assign valid_3_MPORT_283_mask = 1'h1;
  assign valid_3_MPORT_283_en = reset;
  assign valid_3_MPORT_287_data = 1'h0;
  assign valid_3_MPORT_287_addr = 4'h5;
  assign valid_3_MPORT_287_mask = 1'h1;
  assign valid_3_MPORT_287_en = reset;
  assign valid_3_MPORT_291_data = 1'h0;
  assign valid_3_MPORT_291_addr = 4'h6;
  assign valid_3_MPORT_291_mask = 1'h1;
  assign valid_3_MPORT_291_en = reset;
  assign valid_3_MPORT_295_data = 1'h0;
  assign valid_3_MPORT_295_addr = 4'h7;
  assign valid_3_MPORT_295_mask = 1'h1;
  assign valid_3_MPORT_295_en = reset;
  assign valid_3_MPORT_299_data = 1'h0;
  assign valid_3_MPORT_299_addr = 4'h8;
  assign valid_3_MPORT_299_mask = 1'h1;
  assign valid_3_MPORT_299_en = reset;
  assign valid_3_MPORT_303_data = 1'h0;
  assign valid_3_MPORT_303_addr = 4'h9;
  assign valid_3_MPORT_303_mask = 1'h1;
  assign valid_3_MPORT_303_en = reset;
  assign valid_3_MPORT_307_data = 1'h0;
  assign valid_3_MPORT_307_addr = 4'ha;
  assign valid_3_MPORT_307_mask = 1'h1;
  assign valid_3_MPORT_307_en = reset;
  assign valid_3_MPORT_311_data = 1'h0;
  assign valid_3_MPORT_311_addr = 4'hb;
  assign valid_3_MPORT_311_mask = 1'h1;
  assign valid_3_MPORT_311_en = reset;
  assign valid_3_MPORT_315_data = 1'h0;
  assign valid_3_MPORT_315_addr = 4'hc;
  assign valid_3_MPORT_315_mask = 1'h1;
  assign valid_3_MPORT_315_en = reset;
  assign valid_3_MPORT_319_data = 1'h0;
  assign valid_3_MPORT_319_addr = 4'hd;
  assign valid_3_MPORT_319_mask = 1'h1;
  assign valid_3_MPORT_319_en = reset;
  assign valid_3_MPORT_323_data = 1'h0;
  assign valid_3_MPORT_323_addr = 4'he;
  assign valid_3_MPORT_323_mask = 1'h1;
  assign valid_3_MPORT_323_en = reset;
  assign valid_3_MPORT_327_data = 1'h0;
  assign valid_3_MPORT_327_addr = 4'hf;
  assign valid_3_MPORT_327_mask = 1'h1;
  assign valid_3_MPORT_327_en = reset;
  assign io_rhit_0 = REG__3 & _WIRE_8_3_tag == REG_10 | (REG__2 & _WIRE_8_2_tag == REG_7 | (REG__1 & _WIRE_8_1_tag ==
    REG_4 | REG__0 & _WIRE_8_0_tag == REG_1)); // @[BranchTargetBuffer.scala 133:66 134:20]
  assign io_rhit_1 = REG_13_3 & _WIRE_27_3_tag == REG_23 | (REG_13_2 & _WIRE_27_2_tag == REG_20 | (REG_13_1 &
    _WIRE_27_1_tag == REG_17 | REG_13_0 & _WIRE_27_0_tag == REG_14)); // @[BranchTargetBuffer.scala 133:66 134:20]
  assign io_rtarget_0 = REG__3 & _WIRE_8_3_tag == REG_10 ? _WIRE_8_3_target : _GEN_499; // @[BranchTargetBuffer.scala 133:66 135:23]
  assign io_rtarget_1 = REG_13_3 & _WIRE_27_3_tag == REG_23 ? _WIRE_27_3_target : _GEN_1228; // @[BranchTargetBuffer.scala 133:66 135:23]
  always @(posedge clock) begin
    if (btb_tag_0_MPORT_44_en & btb_tag_0_MPORT_44_mask) begin
      btb_tag_0[btb_tag_0_MPORT_44_addr] <= btb_tag_0_MPORT_44_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_56_en & btb_tag_0_MPORT_56_mask) begin
      btb_tag_0[btb_tag_0_MPORT_56_addr] <= btb_tag_0_MPORT_56_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_72_en & btb_tag_0_MPORT_72_mask) begin
      btb_tag_0[btb_tag_0_MPORT_72_addr] <= btb_tag_0_MPORT_72_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_76_en & btb_tag_0_MPORT_76_mask) begin
      btb_tag_0[btb_tag_0_MPORT_76_addr] <= btb_tag_0_MPORT_76_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_80_en & btb_tag_0_MPORT_80_mask) begin
      btb_tag_0[btb_tag_0_MPORT_80_addr] <= btb_tag_0_MPORT_80_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_84_en & btb_tag_0_MPORT_84_mask) begin
      btb_tag_0[btb_tag_0_MPORT_84_addr] <= btb_tag_0_MPORT_84_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_88_en & btb_tag_0_MPORT_88_mask) begin
      btb_tag_0[btb_tag_0_MPORT_88_addr] <= btb_tag_0_MPORT_88_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_92_en & btb_tag_0_MPORT_92_mask) begin
      btb_tag_0[btb_tag_0_MPORT_92_addr] <= btb_tag_0_MPORT_92_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_96_en & btb_tag_0_MPORT_96_mask) begin
      btb_tag_0[btb_tag_0_MPORT_96_addr] <= btb_tag_0_MPORT_96_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_100_en & btb_tag_0_MPORT_100_mask) begin
      btb_tag_0[btb_tag_0_MPORT_100_addr] <= btb_tag_0_MPORT_100_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_104_en & btb_tag_0_MPORT_104_mask) begin
      btb_tag_0[btb_tag_0_MPORT_104_addr] <= btb_tag_0_MPORT_104_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_108_en & btb_tag_0_MPORT_108_mask) begin
      btb_tag_0[btb_tag_0_MPORT_108_addr] <= btb_tag_0_MPORT_108_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_112_en & btb_tag_0_MPORT_112_mask) begin
      btb_tag_0[btb_tag_0_MPORT_112_addr] <= btb_tag_0_MPORT_112_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_116_en & btb_tag_0_MPORT_116_mask) begin
      btb_tag_0[btb_tag_0_MPORT_116_addr] <= btb_tag_0_MPORT_116_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_120_en & btb_tag_0_MPORT_120_mask) begin
      btb_tag_0[btb_tag_0_MPORT_120_addr] <= btb_tag_0_MPORT_120_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_124_en & btb_tag_0_MPORT_124_mask) begin
      btb_tag_0[btb_tag_0_MPORT_124_addr] <= btb_tag_0_MPORT_124_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_128_en & btb_tag_0_MPORT_128_mask) begin
      btb_tag_0[btb_tag_0_MPORT_128_addr] <= btb_tag_0_MPORT_128_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_0_MPORT_132_en & btb_tag_0_MPORT_132_mask) begin
      btb_tag_0[btb_tag_0_MPORT_132_addr] <= btb_tag_0_MPORT_132_data; // @[BranchTargetBuffer.scala 90:30]
    end
//     btb_tag_0_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_tag_0_MPORT_addr_pipe_0 <= io_raddr_0;
    end
//     btb_tag_0_MPORT_16_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_tag_0_MPORT_16_addr_pipe_0 <= io_raddr_1;
    end
//     btb_tag_0_MPORT_32_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_tag_0_MPORT_32_addr_pipe_0 <= io_waddr;
    end
    if (btb_tag_1_MPORT_47_en & btb_tag_1_MPORT_47_mask) begin
      btb_tag_1[btb_tag_1_MPORT_47_addr] <= btb_tag_1_MPORT_47_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_60_en & btb_tag_1_MPORT_60_mask) begin
      btb_tag_1[btb_tag_1_MPORT_60_addr] <= btb_tag_1_MPORT_60_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_136_en & btb_tag_1_MPORT_136_mask) begin
      btb_tag_1[btb_tag_1_MPORT_136_addr] <= btb_tag_1_MPORT_136_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_140_en & btb_tag_1_MPORT_140_mask) begin
      btb_tag_1[btb_tag_1_MPORT_140_addr] <= btb_tag_1_MPORT_140_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_144_en & btb_tag_1_MPORT_144_mask) begin
      btb_tag_1[btb_tag_1_MPORT_144_addr] <= btb_tag_1_MPORT_144_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_148_en & btb_tag_1_MPORT_148_mask) begin
      btb_tag_1[btb_tag_1_MPORT_148_addr] <= btb_tag_1_MPORT_148_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_152_en & btb_tag_1_MPORT_152_mask) begin
      btb_tag_1[btb_tag_1_MPORT_152_addr] <= btb_tag_1_MPORT_152_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_156_en & btb_tag_1_MPORT_156_mask) begin
      btb_tag_1[btb_tag_1_MPORT_156_addr] <= btb_tag_1_MPORT_156_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_160_en & btb_tag_1_MPORT_160_mask) begin
      btb_tag_1[btb_tag_1_MPORT_160_addr] <= btb_tag_1_MPORT_160_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_164_en & btb_tag_1_MPORT_164_mask) begin
      btb_tag_1[btb_tag_1_MPORT_164_addr] <= btb_tag_1_MPORT_164_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_168_en & btb_tag_1_MPORT_168_mask) begin
      btb_tag_1[btb_tag_1_MPORT_168_addr] <= btb_tag_1_MPORT_168_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_172_en & btb_tag_1_MPORT_172_mask) begin
      btb_tag_1[btb_tag_1_MPORT_172_addr] <= btb_tag_1_MPORT_172_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_176_en & btb_tag_1_MPORT_176_mask) begin
      btb_tag_1[btb_tag_1_MPORT_176_addr] <= btb_tag_1_MPORT_176_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_180_en & btb_tag_1_MPORT_180_mask) begin
      btb_tag_1[btb_tag_1_MPORT_180_addr] <= btb_tag_1_MPORT_180_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_184_en & btb_tag_1_MPORT_184_mask) begin
      btb_tag_1[btb_tag_1_MPORT_184_addr] <= btb_tag_1_MPORT_184_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_188_en & btb_tag_1_MPORT_188_mask) begin
      btb_tag_1[btb_tag_1_MPORT_188_addr] <= btb_tag_1_MPORT_188_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_192_en & btb_tag_1_MPORT_192_mask) begin
      btb_tag_1[btb_tag_1_MPORT_192_addr] <= btb_tag_1_MPORT_192_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_1_MPORT_196_en & btb_tag_1_MPORT_196_mask) begin
      btb_tag_1[btb_tag_1_MPORT_196_addr] <= btb_tag_1_MPORT_196_data; // @[BranchTargetBuffer.scala 90:30]
    end
//     btb_tag_1_MPORT_4_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_tag_1_MPORT_4_addr_pipe_0 <= io_raddr_0;
    end
//     btb_tag_1_MPORT_20_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_tag_1_MPORT_20_addr_pipe_0 <= io_raddr_1;
    end
//     btb_tag_1_MPORT_35_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_tag_1_MPORT_35_addr_pipe_0 <= io_waddr;
    end
    if (btb_tag_2_MPORT_50_en & btb_tag_2_MPORT_50_mask) begin
      btb_tag_2[btb_tag_2_MPORT_50_addr] <= btb_tag_2_MPORT_50_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_64_en & btb_tag_2_MPORT_64_mask) begin
      btb_tag_2[btb_tag_2_MPORT_64_addr] <= btb_tag_2_MPORT_64_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_200_en & btb_tag_2_MPORT_200_mask) begin
      btb_tag_2[btb_tag_2_MPORT_200_addr] <= btb_tag_2_MPORT_200_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_204_en & btb_tag_2_MPORT_204_mask) begin
      btb_tag_2[btb_tag_2_MPORT_204_addr] <= btb_tag_2_MPORT_204_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_208_en & btb_tag_2_MPORT_208_mask) begin
      btb_tag_2[btb_tag_2_MPORT_208_addr] <= btb_tag_2_MPORT_208_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_212_en & btb_tag_2_MPORT_212_mask) begin
      btb_tag_2[btb_tag_2_MPORT_212_addr] <= btb_tag_2_MPORT_212_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_216_en & btb_tag_2_MPORT_216_mask) begin
      btb_tag_2[btb_tag_2_MPORT_216_addr] <= btb_tag_2_MPORT_216_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_220_en & btb_tag_2_MPORT_220_mask) begin
      btb_tag_2[btb_tag_2_MPORT_220_addr] <= btb_tag_2_MPORT_220_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_224_en & btb_tag_2_MPORT_224_mask) begin
      btb_tag_2[btb_tag_2_MPORT_224_addr] <= btb_tag_2_MPORT_224_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_228_en & btb_tag_2_MPORT_228_mask) begin
      btb_tag_2[btb_tag_2_MPORT_228_addr] <= btb_tag_2_MPORT_228_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_232_en & btb_tag_2_MPORT_232_mask) begin
      btb_tag_2[btb_tag_2_MPORT_232_addr] <= btb_tag_2_MPORT_232_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_236_en & btb_tag_2_MPORT_236_mask) begin
      btb_tag_2[btb_tag_2_MPORT_236_addr] <= btb_tag_2_MPORT_236_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_240_en & btb_tag_2_MPORT_240_mask) begin
      btb_tag_2[btb_tag_2_MPORT_240_addr] <= btb_tag_2_MPORT_240_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_244_en & btb_tag_2_MPORT_244_mask) begin
      btb_tag_2[btb_tag_2_MPORT_244_addr] <= btb_tag_2_MPORT_244_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_248_en & btb_tag_2_MPORT_248_mask) begin
      btb_tag_2[btb_tag_2_MPORT_248_addr] <= btb_tag_2_MPORT_248_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_252_en & btb_tag_2_MPORT_252_mask) begin
      btb_tag_2[btb_tag_2_MPORT_252_addr] <= btb_tag_2_MPORT_252_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_256_en & btb_tag_2_MPORT_256_mask) begin
      btb_tag_2[btb_tag_2_MPORT_256_addr] <= btb_tag_2_MPORT_256_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_2_MPORT_260_en & btb_tag_2_MPORT_260_mask) begin
      btb_tag_2[btb_tag_2_MPORT_260_addr] <= btb_tag_2_MPORT_260_data; // @[BranchTargetBuffer.scala 90:30]
    end
//     btb_tag_2_MPORT_8_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_tag_2_MPORT_8_addr_pipe_0 <= io_raddr_0;
    end
//     btb_tag_2_MPORT_24_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_tag_2_MPORT_24_addr_pipe_0 <= io_raddr_1;
    end
//     btb_tag_2_MPORT_38_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_tag_2_MPORT_38_addr_pipe_0 <= io_waddr;
    end
    if (btb_tag_3_MPORT_53_en & btb_tag_3_MPORT_53_mask) begin
      btb_tag_3[btb_tag_3_MPORT_53_addr] <= btb_tag_3_MPORT_53_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_68_en & btb_tag_3_MPORT_68_mask) begin
      btb_tag_3[btb_tag_3_MPORT_68_addr] <= btb_tag_3_MPORT_68_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_264_en & btb_tag_3_MPORT_264_mask) begin
      btb_tag_3[btb_tag_3_MPORT_264_addr] <= btb_tag_3_MPORT_264_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_268_en & btb_tag_3_MPORT_268_mask) begin
      btb_tag_3[btb_tag_3_MPORT_268_addr] <= btb_tag_3_MPORT_268_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_272_en & btb_tag_3_MPORT_272_mask) begin
      btb_tag_3[btb_tag_3_MPORT_272_addr] <= btb_tag_3_MPORT_272_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_276_en & btb_tag_3_MPORT_276_mask) begin
      btb_tag_3[btb_tag_3_MPORT_276_addr] <= btb_tag_3_MPORT_276_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_280_en & btb_tag_3_MPORT_280_mask) begin
      btb_tag_3[btb_tag_3_MPORT_280_addr] <= btb_tag_3_MPORT_280_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_284_en & btb_tag_3_MPORT_284_mask) begin
      btb_tag_3[btb_tag_3_MPORT_284_addr] <= btb_tag_3_MPORT_284_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_288_en & btb_tag_3_MPORT_288_mask) begin
      btb_tag_3[btb_tag_3_MPORT_288_addr] <= btb_tag_3_MPORT_288_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_292_en & btb_tag_3_MPORT_292_mask) begin
      btb_tag_3[btb_tag_3_MPORT_292_addr] <= btb_tag_3_MPORT_292_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_296_en & btb_tag_3_MPORT_296_mask) begin
      btb_tag_3[btb_tag_3_MPORT_296_addr] <= btb_tag_3_MPORT_296_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_300_en & btb_tag_3_MPORT_300_mask) begin
      btb_tag_3[btb_tag_3_MPORT_300_addr] <= btb_tag_3_MPORT_300_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_304_en & btb_tag_3_MPORT_304_mask) begin
      btb_tag_3[btb_tag_3_MPORT_304_addr] <= btb_tag_3_MPORT_304_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_308_en & btb_tag_3_MPORT_308_mask) begin
      btb_tag_3[btb_tag_3_MPORT_308_addr] <= btb_tag_3_MPORT_308_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_312_en & btb_tag_3_MPORT_312_mask) begin
      btb_tag_3[btb_tag_3_MPORT_312_addr] <= btb_tag_3_MPORT_312_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_316_en & btb_tag_3_MPORT_316_mask) begin
      btb_tag_3[btb_tag_3_MPORT_316_addr] <= btb_tag_3_MPORT_316_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_320_en & btb_tag_3_MPORT_320_mask) begin
      btb_tag_3[btb_tag_3_MPORT_320_addr] <= btb_tag_3_MPORT_320_data; // @[BranchTargetBuffer.scala 90:30]
    end
    if (btb_tag_3_MPORT_324_en & btb_tag_3_MPORT_324_mask) begin
      btb_tag_3[btb_tag_3_MPORT_324_addr] <= btb_tag_3_MPORT_324_data; // @[BranchTargetBuffer.scala 90:30]
    end
//     btb_tag_3_MPORT_12_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_tag_3_MPORT_12_addr_pipe_0 <= io_raddr_0;
    end
//     btb_tag_3_MPORT_28_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_tag_3_MPORT_28_addr_pipe_0 <= io_raddr_1;
    end
//     btb_tag_3_MPORT_41_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_tag_3_MPORT_41_addr_pipe_0 <= io_waddr;
    end
    if (btb_target_0_MPORT_45_en & btb_target_0_MPORT_45_mask) begin
      btb_target_0[btb_target_0_MPORT_45_addr] <= btb_target_0_MPORT_45_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_57_en & btb_target_0_MPORT_57_mask) begin
      btb_target_0[btb_target_0_MPORT_57_addr] <= btb_target_0_MPORT_57_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_73_en & btb_target_0_MPORT_73_mask) begin
      btb_target_0[btb_target_0_MPORT_73_addr] <= btb_target_0_MPORT_73_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_77_en & btb_target_0_MPORT_77_mask) begin
      btb_target_0[btb_target_0_MPORT_77_addr] <= btb_target_0_MPORT_77_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_81_en & btb_target_0_MPORT_81_mask) begin
      btb_target_0[btb_target_0_MPORT_81_addr] <= btb_target_0_MPORT_81_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_85_en & btb_target_0_MPORT_85_mask) begin
      btb_target_0[btb_target_0_MPORT_85_addr] <= btb_target_0_MPORT_85_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_89_en & btb_target_0_MPORT_89_mask) begin
      btb_target_0[btb_target_0_MPORT_89_addr] <= btb_target_0_MPORT_89_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_93_en & btb_target_0_MPORT_93_mask) begin
      btb_target_0[btb_target_0_MPORT_93_addr] <= btb_target_0_MPORT_93_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_97_en & btb_target_0_MPORT_97_mask) begin
      btb_target_0[btb_target_0_MPORT_97_addr] <= btb_target_0_MPORT_97_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_101_en & btb_target_0_MPORT_101_mask) begin
      btb_target_0[btb_target_0_MPORT_101_addr] <= btb_target_0_MPORT_101_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_105_en & btb_target_0_MPORT_105_mask) begin
      btb_target_0[btb_target_0_MPORT_105_addr] <= btb_target_0_MPORT_105_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_109_en & btb_target_0_MPORT_109_mask) begin
      btb_target_0[btb_target_0_MPORT_109_addr] <= btb_target_0_MPORT_109_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_113_en & btb_target_0_MPORT_113_mask) begin
      btb_target_0[btb_target_0_MPORT_113_addr] <= btb_target_0_MPORT_113_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_117_en & btb_target_0_MPORT_117_mask) begin
      btb_target_0[btb_target_0_MPORT_117_addr] <= btb_target_0_MPORT_117_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_121_en & btb_target_0_MPORT_121_mask) begin
      btb_target_0[btb_target_0_MPORT_121_addr] <= btb_target_0_MPORT_121_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_125_en & btb_target_0_MPORT_125_mask) begin
      btb_target_0[btb_target_0_MPORT_125_addr] <= btb_target_0_MPORT_125_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_129_en & btb_target_0_MPORT_129_mask) begin
      btb_target_0[btb_target_0_MPORT_129_addr] <= btb_target_0_MPORT_129_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_0_MPORT_133_en & btb_target_0_MPORT_133_mask) begin
      btb_target_0[btb_target_0_MPORT_133_addr] <= btb_target_0_MPORT_133_data; // @[BranchTargetBuffer.scala 94:33]
    end
//     btb_target_0_MPORT_1_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_target_0_MPORT_1_addr_pipe_0 <= io_raddr_0;
    end
//     btb_target_0_MPORT_17_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_target_0_MPORT_17_addr_pipe_0 <= io_raddr_1;
    end
    if (btb_target_1_MPORT_48_en & btb_target_1_MPORT_48_mask) begin
      btb_target_1[btb_target_1_MPORT_48_addr] <= btb_target_1_MPORT_48_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_61_en & btb_target_1_MPORT_61_mask) begin
      btb_target_1[btb_target_1_MPORT_61_addr] <= btb_target_1_MPORT_61_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_137_en & btb_target_1_MPORT_137_mask) begin
      btb_target_1[btb_target_1_MPORT_137_addr] <= btb_target_1_MPORT_137_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_141_en & btb_target_1_MPORT_141_mask) begin
      btb_target_1[btb_target_1_MPORT_141_addr] <= btb_target_1_MPORT_141_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_145_en & btb_target_1_MPORT_145_mask) begin
      btb_target_1[btb_target_1_MPORT_145_addr] <= btb_target_1_MPORT_145_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_149_en & btb_target_1_MPORT_149_mask) begin
      btb_target_1[btb_target_1_MPORT_149_addr] <= btb_target_1_MPORT_149_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_153_en & btb_target_1_MPORT_153_mask) begin
      btb_target_1[btb_target_1_MPORT_153_addr] <= btb_target_1_MPORT_153_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_157_en & btb_target_1_MPORT_157_mask) begin
      btb_target_1[btb_target_1_MPORT_157_addr] <= btb_target_1_MPORT_157_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_161_en & btb_target_1_MPORT_161_mask) begin
      btb_target_1[btb_target_1_MPORT_161_addr] <= btb_target_1_MPORT_161_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_165_en & btb_target_1_MPORT_165_mask) begin
      btb_target_1[btb_target_1_MPORT_165_addr] <= btb_target_1_MPORT_165_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_169_en & btb_target_1_MPORT_169_mask) begin
      btb_target_1[btb_target_1_MPORT_169_addr] <= btb_target_1_MPORT_169_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_173_en & btb_target_1_MPORT_173_mask) begin
      btb_target_1[btb_target_1_MPORT_173_addr] <= btb_target_1_MPORT_173_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_177_en & btb_target_1_MPORT_177_mask) begin
      btb_target_1[btb_target_1_MPORT_177_addr] <= btb_target_1_MPORT_177_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_181_en & btb_target_1_MPORT_181_mask) begin
      btb_target_1[btb_target_1_MPORT_181_addr] <= btb_target_1_MPORT_181_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_185_en & btb_target_1_MPORT_185_mask) begin
      btb_target_1[btb_target_1_MPORT_185_addr] <= btb_target_1_MPORT_185_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_189_en & btb_target_1_MPORT_189_mask) begin
      btb_target_1[btb_target_1_MPORT_189_addr] <= btb_target_1_MPORT_189_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_193_en & btb_target_1_MPORT_193_mask) begin
      btb_target_1[btb_target_1_MPORT_193_addr] <= btb_target_1_MPORT_193_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_1_MPORT_197_en & btb_target_1_MPORT_197_mask) begin
      btb_target_1[btb_target_1_MPORT_197_addr] <= btb_target_1_MPORT_197_data; // @[BranchTargetBuffer.scala 94:33]
    end
//     btb_target_1_MPORT_5_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_target_1_MPORT_5_addr_pipe_0 <= io_raddr_0;
    end
//     btb_target_1_MPORT_21_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_target_1_MPORT_21_addr_pipe_0 <= io_raddr_1;
    end
    if (btb_target_2_MPORT_51_en & btb_target_2_MPORT_51_mask) begin
      btb_target_2[btb_target_2_MPORT_51_addr] <= btb_target_2_MPORT_51_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_65_en & btb_target_2_MPORT_65_mask) begin
      btb_target_2[btb_target_2_MPORT_65_addr] <= btb_target_2_MPORT_65_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_201_en & btb_target_2_MPORT_201_mask) begin
      btb_target_2[btb_target_2_MPORT_201_addr] <= btb_target_2_MPORT_201_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_205_en & btb_target_2_MPORT_205_mask) begin
      btb_target_2[btb_target_2_MPORT_205_addr] <= btb_target_2_MPORT_205_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_209_en & btb_target_2_MPORT_209_mask) begin
      btb_target_2[btb_target_2_MPORT_209_addr] <= btb_target_2_MPORT_209_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_213_en & btb_target_2_MPORT_213_mask) begin
      btb_target_2[btb_target_2_MPORT_213_addr] <= btb_target_2_MPORT_213_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_217_en & btb_target_2_MPORT_217_mask) begin
      btb_target_2[btb_target_2_MPORT_217_addr] <= btb_target_2_MPORT_217_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_221_en & btb_target_2_MPORT_221_mask) begin
      btb_target_2[btb_target_2_MPORT_221_addr] <= btb_target_2_MPORT_221_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_225_en & btb_target_2_MPORT_225_mask) begin
      btb_target_2[btb_target_2_MPORT_225_addr] <= btb_target_2_MPORT_225_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_229_en & btb_target_2_MPORT_229_mask) begin
      btb_target_2[btb_target_2_MPORT_229_addr] <= btb_target_2_MPORT_229_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_233_en & btb_target_2_MPORT_233_mask) begin
      btb_target_2[btb_target_2_MPORT_233_addr] <= btb_target_2_MPORT_233_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_237_en & btb_target_2_MPORT_237_mask) begin
      btb_target_2[btb_target_2_MPORT_237_addr] <= btb_target_2_MPORT_237_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_241_en & btb_target_2_MPORT_241_mask) begin
      btb_target_2[btb_target_2_MPORT_241_addr] <= btb_target_2_MPORT_241_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_245_en & btb_target_2_MPORT_245_mask) begin
      btb_target_2[btb_target_2_MPORT_245_addr] <= btb_target_2_MPORT_245_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_249_en & btb_target_2_MPORT_249_mask) begin
      btb_target_2[btb_target_2_MPORT_249_addr] <= btb_target_2_MPORT_249_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_253_en & btb_target_2_MPORT_253_mask) begin
      btb_target_2[btb_target_2_MPORT_253_addr] <= btb_target_2_MPORT_253_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_257_en & btb_target_2_MPORT_257_mask) begin
      btb_target_2[btb_target_2_MPORT_257_addr] <= btb_target_2_MPORT_257_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_2_MPORT_261_en & btb_target_2_MPORT_261_mask) begin
      btb_target_2[btb_target_2_MPORT_261_addr] <= btb_target_2_MPORT_261_data; // @[BranchTargetBuffer.scala 94:33]
    end
//     btb_target_2_MPORT_9_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_target_2_MPORT_9_addr_pipe_0 <= io_raddr_0;
    end
//     btb_target_2_MPORT_25_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_target_2_MPORT_25_addr_pipe_0 <= io_raddr_1;
    end
    if (btb_target_3_MPORT_54_en & btb_target_3_MPORT_54_mask) begin
      btb_target_3[btb_target_3_MPORT_54_addr] <= btb_target_3_MPORT_54_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_69_en & btb_target_3_MPORT_69_mask) begin
      btb_target_3[btb_target_3_MPORT_69_addr] <= btb_target_3_MPORT_69_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_265_en & btb_target_3_MPORT_265_mask) begin
      btb_target_3[btb_target_3_MPORT_265_addr] <= btb_target_3_MPORT_265_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_269_en & btb_target_3_MPORT_269_mask) begin
      btb_target_3[btb_target_3_MPORT_269_addr] <= btb_target_3_MPORT_269_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_273_en & btb_target_3_MPORT_273_mask) begin
      btb_target_3[btb_target_3_MPORT_273_addr] <= btb_target_3_MPORT_273_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_277_en & btb_target_3_MPORT_277_mask) begin
      btb_target_3[btb_target_3_MPORT_277_addr] <= btb_target_3_MPORT_277_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_281_en & btb_target_3_MPORT_281_mask) begin
      btb_target_3[btb_target_3_MPORT_281_addr] <= btb_target_3_MPORT_281_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_285_en & btb_target_3_MPORT_285_mask) begin
      btb_target_3[btb_target_3_MPORT_285_addr] <= btb_target_3_MPORT_285_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_289_en & btb_target_3_MPORT_289_mask) begin
      btb_target_3[btb_target_3_MPORT_289_addr] <= btb_target_3_MPORT_289_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_293_en & btb_target_3_MPORT_293_mask) begin
      btb_target_3[btb_target_3_MPORT_293_addr] <= btb_target_3_MPORT_293_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_297_en & btb_target_3_MPORT_297_mask) begin
      btb_target_3[btb_target_3_MPORT_297_addr] <= btb_target_3_MPORT_297_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_301_en & btb_target_3_MPORT_301_mask) begin
      btb_target_3[btb_target_3_MPORT_301_addr] <= btb_target_3_MPORT_301_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_305_en & btb_target_3_MPORT_305_mask) begin
      btb_target_3[btb_target_3_MPORT_305_addr] <= btb_target_3_MPORT_305_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_309_en & btb_target_3_MPORT_309_mask) begin
      btb_target_3[btb_target_3_MPORT_309_addr] <= btb_target_3_MPORT_309_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_313_en & btb_target_3_MPORT_313_mask) begin
      btb_target_3[btb_target_3_MPORT_313_addr] <= btb_target_3_MPORT_313_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_317_en & btb_target_3_MPORT_317_mask) begin
      btb_target_3[btb_target_3_MPORT_317_addr] <= btb_target_3_MPORT_317_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_321_en & btb_target_3_MPORT_321_mask) begin
      btb_target_3[btb_target_3_MPORT_321_addr] <= btb_target_3_MPORT_321_data; // @[BranchTargetBuffer.scala 94:33]
    end
    if (btb_target_3_MPORT_325_en & btb_target_3_MPORT_325_mask) begin
      btb_target_3[btb_target_3_MPORT_325_addr] <= btb_target_3_MPORT_325_data; // @[BranchTargetBuffer.scala 94:33]
    end
//     btb_target_3_MPORT_13_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_target_3_MPORT_13_addr_pipe_0 <= io_raddr_0;
    end
//     btb_target_3_MPORT_29_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      btb_target_3_MPORT_29_addr_pipe_0 <= io_raddr_1;
    end
    if (valid_0_MPORT_59_en & valid_0_MPORT_59_mask) begin
      valid_0[valid_0_MPORT_59_addr] <= valid_0_MPORT_59_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_75_en & valid_0_MPORT_75_mask) begin
      valid_0[valid_0_MPORT_75_addr] <= valid_0_MPORT_75_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_79_en & valid_0_MPORT_79_mask) begin
      valid_0[valid_0_MPORT_79_addr] <= valid_0_MPORT_79_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_83_en & valid_0_MPORT_83_mask) begin
      valid_0[valid_0_MPORT_83_addr] <= valid_0_MPORT_83_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_87_en & valid_0_MPORT_87_mask) begin
      valid_0[valid_0_MPORT_87_addr] <= valid_0_MPORT_87_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_91_en & valid_0_MPORT_91_mask) begin
      valid_0[valid_0_MPORT_91_addr] <= valid_0_MPORT_91_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_95_en & valid_0_MPORT_95_mask) begin
      valid_0[valid_0_MPORT_95_addr] <= valid_0_MPORT_95_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_99_en & valid_0_MPORT_99_mask) begin
      valid_0[valid_0_MPORT_99_addr] <= valid_0_MPORT_99_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_103_en & valid_0_MPORT_103_mask) begin
      valid_0[valid_0_MPORT_103_addr] <= valid_0_MPORT_103_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_107_en & valid_0_MPORT_107_mask) begin
      valid_0[valid_0_MPORT_107_addr] <= valid_0_MPORT_107_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_111_en & valid_0_MPORT_111_mask) begin
      valid_0[valid_0_MPORT_111_addr] <= valid_0_MPORT_111_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_115_en & valid_0_MPORT_115_mask) begin
      valid_0[valid_0_MPORT_115_addr] <= valid_0_MPORT_115_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_119_en & valid_0_MPORT_119_mask) begin
      valid_0[valid_0_MPORT_119_addr] <= valid_0_MPORT_119_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_123_en & valid_0_MPORT_123_mask) begin
      valid_0[valid_0_MPORT_123_addr] <= valid_0_MPORT_123_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_127_en & valid_0_MPORT_127_mask) begin
      valid_0[valid_0_MPORT_127_addr] <= valid_0_MPORT_127_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_131_en & valid_0_MPORT_131_mask) begin
      valid_0[valid_0_MPORT_131_addr] <= valid_0_MPORT_131_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_0_MPORT_135_en & valid_0_MPORT_135_mask) begin
      valid_0[valid_0_MPORT_135_addr] <= valid_0_MPORT_135_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_63_en & valid_1_MPORT_63_mask) begin
      valid_1[valid_1_MPORT_63_addr] <= valid_1_MPORT_63_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_139_en & valid_1_MPORT_139_mask) begin
      valid_1[valid_1_MPORT_139_addr] <= valid_1_MPORT_139_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_143_en & valid_1_MPORT_143_mask) begin
      valid_1[valid_1_MPORT_143_addr] <= valid_1_MPORT_143_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_147_en & valid_1_MPORT_147_mask) begin
      valid_1[valid_1_MPORT_147_addr] <= valid_1_MPORT_147_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_151_en & valid_1_MPORT_151_mask) begin
      valid_1[valid_1_MPORT_151_addr] <= valid_1_MPORT_151_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_155_en & valid_1_MPORT_155_mask) begin
      valid_1[valid_1_MPORT_155_addr] <= valid_1_MPORT_155_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_159_en & valid_1_MPORT_159_mask) begin
      valid_1[valid_1_MPORT_159_addr] <= valid_1_MPORT_159_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_163_en & valid_1_MPORT_163_mask) begin
      valid_1[valid_1_MPORT_163_addr] <= valid_1_MPORT_163_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_167_en & valid_1_MPORT_167_mask) begin
      valid_1[valid_1_MPORT_167_addr] <= valid_1_MPORT_167_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_171_en & valid_1_MPORT_171_mask) begin
      valid_1[valid_1_MPORT_171_addr] <= valid_1_MPORT_171_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_175_en & valid_1_MPORT_175_mask) begin
      valid_1[valid_1_MPORT_175_addr] <= valid_1_MPORT_175_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_179_en & valid_1_MPORT_179_mask) begin
      valid_1[valid_1_MPORT_179_addr] <= valid_1_MPORT_179_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_183_en & valid_1_MPORT_183_mask) begin
      valid_1[valid_1_MPORT_183_addr] <= valid_1_MPORT_183_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_187_en & valid_1_MPORT_187_mask) begin
      valid_1[valid_1_MPORT_187_addr] <= valid_1_MPORT_187_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_191_en & valid_1_MPORT_191_mask) begin
      valid_1[valid_1_MPORT_191_addr] <= valid_1_MPORT_191_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_195_en & valid_1_MPORT_195_mask) begin
      valid_1[valid_1_MPORT_195_addr] <= valid_1_MPORT_195_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_1_MPORT_199_en & valid_1_MPORT_199_mask) begin
      valid_1[valid_1_MPORT_199_addr] <= valid_1_MPORT_199_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_67_en & valid_2_MPORT_67_mask) begin
      valid_2[valid_2_MPORT_67_addr] <= valid_2_MPORT_67_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_203_en & valid_2_MPORT_203_mask) begin
      valid_2[valid_2_MPORT_203_addr] <= valid_2_MPORT_203_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_207_en & valid_2_MPORT_207_mask) begin
      valid_2[valid_2_MPORT_207_addr] <= valid_2_MPORT_207_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_211_en & valid_2_MPORT_211_mask) begin
      valid_2[valid_2_MPORT_211_addr] <= valid_2_MPORT_211_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_215_en & valid_2_MPORT_215_mask) begin
      valid_2[valid_2_MPORT_215_addr] <= valid_2_MPORT_215_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_219_en & valid_2_MPORT_219_mask) begin
      valid_2[valid_2_MPORT_219_addr] <= valid_2_MPORT_219_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_223_en & valid_2_MPORT_223_mask) begin
      valid_2[valid_2_MPORT_223_addr] <= valid_2_MPORT_223_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_227_en & valid_2_MPORT_227_mask) begin
      valid_2[valid_2_MPORT_227_addr] <= valid_2_MPORT_227_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_231_en & valid_2_MPORT_231_mask) begin
      valid_2[valid_2_MPORT_231_addr] <= valid_2_MPORT_231_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_235_en & valid_2_MPORT_235_mask) begin
      valid_2[valid_2_MPORT_235_addr] <= valid_2_MPORT_235_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_239_en & valid_2_MPORT_239_mask) begin
      valid_2[valid_2_MPORT_239_addr] <= valid_2_MPORT_239_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_243_en & valid_2_MPORT_243_mask) begin
      valid_2[valid_2_MPORT_243_addr] <= valid_2_MPORT_243_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_247_en & valid_2_MPORT_247_mask) begin
      valid_2[valid_2_MPORT_247_addr] <= valid_2_MPORT_247_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_251_en & valid_2_MPORT_251_mask) begin
      valid_2[valid_2_MPORT_251_addr] <= valid_2_MPORT_251_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_255_en & valid_2_MPORT_255_mask) begin
      valid_2[valid_2_MPORT_255_addr] <= valid_2_MPORT_255_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_259_en & valid_2_MPORT_259_mask) begin
      valid_2[valid_2_MPORT_259_addr] <= valid_2_MPORT_259_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_2_MPORT_263_en & valid_2_MPORT_263_mask) begin
      valid_2[valid_2_MPORT_263_addr] <= valid_2_MPORT_263_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_71_en & valid_3_MPORT_71_mask) begin
      valid_3[valid_3_MPORT_71_addr] <= valid_3_MPORT_71_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_267_en & valid_3_MPORT_267_mask) begin
      valid_3[valid_3_MPORT_267_addr] <= valid_3_MPORT_267_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_271_en & valid_3_MPORT_271_mask) begin
      valid_3[valid_3_MPORT_271_addr] <= valid_3_MPORT_271_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_275_en & valid_3_MPORT_275_mask) begin
      valid_3[valid_3_MPORT_275_addr] <= valid_3_MPORT_275_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_279_en & valid_3_MPORT_279_mask) begin
      valid_3[valid_3_MPORT_279_addr] <= valid_3_MPORT_279_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_283_en & valid_3_MPORT_283_mask) begin
      valid_3[valid_3_MPORT_283_addr] <= valid_3_MPORT_283_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_287_en & valid_3_MPORT_287_mask) begin
      valid_3[valid_3_MPORT_287_addr] <= valid_3_MPORT_287_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_291_en & valid_3_MPORT_291_mask) begin
      valid_3[valid_3_MPORT_291_addr] <= valid_3_MPORT_291_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_295_en & valid_3_MPORT_295_mask) begin
      valid_3[valid_3_MPORT_295_addr] <= valid_3_MPORT_295_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_299_en & valid_3_MPORT_299_mask) begin
      valid_3[valid_3_MPORT_299_addr] <= valid_3_MPORT_299_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_303_en & valid_3_MPORT_303_mask) begin
      valid_3[valid_3_MPORT_303_addr] <= valid_3_MPORT_303_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_307_en & valid_3_MPORT_307_mask) begin
      valid_3[valid_3_MPORT_307_addr] <= valid_3_MPORT_307_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_311_en & valid_3_MPORT_311_mask) begin
      valid_3[valid_3_MPORT_311_addr] <= valid_3_MPORT_311_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_315_en & valid_3_MPORT_315_mask) begin
      valid_3[valid_3_MPORT_315_addr] <= valid_3_MPORT_315_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_319_en & valid_3_MPORT_319_mask) begin
      valid_3[valid_3_MPORT_319_addr] <= valid_3_MPORT_319_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_323_en & valid_3_MPORT_323_mask) begin
      valid_3[valid_3_MPORT_323_addr] <= valid_3_MPORT_323_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (valid_3_MPORT_327_en & valid_3_MPORT_327_mask) begin
      valid_3[valid_3_MPORT_327_addr] <= valid_3_MPORT_327_data; // @[BranchTargetBuffer.scala 102:20]
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_0 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_0 <= _GEN_1936;
        end else begin
          plru0_0 <= _GEN_1888;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_0 <= _GEN_2487;
      end else begin
        plru0_0 <= _GEN_2439;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_0 <= _GEN_1281;
      end else begin
        plru0_0 <= _GEN_1230;
      end
    end else begin
      plru0_0 <= _GEN_1230;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_1 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_1 <= _GEN_1937;
        end else begin
          plru0_1 <= _GEN_1889;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_1 <= _GEN_2488;
      end else begin
        plru0_1 <= _GEN_2440;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_1 <= _GEN_1282;
      end else begin
        plru0_1 <= _GEN_1231;
      end
    end else begin
      plru0_1 <= _GEN_1231;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_2 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_2 <= _GEN_1938;
        end else begin
          plru0_2 <= _GEN_1890;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_2 <= _GEN_2489;
      end else begin
        plru0_2 <= _GEN_2441;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_2 <= _GEN_1283;
      end else begin
        plru0_2 <= _GEN_1232;
      end
    end else begin
      plru0_2 <= _GEN_1232;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_3 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_3 <= _GEN_1939;
        end else begin
          plru0_3 <= _GEN_1891;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_3 <= _GEN_2490;
      end else begin
        plru0_3 <= _GEN_2442;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_3 <= _GEN_1284;
      end else begin
        plru0_3 <= _GEN_1233;
      end
    end else begin
      plru0_3 <= _GEN_1233;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_4 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_4 <= _GEN_1940;
        end else begin
          plru0_4 <= _GEN_1892;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_4 <= _GEN_2491;
      end else begin
        plru0_4 <= _GEN_2443;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_4 <= _GEN_1285;
      end else begin
        plru0_4 <= _GEN_1234;
      end
    end else begin
      plru0_4 <= _GEN_1234;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_5 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_5 <= _GEN_1941;
        end else begin
          plru0_5 <= _GEN_1893;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_5 <= _GEN_2492;
      end else begin
        plru0_5 <= _GEN_2444;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_5 <= _GEN_1286;
      end else begin
        plru0_5 <= _GEN_1235;
      end
    end else begin
      plru0_5 <= _GEN_1235;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_6 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_6 <= _GEN_1942;
        end else begin
          plru0_6 <= _GEN_1894;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_6 <= _GEN_2493;
      end else begin
        plru0_6 <= _GEN_2445;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_6 <= _GEN_1287;
      end else begin
        plru0_6 <= _GEN_1236;
      end
    end else begin
      plru0_6 <= _GEN_1236;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_7 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_7 <= _GEN_1943;
        end else begin
          plru0_7 <= _GEN_1895;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_7 <= _GEN_2494;
      end else begin
        plru0_7 <= _GEN_2446;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_7 <= _GEN_1288;
      end else begin
        plru0_7 <= _GEN_1237;
      end
    end else begin
      plru0_7 <= _GEN_1237;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_8 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_8 <= _GEN_1944;
        end else begin
          plru0_8 <= _GEN_1896;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_8 <= _GEN_2495;
      end else begin
        plru0_8 <= _GEN_2447;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_8 <= _GEN_1289;
      end else begin
        plru0_8 <= _GEN_1238;
      end
    end else begin
      plru0_8 <= _GEN_1238;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_9 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_9 <= _GEN_1945;
        end else begin
          plru0_9 <= _GEN_1897;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_9 <= _GEN_2496;
      end else begin
        plru0_9 <= _GEN_2448;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_9 <= _GEN_1290;
      end else begin
        plru0_9 <= _GEN_1239;
      end
    end else begin
      plru0_9 <= _GEN_1239;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_10 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_10 <= _GEN_1946;
        end else begin
          plru0_10 <= _GEN_1898;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_10 <= _GEN_2497;
      end else begin
        plru0_10 <= _GEN_2449;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_10 <= _GEN_1291;
      end else begin
        plru0_10 <= _GEN_1240;
      end
    end else begin
      plru0_10 <= _GEN_1240;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_11 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_11 <= _GEN_1947;
        end else begin
          plru0_11 <= _GEN_1899;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_11 <= _GEN_2498;
      end else begin
        plru0_11 <= _GEN_2450;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_11 <= _GEN_1292;
      end else begin
        plru0_11 <= _GEN_1241;
      end
    end else begin
      plru0_11 <= _GEN_1241;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_12 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_12 <= _GEN_1948;
        end else begin
          plru0_12 <= _GEN_1900;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_12 <= _GEN_2499;
      end else begin
        plru0_12 <= _GEN_2451;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_12 <= _GEN_1293;
      end else begin
        plru0_12 <= _GEN_1242;
      end
    end else begin
      plru0_12 <= _GEN_1242;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_13 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_13 <= _GEN_1949;
        end else begin
          plru0_13 <= _GEN_1901;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_13 <= _GEN_2500;
      end else begin
        plru0_13 <= _GEN_2452;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_13 <= _GEN_1294;
      end else begin
        plru0_13 <= _GEN_1243;
      end
    end else begin
      plru0_13 <= _GEN_1243;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_14 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_14 <= _GEN_1950;
        end else begin
          plru0_14 <= _GEN_1902;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_14 <= _GEN_2501;
      end else begin
        plru0_14 <= _GEN_2453;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_14 <= _GEN_1295;
      end else begin
        plru0_14 <= _GEN_1244;
      end
    end else begin
      plru0_14 <= _GEN_1244;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 107:22]
      plru0_15 <= 1'h0; // @[BranchTargetBuffer.scala 107:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru0_15 <= _GEN_1951;
        end else begin
          plru0_15 <= _GEN_1903;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru0_15 <= _GEN_2502;
      end else begin
        plru0_15 <= _GEN_2454;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru0_15 <= _GEN_1296;
      end else begin
        plru0_15 <= _GEN_1245;
      end
    end else begin
      plru0_15 <= _GEN_1245;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_0 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_0 <= _GEN_1678;
        end else begin
          plru1_0 <= _GEN_1630;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_0 <= _GEN_2227;
      end else begin
        plru1_0 <= _GEN_2179;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_0 <= _GEN_933;
      end else begin
        plru1_0 <= _GEN_882;
      end
    end else begin
      plru1_0 <= _GEN_882;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_1 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_1 <= _GEN_1679;
        end else begin
          plru1_1 <= _GEN_1631;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_1 <= _GEN_2228;
      end else begin
        plru1_1 <= _GEN_2180;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_1 <= _GEN_934;
      end else begin
        plru1_1 <= _GEN_883;
      end
    end else begin
      plru1_1 <= _GEN_883;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_2 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_2 <= _GEN_1680;
        end else begin
          plru1_2 <= _GEN_1632;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_2 <= _GEN_2229;
      end else begin
        plru1_2 <= _GEN_2181;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_2 <= _GEN_935;
      end else begin
        plru1_2 <= _GEN_884;
      end
    end else begin
      plru1_2 <= _GEN_884;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_3 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_3 <= _GEN_1681;
        end else begin
          plru1_3 <= _GEN_1633;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_3 <= _GEN_2230;
      end else begin
        plru1_3 <= _GEN_2182;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_3 <= _GEN_936;
      end else begin
        plru1_3 <= _GEN_885;
      end
    end else begin
      plru1_3 <= _GEN_885;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_4 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_4 <= _GEN_1682;
        end else begin
          plru1_4 <= _GEN_1634;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_4 <= _GEN_2231;
      end else begin
        plru1_4 <= _GEN_2183;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_4 <= _GEN_937;
      end else begin
        plru1_4 <= _GEN_886;
      end
    end else begin
      plru1_4 <= _GEN_886;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_5 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_5 <= _GEN_1683;
        end else begin
          plru1_5 <= _GEN_1635;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_5 <= _GEN_2232;
      end else begin
        plru1_5 <= _GEN_2184;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_5 <= _GEN_938;
      end else begin
        plru1_5 <= _GEN_887;
      end
    end else begin
      plru1_5 <= _GEN_887;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_6 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_6 <= _GEN_1684;
        end else begin
          plru1_6 <= _GEN_1636;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_6 <= _GEN_2233;
      end else begin
        plru1_6 <= _GEN_2185;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_6 <= _GEN_939;
      end else begin
        plru1_6 <= _GEN_888;
      end
    end else begin
      plru1_6 <= _GEN_888;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_7 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_7 <= _GEN_1685;
        end else begin
          plru1_7 <= _GEN_1637;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_7 <= _GEN_2234;
      end else begin
        plru1_7 <= _GEN_2186;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_7 <= _GEN_940;
      end else begin
        plru1_7 <= _GEN_889;
      end
    end else begin
      plru1_7 <= _GEN_889;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_8 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_8 <= _GEN_1686;
        end else begin
          plru1_8 <= _GEN_1638;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_8 <= _GEN_2235;
      end else begin
        plru1_8 <= _GEN_2187;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_8 <= _GEN_941;
      end else begin
        plru1_8 <= _GEN_890;
      end
    end else begin
      plru1_8 <= _GEN_890;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_9 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_9 <= _GEN_1687;
        end else begin
          plru1_9 <= _GEN_1639;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_9 <= _GEN_2236;
      end else begin
        plru1_9 <= _GEN_2188;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_9 <= _GEN_942;
      end else begin
        plru1_9 <= _GEN_891;
      end
    end else begin
      plru1_9 <= _GEN_891;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_10 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_10 <= _GEN_1688;
        end else begin
          plru1_10 <= _GEN_1640;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_10 <= _GEN_2237;
      end else begin
        plru1_10 <= _GEN_2189;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_10 <= _GEN_943;
      end else begin
        plru1_10 <= _GEN_892;
      end
    end else begin
      plru1_10 <= _GEN_892;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_11 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_11 <= _GEN_1689;
        end else begin
          plru1_11 <= _GEN_1641;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_11 <= _GEN_2238;
      end else begin
        plru1_11 <= _GEN_2190;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_11 <= _GEN_944;
      end else begin
        plru1_11 <= _GEN_893;
      end
    end else begin
      plru1_11 <= _GEN_893;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_12 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_12 <= _GEN_1690;
        end else begin
          plru1_12 <= _GEN_1642;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_12 <= _GEN_2239;
      end else begin
        plru1_12 <= _GEN_2191;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_12 <= _GEN_945;
      end else begin
        plru1_12 <= _GEN_894;
      end
    end else begin
      plru1_12 <= _GEN_894;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_13 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_13 <= _GEN_1691;
        end else begin
          plru1_13 <= _GEN_1643;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_13 <= _GEN_2240;
      end else begin
        plru1_13 <= _GEN_2192;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_13 <= _GEN_946;
      end else begin
        plru1_13 <= _GEN_895;
      end
    end else begin
      plru1_13 <= _GEN_895;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_14 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_14 <= _GEN_1692;
        end else begin
          plru1_14 <= _GEN_1644;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_14 <= _GEN_2241;
      end else begin
        plru1_14 <= _GEN_2193;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_14 <= _GEN_947;
      end else begin
        plru1_14 <= _GEN_896;
      end
    end else begin
      plru1_14 <= _GEN_896;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 109:22]
      plru1_15 <= 1'h0; // @[BranchTargetBuffer.scala 109:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h1) begin // @[BranchTargetBuffer.scala 175:30]
          plru1_15 <= _GEN_1693;
        end else begin
          plru1_15 <= _GEN_1645;
        end
      end else if (replace_way == 2'h1) begin // @[BranchTargetBuffer.scala 187:36]
        plru1_15 <= _GEN_2242;
      end else begin
        plru1_15 <= _GEN_2194;
      end
    end else if (REG_13_1 & _WIRE_27_1_tag == REG_17) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_18) begin // @[BranchTargetBuffer.scala 137:35]
        plru1_15 <= _GEN_948;
      end else begin
        plru1_15 <= _GEN_897;
      end
    end else begin
      plru1_15 <= _GEN_897;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_0 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_0 <= _GEN_1968;
        end else begin
          plru2_0 <= _GEN_1920;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_0 <= _GEN_2519;
      end else begin
        plru2_0 <= _GEN_2471;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_0 <= _GEN_1313;
      end else begin
        plru2_0 <= _GEN_1262;
      end
    end else begin
      plru2_0 <= _GEN_1262;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_1 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_1 <= _GEN_1969;
        end else begin
          plru2_1 <= _GEN_1921;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_1 <= _GEN_2520;
      end else begin
        plru2_1 <= _GEN_2472;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_1 <= _GEN_1314;
      end else begin
        plru2_1 <= _GEN_1263;
      end
    end else begin
      plru2_1 <= _GEN_1263;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_2 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_2 <= _GEN_1970;
        end else begin
          plru2_2 <= _GEN_1922;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_2 <= _GEN_2521;
      end else begin
        plru2_2 <= _GEN_2473;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_2 <= _GEN_1315;
      end else begin
        plru2_2 <= _GEN_1264;
      end
    end else begin
      plru2_2 <= _GEN_1264;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_3 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_3 <= _GEN_1971;
        end else begin
          plru2_3 <= _GEN_1923;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_3 <= _GEN_2522;
      end else begin
        plru2_3 <= _GEN_2474;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_3 <= _GEN_1316;
      end else begin
        plru2_3 <= _GEN_1265;
      end
    end else begin
      plru2_3 <= _GEN_1265;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_4 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_4 <= _GEN_1972;
        end else begin
          plru2_4 <= _GEN_1924;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_4 <= _GEN_2523;
      end else begin
        plru2_4 <= _GEN_2475;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_4 <= _GEN_1317;
      end else begin
        plru2_4 <= _GEN_1266;
      end
    end else begin
      plru2_4 <= _GEN_1266;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_5 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_5 <= _GEN_1973;
        end else begin
          plru2_5 <= _GEN_1925;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_5 <= _GEN_2524;
      end else begin
        plru2_5 <= _GEN_2476;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_5 <= _GEN_1318;
      end else begin
        plru2_5 <= _GEN_1267;
      end
    end else begin
      plru2_5 <= _GEN_1267;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_6 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_6 <= _GEN_1974;
        end else begin
          plru2_6 <= _GEN_1926;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_6 <= _GEN_2525;
      end else begin
        plru2_6 <= _GEN_2477;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_6 <= _GEN_1319;
      end else begin
        plru2_6 <= _GEN_1268;
      end
    end else begin
      plru2_6 <= _GEN_1268;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_7 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_7 <= _GEN_1975;
        end else begin
          plru2_7 <= _GEN_1927;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_7 <= _GEN_2526;
      end else begin
        plru2_7 <= _GEN_2478;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_7 <= _GEN_1320;
      end else begin
        plru2_7 <= _GEN_1269;
      end
    end else begin
      plru2_7 <= _GEN_1269;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_8 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_8 <= _GEN_1976;
        end else begin
          plru2_8 <= _GEN_1928;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_8 <= _GEN_2527;
      end else begin
        plru2_8 <= _GEN_2479;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_8 <= _GEN_1321;
      end else begin
        plru2_8 <= _GEN_1270;
      end
    end else begin
      plru2_8 <= _GEN_1270;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_9 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_9 <= _GEN_1977;
        end else begin
          plru2_9 <= _GEN_1929;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_9 <= _GEN_2528;
      end else begin
        plru2_9 <= _GEN_2480;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_9 <= _GEN_1322;
      end else begin
        plru2_9 <= _GEN_1271;
      end
    end else begin
      plru2_9 <= _GEN_1271;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_10 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_10 <= _GEN_1978;
        end else begin
          plru2_10 <= _GEN_1930;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_10 <= _GEN_2529;
      end else begin
        plru2_10 <= _GEN_2481;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_10 <= _GEN_1323;
      end else begin
        plru2_10 <= _GEN_1272;
      end
    end else begin
      plru2_10 <= _GEN_1272;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_11 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_11 <= _GEN_1979;
        end else begin
          plru2_11 <= _GEN_1931;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_11 <= _GEN_2530;
      end else begin
        plru2_11 <= _GEN_2482;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_11 <= _GEN_1324;
      end else begin
        plru2_11 <= _GEN_1273;
      end
    end else begin
      plru2_11 <= _GEN_1273;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_12 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_12 <= _GEN_1980;
        end else begin
          plru2_12 <= _GEN_1932;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_12 <= _GEN_2531;
      end else begin
        plru2_12 <= _GEN_2483;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_12 <= _GEN_1325;
      end else begin
        plru2_12 <= _GEN_1274;
      end
    end else begin
      plru2_12 <= _GEN_1274;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_13 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_13 <= _GEN_1981;
        end else begin
          plru2_13 <= _GEN_1933;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_13 <= _GEN_2532;
      end else begin
        plru2_13 <= _GEN_2484;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_13 <= _GEN_1326;
      end else begin
        plru2_13 <= _GEN_1275;
      end
    end else begin
      plru2_13 <= _GEN_1275;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_14 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_14 <= _GEN_1982;
        end else begin
          plru2_14 <= _GEN_1934;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_14 <= _GEN_2533;
      end else begin
        plru2_14 <= _GEN_2485;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_14 <= _GEN_1327;
      end else begin
        plru2_14 <= _GEN_1276;
      end
    end else begin
      plru2_14 <= _GEN_1276;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 111:22]
      plru2_15 <= 1'h0; // @[BranchTargetBuffer.scala 111:22]
    end else if (REG_30) begin // @[BranchTargetBuffer.scala 172:26]
      if (w_hit) begin // @[BranchTargetBuffer.scala 173:18]
        if (w_way == 2'h3) begin // @[BranchTargetBuffer.scala 175:30]
          plru2_15 <= _GEN_1983;
        end else begin
          plru2_15 <= _GEN_1935;
        end
      end else if (replace_way == 2'h3) begin // @[BranchTargetBuffer.scala 187:36]
        plru2_15 <= _GEN_2534;
      end else begin
        plru2_15 <= _GEN_2486;
      end
    end else if (REG_13_3 & _WIRE_27_3_tag == REG_23) begin // @[BranchTargetBuffer.scala 133:66]
      if (REG_24) begin // @[BranchTargetBuffer.scala 137:35]
        plru2_15 <= _GEN_1328;
      end else begin
        plru2_15 <= _GEN_1277;
      end
    end else begin
      plru2_15 <= _GEN_1277;
    end
    if (reset) begin // @[BranchTargetBuffer.scala 124:25]
      REG__0 <= 1'h0; // @[BranchTargetBuffer.scala 124:25]
    end else begin
      REG__0 <= valid_0_MPORT_3_data; // @[BranchTargetBuffer.scala 132:17]
    end
    if (reset) begin // @[BranchTargetBuffer.scala 124:25]
      REG__1 <= 1'h0; // @[BranchTargetBuffer.scala 124:25]
    end else begin
      REG__1 <= valid_1_MPORT_7_data; // @[BranchTargetBuffer.scala 132:17]
    end
    if (reset) begin // @[BranchTargetBuffer.scala 124:25]
      REG__2 <= 1'h0; // @[BranchTargetBuffer.scala 124:25]
    end else begin
      REG__2 <= valid_2_MPORT_11_data; // @[BranchTargetBuffer.scala 132:17]
    end
    if (reset) begin // @[BranchTargetBuffer.scala 124:25]
      REG__3 <= 1'h0; // @[BranchTargetBuffer.scala 124:25]
    end else begin
      REG__3 <= valid_3_MPORT_15_data; // @[BranchTargetBuffer.scala 132:17]
    end
    REG_1 <= io_rtag_0; // @[BranchTargetBuffer.scala 133:51]
    REG_2 <= io_ren_0; // @[BranchTargetBuffer.scala 137:22]
    REG_3 <= io_raddr_0; // @[BranchTargetBuffer.scala 138:33]
    REG_4 <= io_rtag_0; // @[BranchTargetBuffer.scala 133:51]
    REG_5 <= io_ren_0; // @[BranchTargetBuffer.scala 137:22]
    REG_6 <= io_raddr_0; // @[BranchTargetBuffer.scala 138:33]
    REG_7 <= io_rtag_0; // @[BranchTargetBuffer.scala 133:51]
    REG_8 <= io_ren_0; // @[BranchTargetBuffer.scala 137:22]
    REG_9 <= io_raddr_0; // @[BranchTargetBuffer.scala 138:33]
    REG_10 <= io_rtag_0; // @[BranchTargetBuffer.scala 133:51]
    REG_11 <= io_ren_0; // @[BranchTargetBuffer.scala 137:22]
    REG_12 <= io_raddr_0; // @[BranchTargetBuffer.scala 138:33]
    if (reset) begin // @[BranchTargetBuffer.scala 124:25]
      REG_13_0 <= 1'h0; // @[BranchTargetBuffer.scala 124:25]
    end else begin
      REG_13_0 <= valid_0_MPORT_19_data; // @[BranchTargetBuffer.scala 132:17]
    end
    if (reset) begin // @[BranchTargetBuffer.scala 124:25]
      REG_13_1 <= 1'h0; // @[BranchTargetBuffer.scala 124:25]
    end else begin
      REG_13_1 <= valid_1_MPORT_23_data; // @[BranchTargetBuffer.scala 132:17]
    end
    if (reset) begin // @[BranchTargetBuffer.scala 124:25]
      REG_13_2 <= 1'h0; // @[BranchTargetBuffer.scala 124:25]
    end else begin
      REG_13_2 <= valid_2_MPORT_27_data; // @[BranchTargetBuffer.scala 132:17]
    end
    if (reset) begin // @[BranchTargetBuffer.scala 124:25]
      REG_13_3 <= 1'h0; // @[BranchTargetBuffer.scala 124:25]
    end else begin
      REG_13_3 <= valid_3_MPORT_31_data; // @[BranchTargetBuffer.scala 132:17]
    end
    REG_14 <= io_rtag_1; // @[BranchTargetBuffer.scala 133:51]
    REG_15 <= io_ren_1; // @[BranchTargetBuffer.scala 137:22]
    REG_16 <= io_raddr_1; // @[BranchTargetBuffer.scala 138:33]
    REG_17 <= io_rtag_1; // @[BranchTargetBuffer.scala 133:51]
    REG_18 <= io_ren_1; // @[BranchTargetBuffer.scala 137:22]
    REG_19 <= io_raddr_1; // @[BranchTargetBuffer.scala 138:33]
    REG_20 <= io_rtag_1; // @[BranchTargetBuffer.scala 133:51]
    REG_21 <= io_ren_1; // @[BranchTargetBuffer.scala 137:22]
    REG_22 <= io_raddr_1; // @[BranchTargetBuffer.scala 138:33]
    REG_23 <= io_rtag_1; // @[BranchTargetBuffer.scala 133:51]
    REG_24 <= io_ren_1; // @[BranchTargetBuffer.scala 137:22]
    REG_25 <= io_raddr_1; // @[BranchTargetBuffer.scala 138:33]
    if (reset) begin // @[BranchTargetBuffer.scala 157:25]
      w_rvalid_0 <= 1'h0; // @[BranchTargetBuffer.scala 157:25]
    end else begin
      w_rvalid_0 <= valid_0_MPORT_34_data; // @[BranchTargetBuffer.scala 165:17]
    end
    if (reset) begin // @[BranchTargetBuffer.scala 157:25]
      w_rvalid_1 <= 1'h0; // @[BranchTargetBuffer.scala 157:25]
    end else begin
      w_rvalid_1 <= valid_1_MPORT_37_data; // @[BranchTargetBuffer.scala 165:17]
    end
    if (reset) begin // @[BranchTargetBuffer.scala 157:25]
      w_rvalid_2 <= 1'h0; // @[BranchTargetBuffer.scala 157:25]
    end else begin
      w_rvalid_2 <= valid_2_MPORT_40_data; // @[BranchTargetBuffer.scala 165:17]
    end
    if (reset) begin // @[BranchTargetBuffer.scala 157:25]
      w_rvalid_3 <= 1'h0; // @[BranchTargetBuffer.scala 157:25]
    end else begin
      w_rvalid_3 <= valid_3_MPORT_43_data; // @[BranchTargetBuffer.scala 165:17]
    end
    REG_26 <= io_wtag; // @[BranchTargetBuffer.scala 166:53]
    REG_27 <= io_wtag; // @[BranchTargetBuffer.scala 166:53]
    REG_28 <= io_wtag; // @[BranchTargetBuffer.scala 166:53]
    REG_29 <= io_wtag; // @[BranchTargetBuffer.scala 166:53]
    REG_30 <= io_wen; // @[BranchTargetBuffer.scala 172:16]
    REG_31 <= io_waddr; // @[BranchTargetBuffer.scala 176:35]
    REG_32 <= io_wtag; // @[BranchTargetBuffer.scala 149:20 150:14]
    REG_33 <= io_waddr; // @[BranchTargetBuffer.scala 177:38]
    REG_34 <= io_wtarget; // @[BranchTargetBuffer.scala 149:20 151:17]
    REG_37 <= io_waddr; // @[BranchTargetBuffer.scala 179:33]
    REG_38 <= io_waddr; // @[BranchTargetBuffer.scala 176:35]
    REG_39 <= io_wtag; // @[BranchTargetBuffer.scala 149:20 150:14]
    REG_40 <= io_waddr; // @[BranchTargetBuffer.scala 177:38]
    REG_41 <= io_wtarget; // @[BranchTargetBuffer.scala 149:20 151:17]
    REG_44 <= io_waddr; // @[BranchTargetBuffer.scala 179:33]
    REG_45 <= io_waddr; // @[BranchTargetBuffer.scala 176:35]
    REG_46 <= io_wtag; // @[BranchTargetBuffer.scala 149:20 150:14]
    REG_47 <= io_waddr; // @[BranchTargetBuffer.scala 177:38]
    REG_48 <= io_wtarget; // @[BranchTargetBuffer.scala 149:20 151:17]
    REG_51 <= io_waddr; // @[BranchTargetBuffer.scala 179:33]
    REG_52 <= io_waddr; // @[BranchTargetBuffer.scala 176:35]
    REG_53 <= io_wtag; // @[BranchTargetBuffer.scala 149:20 150:14]
    REG_54 <= io_waddr; // @[BranchTargetBuffer.scala 177:38]
    REG_55 <= io_wtarget; // @[BranchTargetBuffer.scala 149:20 151:17]
    REG_58 <= io_waddr; // @[BranchTargetBuffer.scala 179:33]
    REG_59 <= io_waddr; // @[BranchTargetBuffer.scala 188:35]
    REG_60 <= io_wtag; // @[BranchTargetBuffer.scala 149:20 150:14]
    REG_61 <= io_waddr; // @[BranchTargetBuffer.scala 189:38]
    REG_62 <= io_wtarget; // @[BranchTargetBuffer.scala 149:20 151:17]
    REG_65 <= io_waddr; // @[BranchTargetBuffer.scala 191:27]
    REG_66 <= io_waddr; // @[BranchTargetBuffer.scala 192:33]
    REG_67 <= io_waddr; // @[BranchTargetBuffer.scala 188:35]
    REG_68 <= io_wtag; // @[BranchTargetBuffer.scala 149:20 150:14]
    REG_69 <= io_waddr; // @[BranchTargetBuffer.scala 189:38]
    REG_70 <= io_wtarget; // @[BranchTargetBuffer.scala 149:20 151:17]
    REG_73 <= io_waddr; // @[BranchTargetBuffer.scala 191:27]
    REG_74 <= io_waddr; // @[BranchTargetBuffer.scala 192:33]
    REG_75 <= io_waddr; // @[BranchTargetBuffer.scala 188:35]
    REG_76 <= io_wtag; // @[BranchTargetBuffer.scala 149:20 150:14]
    REG_77 <= io_waddr; // @[BranchTargetBuffer.scala 189:38]
    REG_78 <= io_wtarget; // @[BranchTargetBuffer.scala 149:20 151:17]
    REG_81 <= io_waddr; // @[BranchTargetBuffer.scala 191:27]
    REG_82 <= io_waddr; // @[BranchTargetBuffer.scala 192:33]
    REG_83 <= io_waddr; // @[BranchTargetBuffer.scala 188:35]
    REG_84 <= io_wtag; // @[BranchTargetBuffer.scala 149:20 150:14]
    REG_85 <= io_waddr; // @[BranchTargetBuffer.scala 189:38]
    REG_86 <= io_wtarget; // @[BranchTargetBuffer.scala 149:20 151:17]
    REG_89 <= io_waddr; // @[BranchTargetBuffer.scala 191:27]
    REG_90 <= io_waddr; // @[BranchTargetBuffer.scala 192:33]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    btb_tag_0[initvar] = _RAND_0[25:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    btb_tag_1[initvar] = _RAND_7[25:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    btb_tag_2[initvar] = _RAND_14[25:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    btb_tag_3[initvar] = _RAND_21[25:0];
  _RAND_28 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    btb_target_0[initvar] = _RAND_28[31:0];
  _RAND_33 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    btb_target_1[initvar] = _RAND_33[31:0];
  _RAND_38 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    btb_target_2[initvar] = _RAND_38[31:0];
  _RAND_43 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    btb_target_3[initvar] = _RAND_43[31:0];
  _RAND_48 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    valid_0[initvar] = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    valid_1[initvar] = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    valid_2[initvar] = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    valid_3[initvar] = _RAND_51[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
//   btb_tag_0_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  btb_tag_0_MPORT_addr_pipe_0 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
//   btb_tag_0_MPORT_16_en_pipe_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  btb_tag_0_MPORT_16_addr_pipe_0 = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
//   btb_tag_0_MPORT_32_en_pipe_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  btb_tag_0_MPORT_32_addr_pipe_0 = _RAND_6[3:0];
  _RAND_8 = {1{`RANDOM}};
//   btb_tag_1_MPORT_4_en_pipe_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  btb_tag_1_MPORT_4_addr_pipe_0 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
//   btb_tag_1_MPORT_20_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  btb_tag_1_MPORT_20_addr_pipe_0 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
//   btb_tag_1_MPORT_35_en_pipe_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  btb_tag_1_MPORT_35_addr_pipe_0 = _RAND_13[3:0];
  _RAND_15 = {1{`RANDOM}};
//   btb_tag_2_MPORT_8_en_pipe_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  btb_tag_2_MPORT_8_addr_pipe_0 = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
//   btb_tag_2_MPORT_24_en_pipe_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  btb_tag_2_MPORT_24_addr_pipe_0 = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
//   btb_tag_2_MPORT_38_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  btb_tag_2_MPORT_38_addr_pipe_0 = _RAND_20[3:0];
  _RAND_22 = {1{`RANDOM}};
//   btb_tag_3_MPORT_12_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  btb_tag_3_MPORT_12_addr_pipe_0 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
//   btb_tag_3_MPORT_28_en_pipe_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  btb_tag_3_MPORT_28_addr_pipe_0 = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
//   btb_tag_3_MPORT_41_en_pipe_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  btb_tag_3_MPORT_41_addr_pipe_0 = _RAND_27[3:0];
  _RAND_29 = {1{`RANDOM}};
//   btb_target_0_MPORT_1_en_pipe_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  btb_target_0_MPORT_1_addr_pipe_0 = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
//   btb_target_0_MPORT_17_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  btb_target_0_MPORT_17_addr_pipe_0 = _RAND_32[3:0];
  _RAND_34 = {1{`RANDOM}};
//   btb_target_1_MPORT_5_en_pipe_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  btb_target_1_MPORT_5_addr_pipe_0 = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
//   btb_target_1_MPORT_21_en_pipe_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  btb_target_1_MPORT_21_addr_pipe_0 = _RAND_37[3:0];
  _RAND_39 = {1{`RANDOM}};
//   btb_target_2_MPORT_9_en_pipe_0 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  btb_target_2_MPORT_9_addr_pipe_0 = _RAND_40[3:0];
  _RAND_41 = {1{`RANDOM}};
//   btb_target_2_MPORT_25_en_pipe_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  btb_target_2_MPORT_25_addr_pipe_0 = _RAND_42[3:0];
  _RAND_44 = {1{`RANDOM}};
//   btb_target_3_MPORT_13_en_pipe_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  btb_target_3_MPORT_13_addr_pipe_0 = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
//   btb_target_3_MPORT_29_en_pipe_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  btb_target_3_MPORT_29_addr_pipe_0 = _RAND_47[3:0];
  _RAND_52 = {1{`RANDOM}};
  plru0_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  plru0_1 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  plru0_2 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  plru0_3 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  plru0_4 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  plru0_5 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  plru0_6 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  plru0_7 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  plru0_8 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  plru0_9 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  plru0_10 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  plru0_11 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  plru0_12 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  plru0_13 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  plru0_14 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  plru0_15 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  plru1_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  plru1_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  plru1_2 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  plru1_3 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  plru1_4 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  plru1_5 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  plru1_6 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  plru1_7 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  plru1_8 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  plru1_9 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  plru1_10 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  plru1_11 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  plru1_12 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  plru1_13 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  plru1_14 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  plru1_15 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  plru2_0 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  plru2_1 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  plru2_2 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  plru2_3 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  plru2_4 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  plru2_5 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  plru2_6 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  plru2_7 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  plru2_8 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  plru2_9 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  plru2_10 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  plru2_11 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  plru2_12 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  plru2_13 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  plru2_14 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  plru2_15 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  REG__0 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  REG__1 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  REG__2 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  REG__3 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  REG_1 = _RAND_104[25:0];
  _RAND_105 = {1{`RANDOM}};
  REG_2 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  REG_3 = _RAND_106[3:0];
  _RAND_107 = {1{`RANDOM}};
  REG_4 = _RAND_107[25:0];
  _RAND_108 = {1{`RANDOM}};
  REG_5 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  REG_6 = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  REG_7 = _RAND_110[25:0];
  _RAND_111 = {1{`RANDOM}};
  REG_8 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  REG_9 = _RAND_112[3:0];
  _RAND_113 = {1{`RANDOM}};
  REG_10 = _RAND_113[25:0];
  _RAND_114 = {1{`RANDOM}};
  REG_11 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  REG_12 = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  REG_13_0 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  REG_13_1 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  REG_13_2 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  REG_13_3 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  REG_14 = _RAND_120[25:0];
  _RAND_121 = {1{`RANDOM}};
  REG_15 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  REG_16 = _RAND_122[3:0];
  _RAND_123 = {1{`RANDOM}};
  REG_17 = _RAND_123[25:0];
  _RAND_124 = {1{`RANDOM}};
  REG_18 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  REG_19 = _RAND_125[3:0];
  _RAND_126 = {1{`RANDOM}};
  REG_20 = _RAND_126[25:0];
  _RAND_127 = {1{`RANDOM}};
  REG_21 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  REG_22 = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  REG_23 = _RAND_129[25:0];
  _RAND_130 = {1{`RANDOM}};
  REG_24 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  REG_25 = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  w_rvalid_0 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  w_rvalid_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  w_rvalid_2 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  w_rvalid_3 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  REG_26 = _RAND_136[25:0];
  _RAND_137 = {1{`RANDOM}};
  REG_27 = _RAND_137[25:0];
  _RAND_138 = {1{`RANDOM}};
  REG_28 = _RAND_138[25:0];
  _RAND_139 = {1{`RANDOM}};
  REG_29 = _RAND_139[25:0];
  _RAND_140 = {1{`RANDOM}};
  REG_30 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  REG_31 = _RAND_141[3:0];
  _RAND_142 = {1{`RANDOM}};
  REG_32 = _RAND_142[25:0];
  _RAND_143 = {1{`RANDOM}};
  REG_33 = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  REG_34 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  REG_37 = _RAND_145[3:0];
  _RAND_146 = {1{`RANDOM}};
  REG_38 = _RAND_146[3:0];
  _RAND_147 = {1{`RANDOM}};
  REG_39 = _RAND_147[25:0];
  _RAND_148 = {1{`RANDOM}};
  REG_40 = _RAND_148[3:0];
  _RAND_149 = {1{`RANDOM}};
  REG_41 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  REG_44 = _RAND_150[3:0];
  _RAND_151 = {1{`RANDOM}};
  REG_45 = _RAND_151[3:0];
  _RAND_152 = {1{`RANDOM}};
  REG_46 = _RAND_152[25:0];
  _RAND_153 = {1{`RANDOM}};
  REG_47 = _RAND_153[3:0];
  _RAND_154 = {1{`RANDOM}};
  REG_48 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  REG_51 = _RAND_155[3:0];
  _RAND_156 = {1{`RANDOM}};
  REG_52 = _RAND_156[3:0];
  _RAND_157 = {1{`RANDOM}};
  REG_53 = _RAND_157[25:0];
  _RAND_158 = {1{`RANDOM}};
  REG_54 = _RAND_158[3:0];
  _RAND_159 = {1{`RANDOM}};
  REG_55 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  REG_58 = _RAND_160[3:0];
  _RAND_161 = {1{`RANDOM}};
  REG_59 = _RAND_161[3:0];
  _RAND_162 = {1{`RANDOM}};
  REG_60 = _RAND_162[25:0];
  _RAND_163 = {1{`RANDOM}};
  REG_61 = _RAND_163[3:0];
  _RAND_164 = {1{`RANDOM}};
  REG_62 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  REG_65 = _RAND_165[3:0];
  _RAND_166 = {1{`RANDOM}};
  REG_66 = _RAND_166[3:0];
  _RAND_167 = {1{`RANDOM}};
  REG_67 = _RAND_167[3:0];
  _RAND_168 = {1{`RANDOM}};
  REG_68 = _RAND_168[25:0];
  _RAND_169 = {1{`RANDOM}};
  REG_69 = _RAND_169[3:0];
  _RAND_170 = {1{`RANDOM}};
  REG_70 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  REG_73 = _RAND_171[3:0];
  _RAND_172 = {1{`RANDOM}};
  REG_74 = _RAND_172[3:0];
  _RAND_173 = {1{`RANDOM}};
  REG_75 = _RAND_173[3:0];
  _RAND_174 = {1{`RANDOM}};
  REG_76 = _RAND_174[25:0];
  _RAND_175 = {1{`RANDOM}};
  REG_77 = _RAND_175[3:0];
  _RAND_176 = {1{`RANDOM}};
  REG_78 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  REG_81 = _RAND_177[3:0];
  _RAND_178 = {1{`RANDOM}};
  REG_82 = _RAND_178[3:0];
  _RAND_179 = {1{`RANDOM}};
  REG_83 = _RAND_179[3:0];
  _RAND_180 = {1{`RANDOM}};
  REG_84 = _RAND_180[25:0];
  _RAND_181 = {1{`RANDOM}};
  REG_85 = _RAND_181[3:0];
  _RAND_182 = {1{`RANDOM}};
  REG_86 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  REG_89 = _RAND_183[3:0];
  _RAND_184 = {1{`RANDOM}};
  REG_90 = _RAND_184[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_BranchPredictor(
  input         clock,
  input         reset,
  input  [31:0] io_pc,
  input         io_pc_en,
  input         io_jmp_packet_valid,
  input  [31:0] io_jmp_packet_inst_pc,
  input         io_jmp_packet_jmp,
  input  [31:0] io_jmp_packet_jmp_pc,
  input         io_jmp_packet_mis,
  input         io_jmp_packet_sys,
  output        io_pred_br_0,
  output        io_pred_br_1,
  output [31:0] io_pred_bpc,
  output        io_pred_valid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [5:0] bht [0:63]; // @[BranchPredictor.scala 68:16]
//   wire  bht_bht_rdata_0_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_bht_rdata_0_addr; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_bht_rdata_0_data; // @[BranchPredictor.scala 68:16]
//   wire  bht_bht_rdata_1_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_bht_rdata_1_addr; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_bht_rdata_1_data; // @[BranchPredictor.scala 68:16]
//   wire  bht_bht_wrdata_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_bht_wrdata_addr; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_bht_wrdata_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_1_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_1_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_1_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_1_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_2_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_2_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_2_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_2_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_3_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_3_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_3_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_3_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_4_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_4_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_4_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_4_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_5_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_5_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_5_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_5_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_6_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_6_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_6_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_6_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_7_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_7_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_7_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_7_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_8_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_8_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_8_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_8_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_9_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_9_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_9_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_9_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_10_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_10_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_10_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_10_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_11_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_11_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_11_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_11_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_12_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_12_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_12_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_12_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_13_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_13_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_13_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_13_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_14_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_14_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_14_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_14_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_15_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_15_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_15_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_15_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_16_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_16_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_16_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_16_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_17_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_17_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_17_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_17_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_18_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_18_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_18_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_18_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_19_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_19_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_19_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_19_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_20_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_20_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_20_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_20_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_21_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_21_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_21_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_21_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_22_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_22_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_22_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_22_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_23_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_23_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_23_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_23_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_24_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_24_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_24_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_24_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_25_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_25_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_25_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_25_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_26_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_26_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_26_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_26_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_27_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_27_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_27_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_27_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_28_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_28_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_28_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_28_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_29_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_29_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_29_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_29_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_30_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_30_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_30_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_30_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_31_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_31_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_31_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_31_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_32_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_32_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_32_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_32_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_33_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_33_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_33_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_33_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_34_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_34_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_34_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_34_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_35_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_35_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_35_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_35_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_36_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_36_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_36_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_36_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_37_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_37_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_37_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_37_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_38_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_38_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_38_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_38_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_39_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_39_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_39_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_39_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_40_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_40_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_40_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_40_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_41_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_41_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_41_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_41_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_42_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_42_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_42_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_42_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_43_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_43_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_43_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_43_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_44_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_44_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_44_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_44_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_45_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_45_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_45_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_45_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_46_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_46_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_46_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_46_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_47_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_47_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_47_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_47_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_48_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_48_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_48_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_48_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_49_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_49_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_49_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_49_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_50_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_50_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_50_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_50_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_51_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_51_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_51_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_51_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_52_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_52_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_52_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_52_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_53_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_53_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_53_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_53_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_54_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_54_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_54_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_54_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_55_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_55_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_55_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_55_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_56_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_56_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_56_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_56_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_57_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_57_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_57_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_57_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_58_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_58_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_58_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_58_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_59_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_59_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_59_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_59_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_60_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_60_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_60_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_60_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_61_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_61_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_61_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_61_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_62_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_62_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_62_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_62_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_63_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_63_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_63_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_63_en; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_64_data; // @[BranchPredictor.scala 68:16]
  wire [5:0] bht_MPORT_64_addr; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_64_mask; // @[BranchPredictor.scala 68:16]
  wire  bht_MPORT_64_en; // @[BranchPredictor.scala 68:16]
  wire  pht_clock; // @[BranchPredictor.scala 101:19]
  wire  pht_reset; // @[BranchPredictor.scala 101:19]
  wire [2:0] pht_io_rindex_0; // @[BranchPredictor.scala 101:19]
  wire [2:0] pht_io_rindex_1; // @[BranchPredictor.scala 101:19]
  wire [5:0] pht_io_raddr_0; // @[BranchPredictor.scala 101:19]
  wire [5:0] pht_io_raddr_1; // @[BranchPredictor.scala 101:19]
  wire  pht_io_rdirect_0; // @[BranchPredictor.scala 101:19]
  wire  pht_io_rdirect_1; // @[BranchPredictor.scala 101:19]
  wire [2:0] pht_io_windex; // @[BranchPredictor.scala 101:19]
  wire [5:0] pht_io_waddr; // @[BranchPredictor.scala 101:19]
  wire  pht_io_wen; // @[BranchPredictor.scala 101:19]
  wire  pht_io_wjmp; // @[BranchPredictor.scala 101:19]
  wire  btb_clock; // @[BranchPredictor.scala 121:19]
  wire  btb_reset; // @[BranchPredictor.scala 121:19]
  wire [3:0] btb_io_raddr_0; // @[BranchPredictor.scala 121:19]
  wire [3:0] btb_io_raddr_1; // @[BranchPredictor.scala 121:19]
  wire  btb_io_ren_0; // @[BranchPredictor.scala 121:19]
  wire  btb_io_ren_1; // @[BranchPredictor.scala 121:19]
  wire [25:0] btb_io_rtag_0; // @[BranchPredictor.scala 121:19]
  wire [25:0] btb_io_rtag_1; // @[BranchPredictor.scala 121:19]
  wire  btb_io_rhit_0; // @[BranchPredictor.scala 121:19]
  wire  btb_io_rhit_1; // @[BranchPredictor.scala 121:19]
  wire [31:0] btb_io_rtarget_0; // @[BranchPredictor.scala 121:19]
  wire [31:0] btb_io_rtarget_1; // @[BranchPredictor.scala 121:19]
  wire [3:0] btb_io_waddr; // @[BranchPredictor.scala 121:19]
  wire  btb_io_wen; // @[BranchPredictor.scala 121:19]
  wire [25:0] btb_io_wtag; // @[BranchPredictor.scala 121:19]
  wire [31:0] btb_io_wtarget; // @[BranchPredictor.scala 121:19]
  wire [31:0] pc_base = {io_pc[31:3],3'h0}; // @[Cat.scala 30:58]
  wire [32:0] _T_2 = {{1'd0}, pc_base}; // @[BranchPredictor.scala 50:22]
  wire [31:0] pc_0 = _T_2[31:0]; // @[BranchPredictor.scala 50:22]
  wire [31:0] pc_1 = pc_base + 32'h4; // @[BranchPredictor.scala 50:22]
  reg  pc_en_0; // @[BranchPredictor.scala 55:22]
  reg  pc_en_1; // @[BranchPredictor.scala 55:22]
  wire  _T_10 = ~io_jmp_packet_sys; // @[BranchPredictor.scala 62:46]
  wire  jmp_packet_valid = io_jmp_packet_valid & ~io_jmp_packet_sys; // @[BranchPredictor.scala 62:43]
  wire [5:0] bht_raddr_0 = pc_0[7:2]; // @[BranchPredictor.scala 69:34]
  wire [5:0] bht_raddr_1 = pc_1[7:2]; // @[BranchPredictor.scala 69:34]
  wire [5:0] bht_waddr = io_jmp_packet_inst_pc[7:2]; // @[BranchPredictor.scala 69:34]
  wire  btb_rhit_1 = btb_io_rhit_1;
  wire  btb_rhit_0 = btb_io_rhit_0;
  wire  pht_rdirect_1 = pht_io_rdirect_1;
  wire  pht_rdirect_0 = pht_io_rdirect_0;
  wire [31:0] _T_63 = io_jmp_packet_inst_pc + 32'h4; // @[BranchPredictor.scala 163:42]
  wire [31:0] _T_97 = io_jmp_packet_jmp ? io_jmp_packet_jmp_pc : _T_63; // @[BranchPredictor.scala 187:25]
  reg [31:0] REG_4; // @[BranchPredictor.scala 191:64]
  wire [31:0] btb_rtarget_0 = btb_io_rtarget_0;
  wire [31:0] _T_98 = btb_rhit_0 ? btb_rtarget_0 : REG_4; // @[BranchPredictor.scala 191:27]
  reg [31:0] REG_5; // @[BranchPredictor.scala 194:31]
  wire  _GEN_79 = pht_rdirect_0 & btb_rhit_0; // @[BranchPredictor.scala 189:29 190:20 193:20]
  wire [31:0] _GEN_80 = pht_rdirect_0 ? _T_98 : REG_5; // @[BranchPredictor.scala 189:29 191:21 194:21]
  wire  pred_br_0 = jmp_packet_valid & io_jmp_packet_mis ? 1'h0 : _GEN_79; // @[BranchPredictor.scala 185:47 186:18]
  wire [31:0] pred_bpc_0 = jmp_packet_valid & io_jmp_packet_mis ? _T_97 : _GEN_80; // @[BranchPredictor.scala 185:47 187:19]
  reg [31:0] REG_6; // @[BranchPredictor.scala 191:64]
  wire [31:0] btb_rtarget_1 = btb_io_rtarget_1;
  wire [31:0] _T_103 = btb_rhit_1 ? btb_rtarget_1 : REG_6; // @[BranchPredictor.scala 191:27]
  reg [31:0] REG_7; // @[BranchPredictor.scala 194:31]
  wire  _GEN_83 = pht_rdirect_1 & btb_rhit_1; // @[BranchPredictor.scala 189:29 190:20 193:20]
  wire [31:0] _GEN_84 = pht_rdirect_1 ? _T_103 : REG_7; // @[BranchPredictor.scala 189:29 191:21 194:21]
  wire  pred_br_1 = jmp_packet_valid & io_jmp_packet_mis ? 1'h0 : _GEN_83; // @[BranchPredictor.scala 185:47 186:18]
  wire [31:0] pred_bpc_1 = jmp_packet_valid & io_jmp_packet_mis ? _T_97 : _GEN_84; // @[BranchPredictor.scala 185:47 187:19]
  wire [1:0] _T_106 = {pred_br_1,pred_br_0}; // @[Cat.scala 30:58]
  wire [31:0] _T_108 = 2'h3 == _T_106 ? pred_bpc_0 : 32'h0; // @[Mux.scala 80:57]
  wire [31:0] _T_110 = 2'h1 == _T_106 ? pred_bpc_0 : _T_108; // @[Mux.scala 80:57]
  reg  REG_8; // @[BranchPredictor.scala 214:27]
  ysyx_210128_PatternHistoryTableLocal pht ( // @[BranchPredictor.scala 101:19]
    .clock(pht_clock),
    .reset(pht_reset),
    .io_rindex_0(pht_io_rindex_0),
    .io_rindex_1(pht_io_rindex_1),
    .io_raddr_0(pht_io_raddr_0),
    .io_raddr_1(pht_io_raddr_1),
    .io_rdirect_0(pht_io_rdirect_0),
    .io_rdirect_1(pht_io_rdirect_1),
    .io_windex(pht_io_windex),
    .io_waddr(pht_io_waddr),
    .io_wen(pht_io_wen),
    .io_wjmp(pht_io_wjmp)
  );
  ysyx_210128_BranchTargetBuffer4WayAssociative btb ( // @[BranchPredictor.scala 121:19]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_raddr_0(btb_io_raddr_0),
    .io_raddr_1(btb_io_raddr_1),
    .io_ren_0(btb_io_ren_0),
    .io_ren_1(btb_io_ren_1),
    .io_rtag_0(btb_io_rtag_0),
    .io_rtag_1(btb_io_rtag_1),
    .io_rhit_0(btb_io_rhit_0),
    .io_rhit_1(btb_io_rhit_1),
    .io_rtarget_0(btb_io_rtarget_0),
    .io_rtarget_1(btb_io_rtarget_1),
    .io_waddr(btb_io_waddr),
    .io_wen(btb_io_wen),
    .io_wtag(btb_io_wtag),
    .io_wtarget(btb_io_wtarget)
  );
//   assign bht_bht_rdata_0_en = 1'h1;
  assign bht_bht_rdata_0_addr = pc_0[7:2];
  assign bht_bht_rdata_0_data = bht[bht_bht_rdata_0_addr]; // @[BranchPredictor.scala 68:16]
//   assign bht_bht_rdata_1_en = 1'h1;
  assign bht_bht_rdata_1_addr = pc_1[7:2];
  assign bht_bht_rdata_1_data = bht[bht_bht_rdata_1_addr]; // @[BranchPredictor.scala 68:16]
//   assign bht_bht_wrdata_en = 1'h1;
  assign bht_bht_wrdata_addr = io_jmp_packet_inst_pc[7:2];
  assign bht_bht_wrdata_data = bht[bht_bht_wrdata_addr]; // @[BranchPredictor.scala 68:16]
  assign bht_MPORT_data = {io_jmp_packet_jmp,bht_bht_wrdata_data[5:1]};
  assign bht_MPORT_addr = io_jmp_packet_inst_pc[7:2];
  assign bht_MPORT_mask = 1'h1;
  assign bht_MPORT_en = io_jmp_packet_valid & _T_10;
  assign bht_MPORT_1_data = 6'h0;
  assign bht_MPORT_1_addr = 6'h0;
  assign bht_MPORT_1_mask = 1'h1;
  assign bht_MPORT_1_en = reset;
  assign bht_MPORT_2_data = 6'h0;
  assign bht_MPORT_2_addr = 6'h1;
  assign bht_MPORT_2_mask = 1'h1;
  assign bht_MPORT_2_en = reset;
  assign bht_MPORT_3_data = 6'h0;
  assign bht_MPORT_3_addr = 6'h2;
  assign bht_MPORT_3_mask = 1'h1;
  assign bht_MPORT_3_en = reset;
  assign bht_MPORT_4_data = 6'h0;
  assign bht_MPORT_4_addr = 6'h3;
  assign bht_MPORT_4_mask = 1'h1;
  assign bht_MPORT_4_en = reset;
  assign bht_MPORT_5_data = 6'h0;
  assign bht_MPORT_5_addr = 6'h4;
  assign bht_MPORT_5_mask = 1'h1;
  assign bht_MPORT_5_en = reset;
  assign bht_MPORT_6_data = 6'h0;
  assign bht_MPORT_6_addr = 6'h5;
  assign bht_MPORT_6_mask = 1'h1;
  assign bht_MPORT_6_en = reset;
  assign bht_MPORT_7_data = 6'h0;
  assign bht_MPORT_7_addr = 6'h6;
  assign bht_MPORT_7_mask = 1'h1;
  assign bht_MPORT_7_en = reset;
  assign bht_MPORT_8_data = 6'h0;
  assign bht_MPORT_8_addr = 6'h7;
  assign bht_MPORT_8_mask = 1'h1;
  assign bht_MPORT_8_en = reset;
  assign bht_MPORT_9_data = 6'h0;
  assign bht_MPORT_9_addr = 6'h8;
  assign bht_MPORT_9_mask = 1'h1;
  assign bht_MPORT_9_en = reset;
  assign bht_MPORT_10_data = 6'h0;
  assign bht_MPORT_10_addr = 6'h9;
  assign bht_MPORT_10_mask = 1'h1;
  assign bht_MPORT_10_en = reset;
  assign bht_MPORT_11_data = 6'h0;
  assign bht_MPORT_11_addr = 6'ha;
  assign bht_MPORT_11_mask = 1'h1;
  assign bht_MPORT_11_en = reset;
  assign bht_MPORT_12_data = 6'h0;
  assign bht_MPORT_12_addr = 6'hb;
  assign bht_MPORT_12_mask = 1'h1;
  assign bht_MPORT_12_en = reset;
  assign bht_MPORT_13_data = 6'h0;
  assign bht_MPORT_13_addr = 6'hc;
  assign bht_MPORT_13_mask = 1'h1;
  assign bht_MPORT_13_en = reset;
  assign bht_MPORT_14_data = 6'h0;
  assign bht_MPORT_14_addr = 6'hd;
  assign bht_MPORT_14_mask = 1'h1;
  assign bht_MPORT_14_en = reset;
  assign bht_MPORT_15_data = 6'h0;
  assign bht_MPORT_15_addr = 6'he;
  assign bht_MPORT_15_mask = 1'h1;
  assign bht_MPORT_15_en = reset;
  assign bht_MPORT_16_data = 6'h0;
  assign bht_MPORT_16_addr = 6'hf;
  assign bht_MPORT_16_mask = 1'h1;
  assign bht_MPORT_16_en = reset;
  assign bht_MPORT_17_data = 6'h0;
  assign bht_MPORT_17_addr = 6'h10;
  assign bht_MPORT_17_mask = 1'h1;
  assign bht_MPORT_17_en = reset;
  assign bht_MPORT_18_data = 6'h0;
  assign bht_MPORT_18_addr = 6'h11;
  assign bht_MPORT_18_mask = 1'h1;
  assign bht_MPORT_18_en = reset;
  assign bht_MPORT_19_data = 6'h0;
  assign bht_MPORT_19_addr = 6'h12;
  assign bht_MPORT_19_mask = 1'h1;
  assign bht_MPORT_19_en = reset;
  assign bht_MPORT_20_data = 6'h0;
  assign bht_MPORT_20_addr = 6'h13;
  assign bht_MPORT_20_mask = 1'h1;
  assign bht_MPORT_20_en = reset;
  assign bht_MPORT_21_data = 6'h0;
  assign bht_MPORT_21_addr = 6'h14;
  assign bht_MPORT_21_mask = 1'h1;
  assign bht_MPORT_21_en = reset;
  assign bht_MPORT_22_data = 6'h0;
  assign bht_MPORT_22_addr = 6'h15;
  assign bht_MPORT_22_mask = 1'h1;
  assign bht_MPORT_22_en = reset;
  assign bht_MPORT_23_data = 6'h0;
  assign bht_MPORT_23_addr = 6'h16;
  assign bht_MPORT_23_mask = 1'h1;
  assign bht_MPORT_23_en = reset;
  assign bht_MPORT_24_data = 6'h0;
  assign bht_MPORT_24_addr = 6'h17;
  assign bht_MPORT_24_mask = 1'h1;
  assign bht_MPORT_24_en = reset;
  assign bht_MPORT_25_data = 6'h0;
  assign bht_MPORT_25_addr = 6'h18;
  assign bht_MPORT_25_mask = 1'h1;
  assign bht_MPORT_25_en = reset;
  assign bht_MPORT_26_data = 6'h0;
  assign bht_MPORT_26_addr = 6'h19;
  assign bht_MPORT_26_mask = 1'h1;
  assign bht_MPORT_26_en = reset;
  assign bht_MPORT_27_data = 6'h0;
  assign bht_MPORT_27_addr = 6'h1a;
  assign bht_MPORT_27_mask = 1'h1;
  assign bht_MPORT_27_en = reset;
  assign bht_MPORT_28_data = 6'h0;
  assign bht_MPORT_28_addr = 6'h1b;
  assign bht_MPORT_28_mask = 1'h1;
  assign bht_MPORT_28_en = reset;
  assign bht_MPORT_29_data = 6'h0;
  assign bht_MPORT_29_addr = 6'h1c;
  assign bht_MPORT_29_mask = 1'h1;
  assign bht_MPORT_29_en = reset;
  assign bht_MPORT_30_data = 6'h0;
  assign bht_MPORT_30_addr = 6'h1d;
  assign bht_MPORT_30_mask = 1'h1;
  assign bht_MPORT_30_en = reset;
  assign bht_MPORT_31_data = 6'h0;
  assign bht_MPORT_31_addr = 6'h1e;
  assign bht_MPORT_31_mask = 1'h1;
  assign bht_MPORT_31_en = reset;
  assign bht_MPORT_32_data = 6'h0;
  assign bht_MPORT_32_addr = 6'h1f;
  assign bht_MPORT_32_mask = 1'h1;
  assign bht_MPORT_32_en = reset;
  assign bht_MPORT_33_data = 6'h0;
  assign bht_MPORT_33_addr = 6'h20;
  assign bht_MPORT_33_mask = 1'h1;
  assign bht_MPORT_33_en = reset;
  assign bht_MPORT_34_data = 6'h0;
  assign bht_MPORT_34_addr = 6'h21;
  assign bht_MPORT_34_mask = 1'h1;
  assign bht_MPORT_34_en = reset;
  assign bht_MPORT_35_data = 6'h0;
  assign bht_MPORT_35_addr = 6'h22;
  assign bht_MPORT_35_mask = 1'h1;
  assign bht_MPORT_35_en = reset;
  assign bht_MPORT_36_data = 6'h0;
  assign bht_MPORT_36_addr = 6'h23;
  assign bht_MPORT_36_mask = 1'h1;
  assign bht_MPORT_36_en = reset;
  assign bht_MPORT_37_data = 6'h0;
  assign bht_MPORT_37_addr = 6'h24;
  assign bht_MPORT_37_mask = 1'h1;
  assign bht_MPORT_37_en = reset;
  assign bht_MPORT_38_data = 6'h0;
  assign bht_MPORT_38_addr = 6'h25;
  assign bht_MPORT_38_mask = 1'h1;
  assign bht_MPORT_38_en = reset;
  assign bht_MPORT_39_data = 6'h0;
  assign bht_MPORT_39_addr = 6'h26;
  assign bht_MPORT_39_mask = 1'h1;
  assign bht_MPORT_39_en = reset;
  assign bht_MPORT_40_data = 6'h0;
  assign bht_MPORT_40_addr = 6'h27;
  assign bht_MPORT_40_mask = 1'h1;
  assign bht_MPORT_40_en = reset;
  assign bht_MPORT_41_data = 6'h0;
  assign bht_MPORT_41_addr = 6'h28;
  assign bht_MPORT_41_mask = 1'h1;
  assign bht_MPORT_41_en = reset;
  assign bht_MPORT_42_data = 6'h0;
  assign bht_MPORT_42_addr = 6'h29;
  assign bht_MPORT_42_mask = 1'h1;
  assign bht_MPORT_42_en = reset;
  assign bht_MPORT_43_data = 6'h0;
  assign bht_MPORT_43_addr = 6'h2a;
  assign bht_MPORT_43_mask = 1'h1;
  assign bht_MPORT_43_en = reset;
  assign bht_MPORT_44_data = 6'h0;
  assign bht_MPORT_44_addr = 6'h2b;
  assign bht_MPORT_44_mask = 1'h1;
  assign bht_MPORT_44_en = reset;
  assign bht_MPORT_45_data = 6'h0;
  assign bht_MPORT_45_addr = 6'h2c;
  assign bht_MPORT_45_mask = 1'h1;
  assign bht_MPORT_45_en = reset;
  assign bht_MPORT_46_data = 6'h0;
  assign bht_MPORT_46_addr = 6'h2d;
  assign bht_MPORT_46_mask = 1'h1;
  assign bht_MPORT_46_en = reset;
  assign bht_MPORT_47_data = 6'h0;
  assign bht_MPORT_47_addr = 6'h2e;
  assign bht_MPORT_47_mask = 1'h1;
  assign bht_MPORT_47_en = reset;
  assign bht_MPORT_48_data = 6'h0;
  assign bht_MPORT_48_addr = 6'h2f;
  assign bht_MPORT_48_mask = 1'h1;
  assign bht_MPORT_48_en = reset;
  assign bht_MPORT_49_data = 6'h0;
  assign bht_MPORT_49_addr = 6'h30;
  assign bht_MPORT_49_mask = 1'h1;
  assign bht_MPORT_49_en = reset;
  assign bht_MPORT_50_data = 6'h0;
  assign bht_MPORT_50_addr = 6'h31;
  assign bht_MPORT_50_mask = 1'h1;
  assign bht_MPORT_50_en = reset;
  assign bht_MPORT_51_data = 6'h0;
  assign bht_MPORT_51_addr = 6'h32;
  assign bht_MPORT_51_mask = 1'h1;
  assign bht_MPORT_51_en = reset;
  assign bht_MPORT_52_data = 6'h0;
  assign bht_MPORT_52_addr = 6'h33;
  assign bht_MPORT_52_mask = 1'h1;
  assign bht_MPORT_52_en = reset;
  assign bht_MPORT_53_data = 6'h0;
  assign bht_MPORT_53_addr = 6'h34;
  assign bht_MPORT_53_mask = 1'h1;
  assign bht_MPORT_53_en = reset;
  assign bht_MPORT_54_data = 6'h0;
  assign bht_MPORT_54_addr = 6'h35;
  assign bht_MPORT_54_mask = 1'h1;
  assign bht_MPORT_54_en = reset;
  assign bht_MPORT_55_data = 6'h0;
  assign bht_MPORT_55_addr = 6'h36;
  assign bht_MPORT_55_mask = 1'h1;
  assign bht_MPORT_55_en = reset;
  assign bht_MPORT_56_data = 6'h0;
  assign bht_MPORT_56_addr = 6'h37;
  assign bht_MPORT_56_mask = 1'h1;
  assign bht_MPORT_56_en = reset;
  assign bht_MPORT_57_data = 6'h0;
  assign bht_MPORT_57_addr = 6'h38;
  assign bht_MPORT_57_mask = 1'h1;
  assign bht_MPORT_57_en = reset;
  assign bht_MPORT_58_data = 6'h0;
  assign bht_MPORT_58_addr = 6'h39;
  assign bht_MPORT_58_mask = 1'h1;
  assign bht_MPORT_58_en = reset;
  assign bht_MPORT_59_data = 6'h0;
  assign bht_MPORT_59_addr = 6'h3a;
  assign bht_MPORT_59_mask = 1'h1;
  assign bht_MPORT_59_en = reset;
  assign bht_MPORT_60_data = 6'h0;
  assign bht_MPORT_60_addr = 6'h3b;
  assign bht_MPORT_60_mask = 1'h1;
  assign bht_MPORT_60_en = reset;
  assign bht_MPORT_61_data = 6'h0;
  assign bht_MPORT_61_addr = 6'h3c;
  assign bht_MPORT_61_mask = 1'h1;
  assign bht_MPORT_61_en = reset;
  assign bht_MPORT_62_data = 6'h0;
  assign bht_MPORT_62_addr = 6'h3d;
  assign bht_MPORT_62_mask = 1'h1;
  assign bht_MPORT_62_en = reset;
  assign bht_MPORT_63_data = 6'h0;
  assign bht_MPORT_63_addr = 6'h3e;
  assign bht_MPORT_63_mask = 1'h1;
  assign bht_MPORT_63_en = reset;
  assign bht_MPORT_64_data = 6'h0;
  assign bht_MPORT_64_addr = 6'h3f;
  assign bht_MPORT_64_mask = 1'h1;
  assign bht_MPORT_64_en = reset;
  assign io_pred_br_0 = pc_en_0 & pred_br_0; // @[BranchPredictor.scala 207:25]
  assign io_pred_br_1 = pc_en_1 & pred_br_1; // @[BranchPredictor.scala 207:25]
  assign io_pred_bpc = 2'h2 == _T_106 ? pred_bpc_1 : _T_110; // @[Mux.scala 80:57]
  assign io_pred_valid = REG_8; // @[BranchPredictor.scala 214:17]
  assign pht_clock = clock;
  assign pht_reset = reset;
  assign pht_io_rindex_0 = pc_0[10:8]; // @[BranchPredictor.scala 104:35]
  assign pht_io_rindex_1 = pc_1[10:8]; // @[BranchPredictor.scala 104:35]
  assign pht_io_raddr_0 = bht_bht_rdata_0_data ^ bht_raddr_0; // @[BranchPredictor.scala 103:58]
  assign pht_io_raddr_1 = bht_bht_rdata_1_data ^ bht_raddr_1; // @[BranchPredictor.scala 103:58]
  assign pht_io_windex = io_jmp_packet_inst_pc[10:8]; // @[BranchPredictor.scala 104:35]
  assign pht_io_waddr = bht_bht_wrdata_data ^ bht_waddr; // @[BranchPredictor.scala 103:58]
  assign pht_io_wen = io_jmp_packet_valid & ~io_jmp_packet_sys; // @[BranchPredictor.scala 62:43]
  assign pht_io_wjmp = io_jmp_packet_jmp; // @[BranchPredictor.scala 118:15]
  assign btb_clock = clock;
  assign btb_reset = reset;
  assign btb_io_raddr_0 = pc_0[5:2]; // @[BranchPredictor.scala 123:34]
  assign btb_io_raddr_1 = pc_1[5:2]; // @[BranchPredictor.scala 123:34]
  assign btb_io_ren_0 = pc_en_0; // @[BranchPredictor.scala 132:19]
  assign btb_io_ren_1 = pc_en_1; // @[BranchPredictor.scala 132:19]
  assign btb_io_rtag_0 = pc_0[31:6]; // @[BranchPredictor.scala 124:33]
  assign btb_io_rtag_1 = pc_1[31:6]; // @[BranchPredictor.scala 124:33]
  assign btb_io_waddr = io_jmp_packet_inst_pc[5:2]; // @[BranchPredictor.scala 123:34]
  assign btb_io_wen = jmp_packet_valid & io_jmp_packet_jmp; // @[BranchPredictor.scala 141:34]
  assign btb_io_wtag = io_jmp_packet_inst_pc[31:6]; // @[BranchPredictor.scala 124:33]
  assign btb_io_wtarget = io_jmp_packet_jmp_pc; // @[BranchPredictor.scala 143:18]
  always @(posedge clock) begin
    if (bht_MPORT_en & bht_MPORT_mask) begin
      bht[bht_MPORT_addr] <= bht_MPORT_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_1_en & bht_MPORT_1_mask) begin
      bht[bht_MPORT_1_addr] <= bht_MPORT_1_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_2_en & bht_MPORT_2_mask) begin
      bht[bht_MPORT_2_addr] <= bht_MPORT_2_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_3_en & bht_MPORT_3_mask) begin
      bht[bht_MPORT_3_addr] <= bht_MPORT_3_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_4_en & bht_MPORT_4_mask) begin
      bht[bht_MPORT_4_addr] <= bht_MPORT_4_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_5_en & bht_MPORT_5_mask) begin
      bht[bht_MPORT_5_addr] <= bht_MPORT_5_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_6_en & bht_MPORT_6_mask) begin
      bht[bht_MPORT_6_addr] <= bht_MPORT_6_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_7_en & bht_MPORT_7_mask) begin
      bht[bht_MPORT_7_addr] <= bht_MPORT_7_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_8_en & bht_MPORT_8_mask) begin
      bht[bht_MPORT_8_addr] <= bht_MPORT_8_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_9_en & bht_MPORT_9_mask) begin
      bht[bht_MPORT_9_addr] <= bht_MPORT_9_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_10_en & bht_MPORT_10_mask) begin
      bht[bht_MPORT_10_addr] <= bht_MPORT_10_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_11_en & bht_MPORT_11_mask) begin
      bht[bht_MPORT_11_addr] <= bht_MPORT_11_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_12_en & bht_MPORT_12_mask) begin
      bht[bht_MPORT_12_addr] <= bht_MPORT_12_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_13_en & bht_MPORT_13_mask) begin
      bht[bht_MPORT_13_addr] <= bht_MPORT_13_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_14_en & bht_MPORT_14_mask) begin
      bht[bht_MPORT_14_addr] <= bht_MPORT_14_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_15_en & bht_MPORT_15_mask) begin
      bht[bht_MPORT_15_addr] <= bht_MPORT_15_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_16_en & bht_MPORT_16_mask) begin
      bht[bht_MPORT_16_addr] <= bht_MPORT_16_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_17_en & bht_MPORT_17_mask) begin
      bht[bht_MPORT_17_addr] <= bht_MPORT_17_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_18_en & bht_MPORT_18_mask) begin
      bht[bht_MPORT_18_addr] <= bht_MPORT_18_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_19_en & bht_MPORT_19_mask) begin
      bht[bht_MPORT_19_addr] <= bht_MPORT_19_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_20_en & bht_MPORT_20_mask) begin
      bht[bht_MPORT_20_addr] <= bht_MPORT_20_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_21_en & bht_MPORT_21_mask) begin
      bht[bht_MPORT_21_addr] <= bht_MPORT_21_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_22_en & bht_MPORT_22_mask) begin
      bht[bht_MPORT_22_addr] <= bht_MPORT_22_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_23_en & bht_MPORT_23_mask) begin
      bht[bht_MPORT_23_addr] <= bht_MPORT_23_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_24_en & bht_MPORT_24_mask) begin
      bht[bht_MPORT_24_addr] <= bht_MPORT_24_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_25_en & bht_MPORT_25_mask) begin
      bht[bht_MPORT_25_addr] <= bht_MPORT_25_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_26_en & bht_MPORT_26_mask) begin
      bht[bht_MPORT_26_addr] <= bht_MPORT_26_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_27_en & bht_MPORT_27_mask) begin
      bht[bht_MPORT_27_addr] <= bht_MPORT_27_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_28_en & bht_MPORT_28_mask) begin
      bht[bht_MPORT_28_addr] <= bht_MPORT_28_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_29_en & bht_MPORT_29_mask) begin
      bht[bht_MPORT_29_addr] <= bht_MPORT_29_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_30_en & bht_MPORT_30_mask) begin
      bht[bht_MPORT_30_addr] <= bht_MPORT_30_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_31_en & bht_MPORT_31_mask) begin
      bht[bht_MPORT_31_addr] <= bht_MPORT_31_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_32_en & bht_MPORT_32_mask) begin
      bht[bht_MPORT_32_addr] <= bht_MPORT_32_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_33_en & bht_MPORT_33_mask) begin
      bht[bht_MPORT_33_addr] <= bht_MPORT_33_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_34_en & bht_MPORT_34_mask) begin
      bht[bht_MPORT_34_addr] <= bht_MPORT_34_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_35_en & bht_MPORT_35_mask) begin
      bht[bht_MPORT_35_addr] <= bht_MPORT_35_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_36_en & bht_MPORT_36_mask) begin
      bht[bht_MPORT_36_addr] <= bht_MPORT_36_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_37_en & bht_MPORT_37_mask) begin
      bht[bht_MPORT_37_addr] <= bht_MPORT_37_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_38_en & bht_MPORT_38_mask) begin
      bht[bht_MPORT_38_addr] <= bht_MPORT_38_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_39_en & bht_MPORT_39_mask) begin
      bht[bht_MPORT_39_addr] <= bht_MPORT_39_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_40_en & bht_MPORT_40_mask) begin
      bht[bht_MPORT_40_addr] <= bht_MPORT_40_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_41_en & bht_MPORT_41_mask) begin
      bht[bht_MPORT_41_addr] <= bht_MPORT_41_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_42_en & bht_MPORT_42_mask) begin
      bht[bht_MPORT_42_addr] <= bht_MPORT_42_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_43_en & bht_MPORT_43_mask) begin
      bht[bht_MPORT_43_addr] <= bht_MPORT_43_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_44_en & bht_MPORT_44_mask) begin
      bht[bht_MPORT_44_addr] <= bht_MPORT_44_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_45_en & bht_MPORT_45_mask) begin
      bht[bht_MPORT_45_addr] <= bht_MPORT_45_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_46_en & bht_MPORT_46_mask) begin
      bht[bht_MPORT_46_addr] <= bht_MPORT_46_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_47_en & bht_MPORT_47_mask) begin
      bht[bht_MPORT_47_addr] <= bht_MPORT_47_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_48_en & bht_MPORT_48_mask) begin
      bht[bht_MPORT_48_addr] <= bht_MPORT_48_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_49_en & bht_MPORT_49_mask) begin
      bht[bht_MPORT_49_addr] <= bht_MPORT_49_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_50_en & bht_MPORT_50_mask) begin
      bht[bht_MPORT_50_addr] <= bht_MPORT_50_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_51_en & bht_MPORT_51_mask) begin
      bht[bht_MPORT_51_addr] <= bht_MPORT_51_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_52_en & bht_MPORT_52_mask) begin
      bht[bht_MPORT_52_addr] <= bht_MPORT_52_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_53_en & bht_MPORT_53_mask) begin
      bht[bht_MPORT_53_addr] <= bht_MPORT_53_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_54_en & bht_MPORT_54_mask) begin
      bht[bht_MPORT_54_addr] <= bht_MPORT_54_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_55_en & bht_MPORT_55_mask) begin
      bht[bht_MPORT_55_addr] <= bht_MPORT_55_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_56_en & bht_MPORT_56_mask) begin
      bht[bht_MPORT_56_addr] <= bht_MPORT_56_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_57_en & bht_MPORT_57_mask) begin
      bht[bht_MPORT_57_addr] <= bht_MPORT_57_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_58_en & bht_MPORT_58_mask) begin
      bht[bht_MPORT_58_addr] <= bht_MPORT_58_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_59_en & bht_MPORT_59_mask) begin
      bht[bht_MPORT_59_addr] <= bht_MPORT_59_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_60_en & bht_MPORT_60_mask) begin
      bht[bht_MPORT_60_addr] <= bht_MPORT_60_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_61_en & bht_MPORT_61_mask) begin
      bht[bht_MPORT_61_addr] <= bht_MPORT_61_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_62_en & bht_MPORT_62_mask) begin
      bht[bht_MPORT_62_addr] <= bht_MPORT_62_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_63_en & bht_MPORT_63_mask) begin
      bht[bht_MPORT_63_addr] <= bht_MPORT_63_data; // @[BranchPredictor.scala 68:16]
    end
    if (bht_MPORT_64_en & bht_MPORT_64_mask) begin
      bht[bht_MPORT_64_addr] <= bht_MPORT_64_data; // @[BranchPredictor.scala 68:16]
    end
    if (reset) begin // @[BranchPredictor.scala 55:22]
      pc_en_0 <= 1'h0; // @[BranchPredictor.scala 55:22]
    end else begin
      pc_en_0 <= io_pc_en & ~io_pc[2]; // @[BranchPredictor.scala 56:12]
    end
    if (reset) begin // @[BranchPredictor.scala 55:22]
      pc_en_1 <= 1'h0; // @[BranchPredictor.scala 55:22]
    end else begin
      pc_en_1 <= io_pc_en; // @[BranchPredictor.scala 57:12]
    end
    REG_4 <= pc_base + 32'h8; // @[BranchPredictor.scala 52:21]
    REG_5 <= pc_base + 32'h8; // @[BranchPredictor.scala 52:21]
    REG_6 <= pc_base + 32'h8; // @[BranchPredictor.scala 52:21]
    REG_7 <= pc_base + 32'h8; // @[BranchPredictor.scala 52:21]
    REG_8 <= io_pc_en; // @[BranchPredictor.scala 214:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    bht[initvar] = _RAND_0[5:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  pc_en_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  pc_en_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  REG_4 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  REG_5 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  REG_6 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  REG_7 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  REG_8 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_InstFetch(
  input         clock,
  input         reset,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [31:0] io_imem_req_bits_addr,
  output [67:0] io_imem_req_bits_user,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input  [67:0] io_imem_resp_bits_user,
  input         io_jmp_packet_valid,
  input  [31:0] io_jmp_packet_inst_pc,
  input         io_jmp_packet_jmp,
  input  [31:0] io_jmp_packet_jmp_pc,
  input         io_jmp_packet_mis,
  input         io_jmp_packet_sys,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_vec_0_pc,
  output [31:0] io_out_bits_vec_0_inst,
  output        io_out_bits_vec_0_pred_br,
  output [31:0] io_out_bits_vec_0_pred_bpc,
  output        io_out_bits_vec_0_valid,
  output [31:0] io_out_bits_vec_1_pc,
  output [31:0] io_out_bits_vec_1_inst,
  output        io_out_bits_vec_1_pred_br,
  output [31:0] io_out_bits_vec_1_pred_bpc,
  output        io_out_bits_vec_1_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  bp_clock; // @[InstFetch.scala 38:18]
  wire  bp_reset; // @[InstFetch.scala 38:18]
  wire [31:0] bp_io_pc; // @[InstFetch.scala 38:18]
  wire  bp_io_pc_en; // @[InstFetch.scala 38:18]
  wire  bp_io_jmp_packet_valid; // @[InstFetch.scala 38:18]
  wire [31:0] bp_io_jmp_packet_inst_pc; // @[InstFetch.scala 38:18]
  wire  bp_io_jmp_packet_jmp; // @[InstFetch.scala 38:18]
  wire [31:0] bp_io_jmp_packet_jmp_pc; // @[InstFetch.scala 38:18]
  wire  bp_io_jmp_packet_mis; // @[InstFetch.scala 38:18]
  wire  bp_io_jmp_packet_sys; // @[InstFetch.scala 38:18]
  wire  bp_io_pred_br_0; // @[InstFetch.scala 38:18]
  wire  bp_io_pred_br_1; // @[InstFetch.scala 38:18]
  wire [31:0] bp_io_pred_bpc; // @[InstFetch.scala 38:18]
  wire  bp_io_pred_valid; // @[InstFetch.scala 38:18]
  reg  empty; // @[InstFetch.scala 17:22]
  wire  _T = io_imem_resp_ready & io_imem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_0 = _T | empty; // @[InstFetch.scala 18:22 19:11 17:22]
  wire  _T_1 = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _T_3 = io_jmp_packet_inst_pc + 32'h4; // @[InstFetch.scala 26:83]
  wire [31:0] mis_pc = io_jmp_packet_jmp ? io_jmp_packet_jmp_pc : _T_3; // @[InstFetch.scala 26:19]
  reg  reg_mis; // @[InstFetch.scala 28:24]
  wire  _T_9 = ~io_jmp_packet_mis; // @[InstFetch.scala 31:31]
  reg  REG; // @[InstFetch.scala 33:23]
  wire  _GEN_2 = REG ? 1'h0 : reg_mis; // @[InstFetch.scala 33:60 34:13 28:24]
  wire  _GEN_3 = _T & ~io_jmp_packet_mis ? 1'h0 : _GEN_2; // @[InstFetch.scala 31:37 32:13]
  wire  _GEN_4 = io_jmp_packet_mis & (~empty | _T_1) | _GEN_3; // @[InstFetch.scala 29:40 30:13]
  reg [31:0] pc; // @[InstFetch.scala 43:19]
  wire [31:0] pc_base = {pc[31:3],3'h0}; // @[Cat.scala 30:58]
  reg [1:0] pc_valid; // @[InstFetch.scala 45:25]
  wire [31:0] npc_s = pc_base + 32'h8; // @[InstFetch.scala 48:23]
  reg  REG_1; // @[InstFetch.scala 51:49]
  reg [31:0] r; // @[Reg.scala 27:20]
  wire [31:0] _GEN_5 = REG_1 ? bp_io_pred_bpc : r; // @[Reg.scala 28:19 27:20 28:23]
  wire [1:0] _T_19 = {bp_io_pred_br_1,bp_io_pred_br_0}; // @[Cat.scala 30:58]
  wire  _T_21 = bp_io_pred_valid & _T_9; // @[InstFetch.scala 52:91]
  wire [1:0] _T_23 = _T_21 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_24 = _T_19 & _T_23; // @[InstFetch.scala 52:64]
  reg  REG_2; // @[InstFetch.scala 52:117]
  wire [1:0] _T_25 = io_jmp_packet_mis ? 2'h0 : _T_24; // @[Utils.scala 68:20]
  wire  _T_27 = REG_2 | io_jmp_packet_mis; // @[Utils.scala 69:72]
  reg [1:0] r_1; // @[Reg.scala 27:20]
  wire [1:0] pred_br = REG_2 ? _T_25 : r_1; // @[Utils.scala 69:8]
  wire  _T_28 = |pred_br; // @[InstFetch.scala 56:42]
  wire [31:0] _T_29 = |pred_br ? _GEN_5 : npc_s; // @[InstFetch.scala 56:33]
  wire [31:0] npc = io_jmp_packet_mis ? mis_pc : _T_29; // @[InstFetch.scala 56:16]
  wire [1:0] _GEN_8 = _GEN_5[2] ? 2'h2 : 2'h3; // @[InstFetch.scala 63:29 64:17]
  wire  pc_update = io_jmp_packet_mis | _T_1; // @[InstFetch.scala 73:23]
  wire [63:0] lo = {npc,pc[31:3],3'h0}; // @[Cat.scala 30:58]
  wire [3:0] hi = {pred_br,pc_valid}; // @[Cat.scala 30:58]
  reg  REG_3; // @[InstFetch.scala 108:67]
  ysyx_210128_BranchPredictor bp ( // @[InstFetch.scala 38:18]
    .clock(bp_clock),
    .reset(bp_reset),
    .io_pc(bp_io_pc),
    .io_pc_en(bp_io_pc_en),
    .io_jmp_packet_valid(bp_io_jmp_packet_valid),
    .io_jmp_packet_inst_pc(bp_io_jmp_packet_inst_pc),
    .io_jmp_packet_jmp(bp_io_jmp_packet_jmp),
    .io_jmp_packet_jmp_pc(bp_io_jmp_packet_jmp_pc),
    .io_jmp_packet_mis(bp_io_jmp_packet_mis),
    .io_jmp_packet_sys(bp_io_jmp_packet_sys),
    .io_pred_br_0(bp_io_pred_br_0),
    .io_pred_br_1(bp_io_pred_br_1),
    .io_pred_bpc(bp_io_pred_bpc),
    .io_pred_valid(bp_io_pred_valid)
  );
  assign io_imem_req_valid = io_out_ready; // @[InstFetch.scala 90:18]
  assign io_imem_req_bits_addr = {pc[31:3],3'h0}; // @[Cat.scala 30:58]
  assign io_imem_req_bits_user = {hi,lo}; // @[Cat.scala 30:58]
  assign io_imem_resp_ready = io_out_ready | io_jmp_packet_mis; // @[InstFetch.scala 92:30]
  assign io_out_valid = io_imem_resp_valid & _T_9 & ~reg_mis & REG_3; // @[InstFetch.scala 108:57]
  assign io_out_bits_vec_0_pc = io_imem_resp_bits_user[31:0]; // @[InstFetch.scala 102:40]
  assign io_out_bits_vec_0_inst = io_imem_resp_bits_rdata[31:0]; // @[InstFetch.scala 103:41]
  assign io_out_bits_vec_0_pred_br = io_imem_resp_bits_user[66] & io_out_bits_vec_0_valid; // @[InstFetch.scala 104:45]
  assign io_out_bits_vec_0_pred_bpc = io_out_bits_vec_0_pred_br ? io_imem_resp_bits_user[63:32] : 32'h0; // @[InstFetch.scala 105:29]
  assign io_out_bits_vec_0_valid = io_imem_resp_bits_user[64]; // @[InstFetch.scala 106:40]
  assign io_out_bits_vec_1_pc = io_imem_resp_bits_user[31:0] + 32'h4; // @[InstFetch.scala 96:48]
  assign io_out_bits_vec_1_inst = io_imem_resp_bits_rdata[63:32]; // @[InstFetch.scala 97:41]
  assign io_out_bits_vec_1_pred_br = io_imem_resp_bits_user[67]; // @[InstFetch.scala 98:40]
  assign io_out_bits_vec_1_pred_bpc = io_out_bits_vec_1_pred_br ? io_imem_resp_bits_user[63:32] : 32'h0; // @[InstFetch.scala 99:29]
  assign io_out_bits_vec_1_valid = ~io_out_bits_vec_0_pred_br & io_imem_resp_bits_user[65]; // @[InstFetch.scala 100:46]
  assign bp_clock = clock;
  assign bp_reset = reset;
  assign bp_io_pc = io_jmp_packet_mis ? mis_pc : _T_29; // @[InstFetch.scala 56:16]
  assign bp_io_pc_en = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 40:37]
  assign bp_io_jmp_packet_valid = io_jmp_packet_valid; // @[InstFetch.scala 69:20]
  assign bp_io_jmp_packet_inst_pc = io_jmp_packet_inst_pc; // @[InstFetch.scala 69:20]
  assign bp_io_jmp_packet_jmp = io_jmp_packet_jmp; // @[InstFetch.scala 69:20]
  assign bp_io_jmp_packet_jmp_pc = io_jmp_packet_jmp_pc; // @[InstFetch.scala 69:20]
  assign bp_io_jmp_packet_mis = io_jmp_packet_mis; // @[InstFetch.scala 69:20]
  assign bp_io_jmp_packet_sys = io_jmp_packet_sys; // @[InstFetch.scala 69:20]
  always @(posedge clock) begin
    if (reset) begin // @[InstFetch.scala 17:22]
      empty <= 1'h0; // @[InstFetch.scala 17:22]
    end else if (_T_1) begin // @[InstFetch.scala 21:21]
      empty <= 1'h0; // @[InstFetch.scala 22:11]
    end else begin
      empty <= _GEN_0;
    end
    if (reset) begin // @[InstFetch.scala 28:24]
      reg_mis <= 1'h0; // @[InstFetch.scala 28:24]
    end else begin
      reg_mis <= _GEN_4;
    end
    REG <= _T & ~_T_1 & io_jmp_packet_mis; // @[InstFetch.scala 33:51]
    if (reset) begin // @[InstFetch.scala 43:19]
      pc <= 32'h30000000; // @[InstFetch.scala 43:19]
    end else if (pc_update) begin // @[InstFetch.scala 75:20]
      if (io_jmp_packet_mis) begin // @[InstFetch.scala 56:16]
        if (io_jmp_packet_jmp) begin // @[InstFetch.scala 26:19]
          pc <= io_jmp_packet_jmp_pc;
        end else begin
          pc <= _T_3;
        end
      end else if (|pred_br) begin // @[InstFetch.scala 56:33]
        pc <= _GEN_5;
      end else begin
        pc <= npc_s;
      end
    end
    if (reset) begin // @[InstFetch.scala 45:25]
      pc_valid <= 2'h3; // @[InstFetch.scala 45:25]
    end else if (pc_update) begin // @[InstFetch.scala 75:20]
      if (io_jmp_packet_mis) begin // @[InstFetch.scala 58:14]
        if (mis_pc[2]) begin // @[InstFetch.scala 59:30]
          pc_valid <= 2'h2; // @[InstFetch.scala 60:17]
        end else begin
          pc_valid <= 2'h3;
        end
      end else if (_T_28) begin // @[InstFetch.scala 62:29]
        pc_valid <= _GEN_8;
      end else begin
        pc_valid <= 2'h3;
      end
    end
    REG_1 <= io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 40:37]
    if (reset) begin // @[Reg.scala 27:20]
      r <= 32'h0; // @[Reg.scala 27:20]
    end else if (REG_1) begin // @[Reg.scala 28:19]
      r <= bp_io_pred_bpc; // @[Reg.scala 28:23]
    end
    REG_2 <= io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 40:37]
    if (reset) begin // @[Reg.scala 27:20]
      r_1 <= 2'h0; // @[Reg.scala 27:20]
    end else if (_T_27) begin // @[Reg.scala 28:19]
      if (io_jmp_packet_mis) begin // @[Utils.scala 68:20]
        r_1 <= 2'h0;
      end else begin
        r_1 <= _T_24;
      end
    end
    REG_3 <= ~io_jmp_packet_mis; // @[InstFetch.scala 108:68]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  empty = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_mis = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pc = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  pc_valid = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  REG_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  REG_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  r_1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  REG_3 = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_Sram(
  input          clock,
  input          io_en,
  input          io_wen,
  input  [5:0]   io_addr,
  input  [127:0] io_wdata,
  output [127:0] io_rdata
);
  wire  sram_CLK; // @[Sram.scala 35:20]
  wire  sram_CEN; // @[Sram.scala 35:20]
  wire  sram_WEN; // @[Sram.scala 35:20]
  wire [5:0] sram_A; // @[Sram.scala 35:20]
  wire [127:0] sram_D; // @[Sram.scala 35:20]
  wire [127:0] sram_Q; // @[Sram.scala 35:20]
  S011HD1P_X32Y2D128 sram ( // @[Sram.scala 35:20]
    .CLK(sram_CLK),
    .CEN(sram_CEN),
    .WEN(sram_WEN),
    .A(sram_A),
    .D(sram_D),
    .Q(sram_Q)
  );
  assign io_rdata = sram_Q; // @[Sram.scala 41:12]
  assign sram_CLK = clock; // @[Sram.scala 36:12]
  assign sram_CEN = ~io_en; // @[Sram.scala 37:15]
  assign sram_WEN = ~io_wen; // @[Sram.scala 38:15]
  assign sram_A = io_addr; // @[Sram.scala 39:10]
  assign sram_D = io_wdata; // @[Sram.scala 40:10]
endmodule
module ysyx_210128_Meta(
  input         clock,
  input         reset,
  input  [5:0]  io_idx,
  output [20:0] io_tag_r,
  input  [20:0] io_tag_w,
  input         io_tag_wen,
  output        io_dirty_r_async,
  input         io_dirty_w,
  input         io_dirty_wen,
  output        io_valid_r_async,
  input         io_invalidate
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] tags [0:63]; // @[Cache.scala 33:25]
//   wire  tags_MPORT_1_en; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_1_addr; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_1_data; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_2_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_2_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_2_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_2_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_3_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_3_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_3_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_3_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_4_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_4_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_4_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_4_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_5_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_5_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_5_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_5_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_6_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_6_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_6_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_6_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_7_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_7_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_7_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_7_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_8_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_8_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_8_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_8_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_9_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_9_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_9_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_9_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_10_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_10_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_10_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_10_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_11_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_11_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_11_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_11_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_12_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_12_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_12_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_12_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_13_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_13_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_13_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_13_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_14_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_14_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_14_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_14_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_15_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_15_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_15_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_15_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_16_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_16_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_16_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_16_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_17_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_17_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_17_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_17_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_18_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_18_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_18_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_18_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_19_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_19_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_19_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_19_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_20_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_20_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_20_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_20_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_21_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_21_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_21_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_21_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_22_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_22_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_22_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_22_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_23_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_23_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_23_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_23_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_24_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_24_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_24_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_24_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_25_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_25_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_25_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_25_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_26_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_26_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_26_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_26_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_27_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_27_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_27_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_27_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_28_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_28_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_28_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_28_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_29_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_29_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_29_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_29_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_30_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_30_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_30_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_30_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_31_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_31_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_31_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_31_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_32_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_32_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_32_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_32_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_33_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_33_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_33_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_33_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_34_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_34_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_34_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_34_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_35_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_35_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_35_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_35_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_36_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_36_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_36_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_36_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_37_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_37_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_37_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_37_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_38_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_38_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_38_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_38_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_39_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_39_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_39_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_39_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_40_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_40_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_40_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_40_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_41_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_41_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_41_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_41_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_42_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_42_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_42_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_42_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_43_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_43_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_43_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_43_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_44_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_44_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_44_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_44_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_45_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_45_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_45_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_45_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_46_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_46_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_46_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_46_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_47_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_47_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_47_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_47_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_48_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_48_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_48_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_48_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_49_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_49_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_49_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_49_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_50_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_50_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_50_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_50_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_51_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_51_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_51_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_51_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_52_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_52_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_52_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_52_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_53_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_53_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_53_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_53_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_54_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_54_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_54_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_54_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_55_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_55_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_55_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_55_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_56_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_56_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_56_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_56_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_57_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_57_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_57_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_57_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_58_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_58_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_58_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_58_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_59_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_59_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_59_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_59_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_60_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_60_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_60_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_60_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_61_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_61_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_61_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_61_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_62_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_62_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_62_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_62_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_63_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_63_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_63_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_63_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_64_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_64_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_64_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_64_en; // @[Cache.scala 33:25]
  wire [20:0] tags_MPORT_65_data; // @[Cache.scala 33:25]
  wire [5:0] tags_MPORT_65_addr; // @[Cache.scala 33:25]
  wire  tags_MPORT_65_mask; // @[Cache.scala 33:25]
  wire  tags_MPORT_65_en; // @[Cache.scala 33:25]
//   reg  tags_MPORT_1_en_pipe_0;
  reg [5:0] tags_MPORT_1_addr_pipe_0;
  reg  valid_0; // @[Cache.scala 35:22]
  reg  valid_1; // @[Cache.scala 35:22]
  reg  valid_2; // @[Cache.scala 35:22]
  reg  valid_3; // @[Cache.scala 35:22]
  reg  valid_4; // @[Cache.scala 35:22]
  reg  valid_5; // @[Cache.scala 35:22]
  reg  valid_6; // @[Cache.scala 35:22]
  reg  valid_7; // @[Cache.scala 35:22]
  reg  valid_8; // @[Cache.scala 35:22]
  reg  valid_9; // @[Cache.scala 35:22]
  reg  valid_10; // @[Cache.scala 35:22]
  reg  valid_11; // @[Cache.scala 35:22]
  reg  valid_12; // @[Cache.scala 35:22]
  reg  valid_13; // @[Cache.scala 35:22]
  reg  valid_14; // @[Cache.scala 35:22]
  reg  valid_15; // @[Cache.scala 35:22]
  reg  valid_16; // @[Cache.scala 35:22]
  reg  valid_17; // @[Cache.scala 35:22]
  reg  valid_18; // @[Cache.scala 35:22]
  reg  valid_19; // @[Cache.scala 35:22]
  reg  valid_20; // @[Cache.scala 35:22]
  reg  valid_21; // @[Cache.scala 35:22]
  reg  valid_22; // @[Cache.scala 35:22]
  reg  valid_23; // @[Cache.scala 35:22]
  reg  valid_24; // @[Cache.scala 35:22]
  reg  valid_25; // @[Cache.scala 35:22]
  reg  valid_26; // @[Cache.scala 35:22]
  reg  valid_27; // @[Cache.scala 35:22]
  reg  valid_28; // @[Cache.scala 35:22]
  reg  valid_29; // @[Cache.scala 35:22]
  reg  valid_30; // @[Cache.scala 35:22]
  reg  valid_31; // @[Cache.scala 35:22]
  reg  valid_32; // @[Cache.scala 35:22]
  reg  valid_33; // @[Cache.scala 35:22]
  reg  valid_34; // @[Cache.scala 35:22]
  reg  valid_35; // @[Cache.scala 35:22]
  reg  valid_36; // @[Cache.scala 35:22]
  reg  valid_37; // @[Cache.scala 35:22]
  reg  valid_38; // @[Cache.scala 35:22]
  reg  valid_39; // @[Cache.scala 35:22]
  reg  valid_40; // @[Cache.scala 35:22]
  reg  valid_41; // @[Cache.scala 35:22]
  reg  valid_42; // @[Cache.scala 35:22]
  reg  valid_43; // @[Cache.scala 35:22]
  reg  valid_44; // @[Cache.scala 35:22]
  reg  valid_45; // @[Cache.scala 35:22]
  reg  valid_46; // @[Cache.scala 35:22]
  reg  valid_47; // @[Cache.scala 35:22]
  reg  valid_48; // @[Cache.scala 35:22]
  reg  valid_49; // @[Cache.scala 35:22]
  reg  valid_50; // @[Cache.scala 35:22]
  reg  valid_51; // @[Cache.scala 35:22]
  reg  valid_52; // @[Cache.scala 35:22]
  reg  valid_53; // @[Cache.scala 35:22]
  reg  valid_54; // @[Cache.scala 35:22]
  reg  valid_55; // @[Cache.scala 35:22]
  reg  valid_56; // @[Cache.scala 35:22]
  reg  valid_57; // @[Cache.scala 35:22]
  reg  valid_58; // @[Cache.scala 35:22]
  reg  valid_59; // @[Cache.scala 35:22]
  reg  valid_60; // @[Cache.scala 35:22]
  reg  valid_61; // @[Cache.scala 35:22]
  reg  valid_62; // @[Cache.scala 35:22]
  reg  valid_63; // @[Cache.scala 35:22]
  reg  dirty_0; // @[Cache.scala 39:22]
  reg  dirty_1; // @[Cache.scala 39:22]
  reg  dirty_2; // @[Cache.scala 39:22]
  reg  dirty_3; // @[Cache.scala 39:22]
  reg  dirty_4; // @[Cache.scala 39:22]
  reg  dirty_5; // @[Cache.scala 39:22]
  reg  dirty_6; // @[Cache.scala 39:22]
  reg  dirty_7; // @[Cache.scala 39:22]
  reg  dirty_8; // @[Cache.scala 39:22]
  reg  dirty_9; // @[Cache.scala 39:22]
  reg  dirty_10; // @[Cache.scala 39:22]
  reg  dirty_11; // @[Cache.scala 39:22]
  reg  dirty_12; // @[Cache.scala 39:22]
  reg  dirty_13; // @[Cache.scala 39:22]
  reg  dirty_14; // @[Cache.scala 39:22]
  reg  dirty_15; // @[Cache.scala 39:22]
  reg  dirty_16; // @[Cache.scala 39:22]
  reg  dirty_17; // @[Cache.scala 39:22]
  reg  dirty_18; // @[Cache.scala 39:22]
  reg  dirty_19; // @[Cache.scala 39:22]
  reg  dirty_20; // @[Cache.scala 39:22]
  reg  dirty_21; // @[Cache.scala 39:22]
  reg  dirty_22; // @[Cache.scala 39:22]
  reg  dirty_23; // @[Cache.scala 39:22]
  reg  dirty_24; // @[Cache.scala 39:22]
  reg  dirty_25; // @[Cache.scala 39:22]
  reg  dirty_26; // @[Cache.scala 39:22]
  reg  dirty_27; // @[Cache.scala 39:22]
  reg  dirty_28; // @[Cache.scala 39:22]
  reg  dirty_29; // @[Cache.scala 39:22]
  reg  dirty_30; // @[Cache.scala 39:22]
  reg  dirty_31; // @[Cache.scala 39:22]
  reg  dirty_32; // @[Cache.scala 39:22]
  reg  dirty_33; // @[Cache.scala 39:22]
  reg  dirty_34; // @[Cache.scala 39:22]
  reg  dirty_35; // @[Cache.scala 39:22]
  reg  dirty_36; // @[Cache.scala 39:22]
  reg  dirty_37; // @[Cache.scala 39:22]
  reg  dirty_38; // @[Cache.scala 39:22]
  reg  dirty_39; // @[Cache.scala 39:22]
  reg  dirty_40; // @[Cache.scala 39:22]
  reg  dirty_41; // @[Cache.scala 39:22]
  reg  dirty_42; // @[Cache.scala 39:22]
  reg  dirty_43; // @[Cache.scala 39:22]
  reg  dirty_44; // @[Cache.scala 39:22]
  reg  dirty_45; // @[Cache.scala 39:22]
  reg  dirty_46; // @[Cache.scala 39:22]
  reg  dirty_47; // @[Cache.scala 39:22]
  reg  dirty_48; // @[Cache.scala 39:22]
  reg  dirty_49; // @[Cache.scala 39:22]
  reg  dirty_50; // @[Cache.scala 39:22]
  reg  dirty_51; // @[Cache.scala 39:22]
  reg  dirty_52; // @[Cache.scala 39:22]
  reg  dirty_53; // @[Cache.scala 39:22]
  reg  dirty_54; // @[Cache.scala 39:22]
  reg  dirty_55; // @[Cache.scala 39:22]
  reg  dirty_56; // @[Cache.scala 39:22]
  reg  dirty_57; // @[Cache.scala 39:22]
  reg  dirty_58; // @[Cache.scala 39:22]
  reg  dirty_59; // @[Cache.scala 39:22]
  reg  dirty_60; // @[Cache.scala 39:22]
  reg  dirty_61; // @[Cache.scala 39:22]
  reg  dirty_62; // @[Cache.scala 39:22]
  reg  dirty_63; // @[Cache.scala 39:22]
  wire  _GEN_0 = 6'h0 == io_idx | valid_0; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_1 = 6'h1 == io_idx | valid_1; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_2 = 6'h2 == io_idx | valid_2; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_3 = 6'h3 == io_idx | valid_3; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_4 = 6'h4 == io_idx | valid_4; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_5 = 6'h5 == io_idx | valid_5; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_6 = 6'h6 == io_idx | valid_6; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_7 = 6'h7 == io_idx | valid_7; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_8 = 6'h8 == io_idx | valid_8; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_9 = 6'h9 == io_idx | valid_9; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_10 = 6'ha == io_idx | valid_10; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_11 = 6'hb == io_idx | valid_11; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_12 = 6'hc == io_idx | valid_12; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_13 = 6'hd == io_idx | valid_13; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_14 = 6'he == io_idx | valid_14; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_15 = 6'hf == io_idx | valid_15; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_16 = 6'h10 == io_idx | valid_16; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_17 = 6'h11 == io_idx | valid_17; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_18 = 6'h12 == io_idx | valid_18; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_19 = 6'h13 == io_idx | valid_19; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_20 = 6'h14 == io_idx | valid_20; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_21 = 6'h15 == io_idx | valid_21; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_22 = 6'h16 == io_idx | valid_22; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_23 = 6'h17 == io_idx | valid_23; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_24 = 6'h18 == io_idx | valid_24; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_25 = 6'h19 == io_idx | valid_25; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_26 = 6'h1a == io_idx | valid_26; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_27 = 6'h1b == io_idx | valid_27; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_28 = 6'h1c == io_idx | valid_28; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_29 = 6'h1d == io_idx | valid_29; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_30 = 6'h1e == io_idx | valid_30; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_31 = 6'h1f == io_idx | valid_31; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_32 = 6'h20 == io_idx | valid_32; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_33 = 6'h21 == io_idx | valid_33; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_34 = 6'h22 == io_idx | valid_34; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_35 = 6'h23 == io_idx | valid_35; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_36 = 6'h24 == io_idx | valid_36; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_37 = 6'h25 == io_idx | valid_37; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_38 = 6'h26 == io_idx | valid_38; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_39 = 6'h27 == io_idx | valid_39; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_40 = 6'h28 == io_idx | valid_40; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_41 = 6'h29 == io_idx | valid_41; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_42 = 6'h2a == io_idx | valid_42; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_43 = 6'h2b == io_idx | valid_43; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_44 = 6'h2c == io_idx | valid_44; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_45 = 6'h2d == io_idx | valid_45; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_46 = 6'h2e == io_idx | valid_46; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_47 = 6'h2f == io_idx | valid_47; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_48 = 6'h30 == io_idx | valid_48; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_49 = 6'h31 == io_idx | valid_49; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_50 = 6'h32 == io_idx | valid_50; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_51 = 6'h33 == io_idx | valid_51; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_52 = 6'h34 == io_idx | valid_52; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_53 = 6'h35 == io_idx | valid_53; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_54 = 6'h36 == io_idx | valid_54; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_55 = 6'h37 == io_idx | valid_55; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_56 = 6'h38 == io_idx | valid_56; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_57 = 6'h39 == io_idx | valid_57; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_58 = 6'h3a == io_idx | valid_58; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_59 = 6'h3b == io_idx | valid_59; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_60 = 6'h3c == io_idx | valid_60; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_61 = 6'h3d == io_idx | valid_61; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_62 = 6'h3e == io_idx | valid_62; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_63 = 6'h3f == io_idx | valid_63; // @[Cache.scala 46:{16,16} 35:22]
  wire  _GEN_138 = 6'h1 == io_idx ? dirty_1 : dirty_0; // @[Cache.scala 51:{20,20}]
  wire  _GEN_139 = 6'h2 == io_idx ? dirty_2 : _GEN_138; // @[Cache.scala 51:{20,20}]
  wire  _GEN_140 = 6'h3 == io_idx ? dirty_3 : _GEN_139; // @[Cache.scala 51:{20,20}]
  wire  _GEN_141 = 6'h4 == io_idx ? dirty_4 : _GEN_140; // @[Cache.scala 51:{20,20}]
  wire  _GEN_142 = 6'h5 == io_idx ? dirty_5 : _GEN_141; // @[Cache.scala 51:{20,20}]
  wire  _GEN_143 = 6'h6 == io_idx ? dirty_6 : _GEN_142; // @[Cache.scala 51:{20,20}]
  wire  _GEN_144 = 6'h7 == io_idx ? dirty_7 : _GEN_143; // @[Cache.scala 51:{20,20}]
  wire  _GEN_145 = 6'h8 == io_idx ? dirty_8 : _GEN_144; // @[Cache.scala 51:{20,20}]
  wire  _GEN_146 = 6'h9 == io_idx ? dirty_9 : _GEN_145; // @[Cache.scala 51:{20,20}]
  wire  _GEN_147 = 6'ha == io_idx ? dirty_10 : _GEN_146; // @[Cache.scala 51:{20,20}]
  wire  _GEN_148 = 6'hb == io_idx ? dirty_11 : _GEN_147; // @[Cache.scala 51:{20,20}]
  wire  _GEN_149 = 6'hc == io_idx ? dirty_12 : _GEN_148; // @[Cache.scala 51:{20,20}]
  wire  _GEN_150 = 6'hd == io_idx ? dirty_13 : _GEN_149; // @[Cache.scala 51:{20,20}]
  wire  _GEN_151 = 6'he == io_idx ? dirty_14 : _GEN_150; // @[Cache.scala 51:{20,20}]
  wire  _GEN_152 = 6'hf == io_idx ? dirty_15 : _GEN_151; // @[Cache.scala 51:{20,20}]
  wire  _GEN_153 = 6'h10 == io_idx ? dirty_16 : _GEN_152; // @[Cache.scala 51:{20,20}]
  wire  _GEN_154 = 6'h11 == io_idx ? dirty_17 : _GEN_153; // @[Cache.scala 51:{20,20}]
  wire  _GEN_155 = 6'h12 == io_idx ? dirty_18 : _GEN_154; // @[Cache.scala 51:{20,20}]
  wire  _GEN_156 = 6'h13 == io_idx ? dirty_19 : _GEN_155; // @[Cache.scala 51:{20,20}]
  wire  _GEN_157 = 6'h14 == io_idx ? dirty_20 : _GEN_156; // @[Cache.scala 51:{20,20}]
  wire  _GEN_158 = 6'h15 == io_idx ? dirty_21 : _GEN_157; // @[Cache.scala 51:{20,20}]
  wire  _GEN_159 = 6'h16 == io_idx ? dirty_22 : _GEN_158; // @[Cache.scala 51:{20,20}]
  wire  _GEN_160 = 6'h17 == io_idx ? dirty_23 : _GEN_159; // @[Cache.scala 51:{20,20}]
  wire  _GEN_161 = 6'h18 == io_idx ? dirty_24 : _GEN_160; // @[Cache.scala 51:{20,20}]
  wire  _GEN_162 = 6'h19 == io_idx ? dirty_25 : _GEN_161; // @[Cache.scala 51:{20,20}]
  wire  _GEN_163 = 6'h1a == io_idx ? dirty_26 : _GEN_162; // @[Cache.scala 51:{20,20}]
  wire  _GEN_164 = 6'h1b == io_idx ? dirty_27 : _GEN_163; // @[Cache.scala 51:{20,20}]
  wire  _GEN_165 = 6'h1c == io_idx ? dirty_28 : _GEN_164; // @[Cache.scala 51:{20,20}]
  wire  _GEN_166 = 6'h1d == io_idx ? dirty_29 : _GEN_165; // @[Cache.scala 51:{20,20}]
  wire  _GEN_167 = 6'h1e == io_idx ? dirty_30 : _GEN_166; // @[Cache.scala 51:{20,20}]
  wire  _GEN_168 = 6'h1f == io_idx ? dirty_31 : _GEN_167; // @[Cache.scala 51:{20,20}]
  wire  _GEN_169 = 6'h20 == io_idx ? dirty_32 : _GEN_168; // @[Cache.scala 51:{20,20}]
  wire  _GEN_170 = 6'h21 == io_idx ? dirty_33 : _GEN_169; // @[Cache.scala 51:{20,20}]
  wire  _GEN_171 = 6'h22 == io_idx ? dirty_34 : _GEN_170; // @[Cache.scala 51:{20,20}]
  wire  _GEN_172 = 6'h23 == io_idx ? dirty_35 : _GEN_171; // @[Cache.scala 51:{20,20}]
  wire  _GEN_173 = 6'h24 == io_idx ? dirty_36 : _GEN_172; // @[Cache.scala 51:{20,20}]
  wire  _GEN_174 = 6'h25 == io_idx ? dirty_37 : _GEN_173; // @[Cache.scala 51:{20,20}]
  wire  _GEN_175 = 6'h26 == io_idx ? dirty_38 : _GEN_174; // @[Cache.scala 51:{20,20}]
  wire  _GEN_176 = 6'h27 == io_idx ? dirty_39 : _GEN_175; // @[Cache.scala 51:{20,20}]
  wire  _GEN_177 = 6'h28 == io_idx ? dirty_40 : _GEN_176; // @[Cache.scala 51:{20,20}]
  wire  _GEN_178 = 6'h29 == io_idx ? dirty_41 : _GEN_177; // @[Cache.scala 51:{20,20}]
  wire  _GEN_179 = 6'h2a == io_idx ? dirty_42 : _GEN_178; // @[Cache.scala 51:{20,20}]
  wire  _GEN_180 = 6'h2b == io_idx ? dirty_43 : _GEN_179; // @[Cache.scala 51:{20,20}]
  wire  _GEN_181 = 6'h2c == io_idx ? dirty_44 : _GEN_180; // @[Cache.scala 51:{20,20}]
  wire  _GEN_182 = 6'h2d == io_idx ? dirty_45 : _GEN_181; // @[Cache.scala 51:{20,20}]
  wire  _GEN_183 = 6'h2e == io_idx ? dirty_46 : _GEN_182; // @[Cache.scala 51:{20,20}]
  wire  _GEN_184 = 6'h2f == io_idx ? dirty_47 : _GEN_183; // @[Cache.scala 51:{20,20}]
  wire  _GEN_185 = 6'h30 == io_idx ? dirty_48 : _GEN_184; // @[Cache.scala 51:{20,20}]
  wire  _GEN_186 = 6'h31 == io_idx ? dirty_49 : _GEN_185; // @[Cache.scala 51:{20,20}]
  wire  _GEN_187 = 6'h32 == io_idx ? dirty_50 : _GEN_186; // @[Cache.scala 51:{20,20}]
  wire  _GEN_188 = 6'h33 == io_idx ? dirty_51 : _GEN_187; // @[Cache.scala 51:{20,20}]
  wire  _GEN_189 = 6'h34 == io_idx ? dirty_52 : _GEN_188; // @[Cache.scala 51:{20,20}]
  wire  _GEN_190 = 6'h35 == io_idx ? dirty_53 : _GEN_189; // @[Cache.scala 51:{20,20}]
  wire  _GEN_191 = 6'h36 == io_idx ? dirty_54 : _GEN_190; // @[Cache.scala 51:{20,20}]
  wire  _GEN_192 = 6'h37 == io_idx ? dirty_55 : _GEN_191; // @[Cache.scala 51:{20,20}]
  wire  _GEN_193 = 6'h38 == io_idx ? dirty_56 : _GEN_192; // @[Cache.scala 51:{20,20}]
  wire  _GEN_194 = 6'h39 == io_idx ? dirty_57 : _GEN_193; // @[Cache.scala 51:{20,20}]
  wire  _GEN_195 = 6'h3a == io_idx ? dirty_58 : _GEN_194; // @[Cache.scala 51:{20,20}]
  wire  _GEN_196 = 6'h3b == io_idx ? dirty_59 : _GEN_195; // @[Cache.scala 51:{20,20}]
  wire  _GEN_197 = 6'h3c == io_idx ? dirty_60 : _GEN_196; // @[Cache.scala 51:{20,20}]
  wire  _GEN_198 = 6'h3d == io_idx ? dirty_61 : _GEN_197; // @[Cache.scala 51:{20,20}]
  wire  _GEN_199 = 6'h3e == io_idx ? dirty_62 : _GEN_198; // @[Cache.scala 51:{20,20}]
  wire  _GEN_202 = 6'h1 == io_idx ? valid_1 : valid_0; // @[Cache.scala 52:{20,20}]
  wire  _GEN_203 = 6'h2 == io_idx ? valid_2 : _GEN_202; // @[Cache.scala 52:{20,20}]
  wire  _GEN_204 = 6'h3 == io_idx ? valid_3 : _GEN_203; // @[Cache.scala 52:{20,20}]
  wire  _GEN_205 = 6'h4 == io_idx ? valid_4 : _GEN_204; // @[Cache.scala 52:{20,20}]
  wire  _GEN_206 = 6'h5 == io_idx ? valid_5 : _GEN_205; // @[Cache.scala 52:{20,20}]
  wire  _GEN_207 = 6'h6 == io_idx ? valid_6 : _GEN_206; // @[Cache.scala 52:{20,20}]
  wire  _GEN_208 = 6'h7 == io_idx ? valid_7 : _GEN_207; // @[Cache.scala 52:{20,20}]
  wire  _GEN_209 = 6'h8 == io_idx ? valid_8 : _GEN_208; // @[Cache.scala 52:{20,20}]
  wire  _GEN_210 = 6'h9 == io_idx ? valid_9 : _GEN_209; // @[Cache.scala 52:{20,20}]
  wire  _GEN_211 = 6'ha == io_idx ? valid_10 : _GEN_210; // @[Cache.scala 52:{20,20}]
  wire  _GEN_212 = 6'hb == io_idx ? valid_11 : _GEN_211; // @[Cache.scala 52:{20,20}]
  wire  _GEN_213 = 6'hc == io_idx ? valid_12 : _GEN_212; // @[Cache.scala 52:{20,20}]
  wire  _GEN_214 = 6'hd == io_idx ? valid_13 : _GEN_213; // @[Cache.scala 52:{20,20}]
  wire  _GEN_215 = 6'he == io_idx ? valid_14 : _GEN_214; // @[Cache.scala 52:{20,20}]
  wire  _GEN_216 = 6'hf == io_idx ? valid_15 : _GEN_215; // @[Cache.scala 52:{20,20}]
  wire  _GEN_217 = 6'h10 == io_idx ? valid_16 : _GEN_216; // @[Cache.scala 52:{20,20}]
  wire  _GEN_218 = 6'h11 == io_idx ? valid_17 : _GEN_217; // @[Cache.scala 52:{20,20}]
  wire  _GEN_219 = 6'h12 == io_idx ? valid_18 : _GEN_218; // @[Cache.scala 52:{20,20}]
  wire  _GEN_220 = 6'h13 == io_idx ? valid_19 : _GEN_219; // @[Cache.scala 52:{20,20}]
  wire  _GEN_221 = 6'h14 == io_idx ? valid_20 : _GEN_220; // @[Cache.scala 52:{20,20}]
  wire  _GEN_222 = 6'h15 == io_idx ? valid_21 : _GEN_221; // @[Cache.scala 52:{20,20}]
  wire  _GEN_223 = 6'h16 == io_idx ? valid_22 : _GEN_222; // @[Cache.scala 52:{20,20}]
  wire  _GEN_224 = 6'h17 == io_idx ? valid_23 : _GEN_223; // @[Cache.scala 52:{20,20}]
  wire  _GEN_225 = 6'h18 == io_idx ? valid_24 : _GEN_224; // @[Cache.scala 52:{20,20}]
  wire  _GEN_226 = 6'h19 == io_idx ? valid_25 : _GEN_225; // @[Cache.scala 52:{20,20}]
  wire  _GEN_227 = 6'h1a == io_idx ? valid_26 : _GEN_226; // @[Cache.scala 52:{20,20}]
  wire  _GEN_228 = 6'h1b == io_idx ? valid_27 : _GEN_227; // @[Cache.scala 52:{20,20}]
  wire  _GEN_229 = 6'h1c == io_idx ? valid_28 : _GEN_228; // @[Cache.scala 52:{20,20}]
  wire  _GEN_230 = 6'h1d == io_idx ? valid_29 : _GEN_229; // @[Cache.scala 52:{20,20}]
  wire  _GEN_231 = 6'h1e == io_idx ? valid_30 : _GEN_230; // @[Cache.scala 52:{20,20}]
  wire  _GEN_232 = 6'h1f == io_idx ? valid_31 : _GEN_231; // @[Cache.scala 52:{20,20}]
  wire  _GEN_233 = 6'h20 == io_idx ? valid_32 : _GEN_232; // @[Cache.scala 52:{20,20}]
  wire  _GEN_234 = 6'h21 == io_idx ? valid_33 : _GEN_233; // @[Cache.scala 52:{20,20}]
  wire  _GEN_235 = 6'h22 == io_idx ? valid_34 : _GEN_234; // @[Cache.scala 52:{20,20}]
  wire  _GEN_236 = 6'h23 == io_idx ? valid_35 : _GEN_235; // @[Cache.scala 52:{20,20}]
  wire  _GEN_237 = 6'h24 == io_idx ? valid_36 : _GEN_236; // @[Cache.scala 52:{20,20}]
  wire  _GEN_238 = 6'h25 == io_idx ? valid_37 : _GEN_237; // @[Cache.scala 52:{20,20}]
  wire  _GEN_239 = 6'h26 == io_idx ? valid_38 : _GEN_238; // @[Cache.scala 52:{20,20}]
  wire  _GEN_240 = 6'h27 == io_idx ? valid_39 : _GEN_239; // @[Cache.scala 52:{20,20}]
  wire  _GEN_241 = 6'h28 == io_idx ? valid_40 : _GEN_240; // @[Cache.scala 52:{20,20}]
  wire  _GEN_242 = 6'h29 == io_idx ? valid_41 : _GEN_241; // @[Cache.scala 52:{20,20}]
  wire  _GEN_243 = 6'h2a == io_idx ? valid_42 : _GEN_242; // @[Cache.scala 52:{20,20}]
  wire  _GEN_244 = 6'h2b == io_idx ? valid_43 : _GEN_243; // @[Cache.scala 52:{20,20}]
  wire  _GEN_245 = 6'h2c == io_idx ? valid_44 : _GEN_244; // @[Cache.scala 52:{20,20}]
  wire  _GEN_246 = 6'h2d == io_idx ? valid_45 : _GEN_245; // @[Cache.scala 52:{20,20}]
  wire  _GEN_247 = 6'h2e == io_idx ? valid_46 : _GEN_246; // @[Cache.scala 52:{20,20}]
  wire  _GEN_248 = 6'h2f == io_idx ? valid_47 : _GEN_247; // @[Cache.scala 52:{20,20}]
  wire  _GEN_249 = 6'h30 == io_idx ? valid_48 : _GEN_248; // @[Cache.scala 52:{20,20}]
  wire  _GEN_250 = 6'h31 == io_idx ? valid_49 : _GEN_249; // @[Cache.scala 52:{20,20}]
  wire  _GEN_251 = 6'h32 == io_idx ? valid_50 : _GEN_250; // @[Cache.scala 52:{20,20}]
  wire  _GEN_252 = 6'h33 == io_idx ? valid_51 : _GEN_251; // @[Cache.scala 52:{20,20}]
  wire  _GEN_253 = 6'h34 == io_idx ? valid_52 : _GEN_252; // @[Cache.scala 52:{20,20}]
  wire  _GEN_254 = 6'h35 == io_idx ? valid_53 : _GEN_253; // @[Cache.scala 52:{20,20}]
  wire  _GEN_255 = 6'h36 == io_idx ? valid_54 : _GEN_254; // @[Cache.scala 52:{20,20}]
  wire  _GEN_256 = 6'h37 == io_idx ? valid_55 : _GEN_255; // @[Cache.scala 52:{20,20}]
  wire  _GEN_257 = 6'h38 == io_idx ? valid_56 : _GEN_256; // @[Cache.scala 52:{20,20}]
  wire  _GEN_258 = 6'h39 == io_idx ? valid_57 : _GEN_257; // @[Cache.scala 52:{20,20}]
  wire  _GEN_259 = 6'h3a == io_idx ? valid_58 : _GEN_258; // @[Cache.scala 52:{20,20}]
  wire  _GEN_260 = 6'h3b == io_idx ? valid_59 : _GEN_259; // @[Cache.scala 52:{20,20}]
  wire  _GEN_261 = 6'h3c == io_idx ? valid_60 : _GEN_260; // @[Cache.scala 52:{20,20}]
  wire  _GEN_262 = 6'h3d == io_idx ? valid_61 : _GEN_261; // @[Cache.scala 52:{20,20}]
  wire  _GEN_263 = 6'h3e == io_idx ? valid_62 : _GEN_262; // @[Cache.scala 52:{20,20}]
//   assign tags_MPORT_1_en = tags_MPORT_1_en_pipe_0;
  assign tags_MPORT_1_addr = tags_MPORT_1_addr_pipe_0;
  assign tags_MPORT_1_data = tags[tags_MPORT_1_addr]; // @[Cache.scala 33:25]
  assign tags_MPORT_data = io_tag_w;
  assign tags_MPORT_addr = io_idx;
  assign tags_MPORT_mask = 1'h1;
  assign tags_MPORT_en = io_tag_wen;
  assign tags_MPORT_2_data = 21'h0;
  assign tags_MPORT_2_addr = 6'h0;
  assign tags_MPORT_2_mask = 1'h1;
  assign tags_MPORT_2_en = reset;
  assign tags_MPORT_3_data = 21'h0;
  assign tags_MPORT_3_addr = 6'h1;
  assign tags_MPORT_3_mask = 1'h1;
  assign tags_MPORT_3_en = reset;
  assign tags_MPORT_4_data = 21'h0;
  assign tags_MPORT_4_addr = 6'h2;
  assign tags_MPORT_4_mask = 1'h1;
  assign tags_MPORT_4_en = reset;
  assign tags_MPORT_5_data = 21'h0;
  assign tags_MPORT_5_addr = 6'h3;
  assign tags_MPORT_5_mask = 1'h1;
  assign tags_MPORT_5_en = reset;
  assign tags_MPORT_6_data = 21'h0;
  assign tags_MPORT_6_addr = 6'h4;
  assign tags_MPORT_6_mask = 1'h1;
  assign tags_MPORT_6_en = reset;
  assign tags_MPORT_7_data = 21'h0;
  assign tags_MPORT_7_addr = 6'h5;
  assign tags_MPORT_7_mask = 1'h1;
  assign tags_MPORT_7_en = reset;
  assign tags_MPORT_8_data = 21'h0;
  assign tags_MPORT_8_addr = 6'h6;
  assign tags_MPORT_8_mask = 1'h1;
  assign tags_MPORT_8_en = reset;
  assign tags_MPORT_9_data = 21'h0;
  assign tags_MPORT_9_addr = 6'h7;
  assign tags_MPORT_9_mask = 1'h1;
  assign tags_MPORT_9_en = reset;
  assign tags_MPORT_10_data = 21'h0;
  assign tags_MPORT_10_addr = 6'h8;
  assign tags_MPORT_10_mask = 1'h1;
  assign tags_MPORT_10_en = reset;
  assign tags_MPORT_11_data = 21'h0;
  assign tags_MPORT_11_addr = 6'h9;
  assign tags_MPORT_11_mask = 1'h1;
  assign tags_MPORT_11_en = reset;
  assign tags_MPORT_12_data = 21'h0;
  assign tags_MPORT_12_addr = 6'ha;
  assign tags_MPORT_12_mask = 1'h1;
  assign tags_MPORT_12_en = reset;
  assign tags_MPORT_13_data = 21'h0;
  assign tags_MPORT_13_addr = 6'hb;
  assign tags_MPORT_13_mask = 1'h1;
  assign tags_MPORT_13_en = reset;
  assign tags_MPORT_14_data = 21'h0;
  assign tags_MPORT_14_addr = 6'hc;
  assign tags_MPORT_14_mask = 1'h1;
  assign tags_MPORT_14_en = reset;
  assign tags_MPORT_15_data = 21'h0;
  assign tags_MPORT_15_addr = 6'hd;
  assign tags_MPORT_15_mask = 1'h1;
  assign tags_MPORT_15_en = reset;
  assign tags_MPORT_16_data = 21'h0;
  assign tags_MPORT_16_addr = 6'he;
  assign tags_MPORT_16_mask = 1'h1;
  assign tags_MPORT_16_en = reset;
  assign tags_MPORT_17_data = 21'h0;
  assign tags_MPORT_17_addr = 6'hf;
  assign tags_MPORT_17_mask = 1'h1;
  assign tags_MPORT_17_en = reset;
  assign tags_MPORT_18_data = 21'h0;
  assign tags_MPORT_18_addr = 6'h10;
  assign tags_MPORT_18_mask = 1'h1;
  assign tags_MPORT_18_en = reset;
  assign tags_MPORT_19_data = 21'h0;
  assign tags_MPORT_19_addr = 6'h11;
  assign tags_MPORT_19_mask = 1'h1;
  assign tags_MPORT_19_en = reset;
  assign tags_MPORT_20_data = 21'h0;
  assign tags_MPORT_20_addr = 6'h12;
  assign tags_MPORT_20_mask = 1'h1;
  assign tags_MPORT_20_en = reset;
  assign tags_MPORT_21_data = 21'h0;
  assign tags_MPORT_21_addr = 6'h13;
  assign tags_MPORT_21_mask = 1'h1;
  assign tags_MPORT_21_en = reset;
  assign tags_MPORT_22_data = 21'h0;
  assign tags_MPORT_22_addr = 6'h14;
  assign tags_MPORT_22_mask = 1'h1;
  assign tags_MPORT_22_en = reset;
  assign tags_MPORT_23_data = 21'h0;
  assign tags_MPORT_23_addr = 6'h15;
  assign tags_MPORT_23_mask = 1'h1;
  assign tags_MPORT_23_en = reset;
  assign tags_MPORT_24_data = 21'h0;
  assign tags_MPORT_24_addr = 6'h16;
  assign tags_MPORT_24_mask = 1'h1;
  assign tags_MPORT_24_en = reset;
  assign tags_MPORT_25_data = 21'h0;
  assign tags_MPORT_25_addr = 6'h17;
  assign tags_MPORT_25_mask = 1'h1;
  assign tags_MPORT_25_en = reset;
  assign tags_MPORT_26_data = 21'h0;
  assign tags_MPORT_26_addr = 6'h18;
  assign tags_MPORT_26_mask = 1'h1;
  assign tags_MPORT_26_en = reset;
  assign tags_MPORT_27_data = 21'h0;
  assign tags_MPORT_27_addr = 6'h19;
  assign tags_MPORT_27_mask = 1'h1;
  assign tags_MPORT_27_en = reset;
  assign tags_MPORT_28_data = 21'h0;
  assign tags_MPORT_28_addr = 6'h1a;
  assign tags_MPORT_28_mask = 1'h1;
  assign tags_MPORT_28_en = reset;
  assign tags_MPORT_29_data = 21'h0;
  assign tags_MPORT_29_addr = 6'h1b;
  assign tags_MPORT_29_mask = 1'h1;
  assign tags_MPORT_29_en = reset;
  assign tags_MPORT_30_data = 21'h0;
  assign tags_MPORT_30_addr = 6'h1c;
  assign tags_MPORT_30_mask = 1'h1;
  assign tags_MPORT_30_en = reset;
  assign tags_MPORT_31_data = 21'h0;
  assign tags_MPORT_31_addr = 6'h1d;
  assign tags_MPORT_31_mask = 1'h1;
  assign tags_MPORT_31_en = reset;
  assign tags_MPORT_32_data = 21'h0;
  assign tags_MPORT_32_addr = 6'h1e;
  assign tags_MPORT_32_mask = 1'h1;
  assign tags_MPORT_32_en = reset;
  assign tags_MPORT_33_data = 21'h0;
  assign tags_MPORT_33_addr = 6'h1f;
  assign tags_MPORT_33_mask = 1'h1;
  assign tags_MPORT_33_en = reset;
  assign tags_MPORT_34_data = 21'h0;
  assign tags_MPORT_34_addr = 6'h20;
  assign tags_MPORT_34_mask = 1'h1;
  assign tags_MPORT_34_en = reset;
  assign tags_MPORT_35_data = 21'h0;
  assign tags_MPORT_35_addr = 6'h21;
  assign tags_MPORT_35_mask = 1'h1;
  assign tags_MPORT_35_en = reset;
  assign tags_MPORT_36_data = 21'h0;
  assign tags_MPORT_36_addr = 6'h22;
  assign tags_MPORT_36_mask = 1'h1;
  assign tags_MPORT_36_en = reset;
  assign tags_MPORT_37_data = 21'h0;
  assign tags_MPORT_37_addr = 6'h23;
  assign tags_MPORT_37_mask = 1'h1;
  assign tags_MPORT_37_en = reset;
  assign tags_MPORT_38_data = 21'h0;
  assign tags_MPORT_38_addr = 6'h24;
  assign tags_MPORT_38_mask = 1'h1;
  assign tags_MPORT_38_en = reset;
  assign tags_MPORT_39_data = 21'h0;
  assign tags_MPORT_39_addr = 6'h25;
  assign tags_MPORT_39_mask = 1'h1;
  assign tags_MPORT_39_en = reset;
  assign tags_MPORT_40_data = 21'h0;
  assign tags_MPORT_40_addr = 6'h26;
  assign tags_MPORT_40_mask = 1'h1;
  assign tags_MPORT_40_en = reset;
  assign tags_MPORT_41_data = 21'h0;
  assign tags_MPORT_41_addr = 6'h27;
  assign tags_MPORT_41_mask = 1'h1;
  assign tags_MPORT_41_en = reset;
  assign tags_MPORT_42_data = 21'h0;
  assign tags_MPORT_42_addr = 6'h28;
  assign tags_MPORT_42_mask = 1'h1;
  assign tags_MPORT_42_en = reset;
  assign tags_MPORT_43_data = 21'h0;
  assign tags_MPORT_43_addr = 6'h29;
  assign tags_MPORT_43_mask = 1'h1;
  assign tags_MPORT_43_en = reset;
  assign tags_MPORT_44_data = 21'h0;
  assign tags_MPORT_44_addr = 6'h2a;
  assign tags_MPORT_44_mask = 1'h1;
  assign tags_MPORT_44_en = reset;
  assign tags_MPORT_45_data = 21'h0;
  assign tags_MPORT_45_addr = 6'h2b;
  assign tags_MPORT_45_mask = 1'h1;
  assign tags_MPORT_45_en = reset;
  assign tags_MPORT_46_data = 21'h0;
  assign tags_MPORT_46_addr = 6'h2c;
  assign tags_MPORT_46_mask = 1'h1;
  assign tags_MPORT_46_en = reset;
  assign tags_MPORT_47_data = 21'h0;
  assign tags_MPORT_47_addr = 6'h2d;
  assign tags_MPORT_47_mask = 1'h1;
  assign tags_MPORT_47_en = reset;
  assign tags_MPORT_48_data = 21'h0;
  assign tags_MPORT_48_addr = 6'h2e;
  assign tags_MPORT_48_mask = 1'h1;
  assign tags_MPORT_48_en = reset;
  assign tags_MPORT_49_data = 21'h0;
  assign tags_MPORT_49_addr = 6'h2f;
  assign tags_MPORT_49_mask = 1'h1;
  assign tags_MPORT_49_en = reset;
  assign tags_MPORT_50_data = 21'h0;
  assign tags_MPORT_50_addr = 6'h30;
  assign tags_MPORT_50_mask = 1'h1;
  assign tags_MPORT_50_en = reset;
  assign tags_MPORT_51_data = 21'h0;
  assign tags_MPORT_51_addr = 6'h31;
  assign tags_MPORT_51_mask = 1'h1;
  assign tags_MPORT_51_en = reset;
  assign tags_MPORT_52_data = 21'h0;
  assign tags_MPORT_52_addr = 6'h32;
  assign tags_MPORT_52_mask = 1'h1;
  assign tags_MPORT_52_en = reset;
  assign tags_MPORT_53_data = 21'h0;
  assign tags_MPORT_53_addr = 6'h33;
  assign tags_MPORT_53_mask = 1'h1;
  assign tags_MPORT_53_en = reset;
  assign tags_MPORT_54_data = 21'h0;
  assign tags_MPORT_54_addr = 6'h34;
  assign tags_MPORT_54_mask = 1'h1;
  assign tags_MPORT_54_en = reset;
  assign tags_MPORT_55_data = 21'h0;
  assign tags_MPORT_55_addr = 6'h35;
  assign tags_MPORT_55_mask = 1'h1;
  assign tags_MPORT_55_en = reset;
  assign tags_MPORT_56_data = 21'h0;
  assign tags_MPORT_56_addr = 6'h36;
  assign tags_MPORT_56_mask = 1'h1;
  assign tags_MPORT_56_en = reset;
  assign tags_MPORT_57_data = 21'h0;
  assign tags_MPORT_57_addr = 6'h37;
  assign tags_MPORT_57_mask = 1'h1;
  assign tags_MPORT_57_en = reset;
  assign tags_MPORT_58_data = 21'h0;
  assign tags_MPORT_58_addr = 6'h38;
  assign tags_MPORT_58_mask = 1'h1;
  assign tags_MPORT_58_en = reset;
  assign tags_MPORT_59_data = 21'h0;
  assign tags_MPORT_59_addr = 6'h39;
  assign tags_MPORT_59_mask = 1'h1;
  assign tags_MPORT_59_en = reset;
  assign tags_MPORT_60_data = 21'h0;
  assign tags_MPORT_60_addr = 6'h3a;
  assign tags_MPORT_60_mask = 1'h1;
  assign tags_MPORT_60_en = reset;
  assign tags_MPORT_61_data = 21'h0;
  assign tags_MPORT_61_addr = 6'h3b;
  assign tags_MPORT_61_mask = 1'h1;
  assign tags_MPORT_61_en = reset;
  assign tags_MPORT_62_data = 21'h0;
  assign tags_MPORT_62_addr = 6'h3c;
  assign tags_MPORT_62_mask = 1'h1;
  assign tags_MPORT_62_en = reset;
  assign tags_MPORT_63_data = 21'h0;
  assign tags_MPORT_63_addr = 6'h3d;
  assign tags_MPORT_63_mask = 1'h1;
  assign tags_MPORT_63_en = reset;
  assign tags_MPORT_64_data = 21'h0;
  assign tags_MPORT_64_addr = 6'h3e;
  assign tags_MPORT_64_mask = 1'h1;
  assign tags_MPORT_64_en = reset;
  assign tags_MPORT_65_data = 21'h0;
  assign tags_MPORT_65_addr = 6'h3f;
  assign tags_MPORT_65_mask = 1'h1;
  assign tags_MPORT_65_en = reset;
  assign io_tag_r = tags_MPORT_1_data; // @[Cache.scala 48:12]
  assign io_dirty_r_async = 6'h3f == io_idx ? dirty_63 : _GEN_199; // @[Cache.scala 51:{20,20}]
  assign io_valid_r_async = 6'h3f == io_idx ? valid_63 : _GEN_263; // @[Cache.scala 52:{20,20}]
  always @(posedge clock) begin
    if (tags_MPORT_en & tags_MPORT_mask) begin
      tags[tags_MPORT_addr] <= tags_MPORT_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_2_en & tags_MPORT_2_mask) begin
      tags[tags_MPORT_2_addr] <= tags_MPORT_2_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_3_en & tags_MPORT_3_mask) begin
      tags[tags_MPORT_3_addr] <= tags_MPORT_3_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_4_en & tags_MPORT_4_mask) begin
      tags[tags_MPORT_4_addr] <= tags_MPORT_4_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_5_en & tags_MPORT_5_mask) begin
      tags[tags_MPORT_5_addr] <= tags_MPORT_5_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_6_en & tags_MPORT_6_mask) begin
      tags[tags_MPORT_6_addr] <= tags_MPORT_6_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_7_en & tags_MPORT_7_mask) begin
      tags[tags_MPORT_7_addr] <= tags_MPORT_7_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_8_en & tags_MPORT_8_mask) begin
      tags[tags_MPORT_8_addr] <= tags_MPORT_8_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_9_en & tags_MPORT_9_mask) begin
      tags[tags_MPORT_9_addr] <= tags_MPORT_9_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_10_en & tags_MPORT_10_mask) begin
      tags[tags_MPORT_10_addr] <= tags_MPORT_10_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_11_en & tags_MPORT_11_mask) begin
      tags[tags_MPORT_11_addr] <= tags_MPORT_11_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_12_en & tags_MPORT_12_mask) begin
      tags[tags_MPORT_12_addr] <= tags_MPORT_12_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_13_en & tags_MPORT_13_mask) begin
      tags[tags_MPORT_13_addr] <= tags_MPORT_13_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_14_en & tags_MPORT_14_mask) begin
      tags[tags_MPORT_14_addr] <= tags_MPORT_14_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_15_en & tags_MPORT_15_mask) begin
      tags[tags_MPORT_15_addr] <= tags_MPORT_15_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_16_en & tags_MPORT_16_mask) begin
      tags[tags_MPORT_16_addr] <= tags_MPORT_16_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_17_en & tags_MPORT_17_mask) begin
      tags[tags_MPORT_17_addr] <= tags_MPORT_17_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_18_en & tags_MPORT_18_mask) begin
      tags[tags_MPORT_18_addr] <= tags_MPORT_18_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_19_en & tags_MPORT_19_mask) begin
      tags[tags_MPORT_19_addr] <= tags_MPORT_19_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_20_en & tags_MPORT_20_mask) begin
      tags[tags_MPORT_20_addr] <= tags_MPORT_20_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_21_en & tags_MPORT_21_mask) begin
      tags[tags_MPORT_21_addr] <= tags_MPORT_21_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_22_en & tags_MPORT_22_mask) begin
      tags[tags_MPORT_22_addr] <= tags_MPORT_22_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_23_en & tags_MPORT_23_mask) begin
      tags[tags_MPORT_23_addr] <= tags_MPORT_23_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_24_en & tags_MPORT_24_mask) begin
      tags[tags_MPORT_24_addr] <= tags_MPORT_24_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_25_en & tags_MPORT_25_mask) begin
      tags[tags_MPORT_25_addr] <= tags_MPORT_25_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_26_en & tags_MPORT_26_mask) begin
      tags[tags_MPORT_26_addr] <= tags_MPORT_26_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_27_en & tags_MPORT_27_mask) begin
      tags[tags_MPORT_27_addr] <= tags_MPORT_27_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_28_en & tags_MPORT_28_mask) begin
      tags[tags_MPORT_28_addr] <= tags_MPORT_28_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_29_en & tags_MPORT_29_mask) begin
      tags[tags_MPORT_29_addr] <= tags_MPORT_29_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_30_en & tags_MPORT_30_mask) begin
      tags[tags_MPORT_30_addr] <= tags_MPORT_30_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_31_en & tags_MPORT_31_mask) begin
      tags[tags_MPORT_31_addr] <= tags_MPORT_31_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_32_en & tags_MPORT_32_mask) begin
      tags[tags_MPORT_32_addr] <= tags_MPORT_32_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_33_en & tags_MPORT_33_mask) begin
      tags[tags_MPORT_33_addr] <= tags_MPORT_33_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_34_en & tags_MPORT_34_mask) begin
      tags[tags_MPORT_34_addr] <= tags_MPORT_34_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_35_en & tags_MPORT_35_mask) begin
      tags[tags_MPORT_35_addr] <= tags_MPORT_35_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_36_en & tags_MPORT_36_mask) begin
      tags[tags_MPORT_36_addr] <= tags_MPORT_36_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_37_en & tags_MPORT_37_mask) begin
      tags[tags_MPORT_37_addr] <= tags_MPORT_37_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_38_en & tags_MPORT_38_mask) begin
      tags[tags_MPORT_38_addr] <= tags_MPORT_38_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_39_en & tags_MPORT_39_mask) begin
      tags[tags_MPORT_39_addr] <= tags_MPORT_39_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_40_en & tags_MPORT_40_mask) begin
      tags[tags_MPORT_40_addr] <= tags_MPORT_40_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_41_en & tags_MPORT_41_mask) begin
      tags[tags_MPORT_41_addr] <= tags_MPORT_41_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_42_en & tags_MPORT_42_mask) begin
      tags[tags_MPORT_42_addr] <= tags_MPORT_42_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_43_en & tags_MPORT_43_mask) begin
      tags[tags_MPORT_43_addr] <= tags_MPORT_43_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_44_en & tags_MPORT_44_mask) begin
      tags[tags_MPORT_44_addr] <= tags_MPORT_44_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_45_en & tags_MPORT_45_mask) begin
      tags[tags_MPORT_45_addr] <= tags_MPORT_45_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_46_en & tags_MPORT_46_mask) begin
      tags[tags_MPORT_46_addr] <= tags_MPORT_46_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_47_en & tags_MPORT_47_mask) begin
      tags[tags_MPORT_47_addr] <= tags_MPORT_47_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_48_en & tags_MPORT_48_mask) begin
      tags[tags_MPORT_48_addr] <= tags_MPORT_48_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_49_en & tags_MPORT_49_mask) begin
      tags[tags_MPORT_49_addr] <= tags_MPORT_49_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_50_en & tags_MPORT_50_mask) begin
      tags[tags_MPORT_50_addr] <= tags_MPORT_50_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_51_en & tags_MPORT_51_mask) begin
      tags[tags_MPORT_51_addr] <= tags_MPORT_51_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_52_en & tags_MPORT_52_mask) begin
      tags[tags_MPORT_52_addr] <= tags_MPORT_52_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_53_en & tags_MPORT_53_mask) begin
      tags[tags_MPORT_53_addr] <= tags_MPORT_53_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_54_en & tags_MPORT_54_mask) begin
      tags[tags_MPORT_54_addr] <= tags_MPORT_54_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_55_en & tags_MPORT_55_mask) begin
      tags[tags_MPORT_55_addr] <= tags_MPORT_55_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_56_en & tags_MPORT_56_mask) begin
      tags[tags_MPORT_56_addr] <= tags_MPORT_56_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_57_en & tags_MPORT_57_mask) begin
      tags[tags_MPORT_57_addr] <= tags_MPORT_57_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_58_en & tags_MPORT_58_mask) begin
      tags[tags_MPORT_58_addr] <= tags_MPORT_58_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_59_en & tags_MPORT_59_mask) begin
      tags[tags_MPORT_59_addr] <= tags_MPORT_59_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_60_en & tags_MPORT_60_mask) begin
      tags[tags_MPORT_60_addr] <= tags_MPORT_60_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_61_en & tags_MPORT_61_mask) begin
      tags[tags_MPORT_61_addr] <= tags_MPORT_61_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_62_en & tags_MPORT_62_mask) begin
      tags[tags_MPORT_62_addr] <= tags_MPORT_62_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_63_en & tags_MPORT_63_mask) begin
      tags[tags_MPORT_63_addr] <= tags_MPORT_63_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_64_en & tags_MPORT_64_mask) begin
      tags[tags_MPORT_64_addr] <= tags_MPORT_64_data; // @[Cache.scala 33:25]
    end
    if (tags_MPORT_65_en & tags_MPORT_65_mask) begin
      tags[tags_MPORT_65_addr] <= tags_MPORT_65_data; // @[Cache.scala 33:25]
    end
//     tags_MPORT_1_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      tags_MPORT_1_addr_pipe_0 <= io_idx;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_0 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_0 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_0 <= _GEN_0;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_1 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_1 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_1 <= _GEN_1;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_2 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_2 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_2 <= _GEN_2;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_3 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_3 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_3 <= _GEN_3;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_4 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_4 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_4 <= _GEN_4;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_5 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_5 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_5 <= _GEN_5;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_6 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_6 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_6 <= _GEN_6;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_7 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_7 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_7 <= _GEN_7;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_8 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_8 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_8 <= _GEN_8;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_9 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_9 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_9 <= _GEN_9;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_10 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_10 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_10 <= _GEN_10;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_11 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_11 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_11 <= _GEN_11;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_12 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_12 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_12 <= _GEN_12;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_13 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_13 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_13 <= _GEN_13;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_14 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_14 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_14 <= _GEN_14;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_15 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_15 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_15 <= _GEN_15;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_16 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_16 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_16 <= _GEN_16;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_17 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_17 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_17 <= _GEN_17;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_18 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_18 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_18 <= _GEN_18;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_19 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_19 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_19 <= _GEN_19;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_20 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_20 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_20 <= _GEN_20;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_21 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_21 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_21 <= _GEN_21;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_22 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_22 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_22 <= _GEN_22;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_23 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_23 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_23 <= _GEN_23;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_24 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_24 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_24 <= _GEN_24;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_25 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_25 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_25 <= _GEN_25;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_26 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_26 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_26 <= _GEN_26;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_27 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_27 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_27 <= _GEN_27;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_28 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_28 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_28 <= _GEN_28;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_29 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_29 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_29 <= _GEN_29;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_30 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_30 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_30 <= _GEN_30;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_31 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_31 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_31 <= _GEN_31;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_32 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_32 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_32 <= _GEN_32;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_33 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_33 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_33 <= _GEN_33;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_34 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_34 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_34 <= _GEN_34;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_35 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_35 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_35 <= _GEN_35;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_36 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_36 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_36 <= _GEN_36;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_37 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_37 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_37 <= _GEN_37;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_38 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_38 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_38 <= _GEN_38;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_39 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_39 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_39 <= _GEN_39;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_40 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_40 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_40 <= _GEN_40;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_41 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_41 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_41 <= _GEN_41;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_42 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_42 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_42 <= _GEN_42;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_43 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_43 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_43 <= _GEN_43;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_44 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_44 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_44 <= _GEN_44;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_45 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_45 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_45 <= _GEN_45;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_46 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_46 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_46 <= _GEN_46;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_47 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_47 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_47 <= _GEN_47;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_48 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_48 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_48 <= _GEN_48;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_49 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_49 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_49 <= _GEN_49;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_50 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_50 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_50 <= _GEN_50;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_51 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_51 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_51 <= _GEN_51;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_52 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_52 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_52 <= _GEN_52;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_53 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_53 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_53 <= _GEN_53;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_54 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_54 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_54 <= _GEN_54;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_55 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_55 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_55 <= _GEN_55;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_56 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_56 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_56 <= _GEN_56;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_57 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_57 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_57 <= _GEN_57;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_58 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_58 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_58 <= _GEN_58;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_59 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_59 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_59 <= _GEN_59;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_60 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_60 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_60 <= _GEN_60;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_61 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_61 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_61 <= _GEN_61;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_62 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_62 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_62 <= _GEN_62;
    end
    if (reset) begin // @[Cache.scala 35:22]
      valid_63 <= 1'h0; // @[Cache.scala 35:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      valid_63 <= 1'h0; // @[Cache.scala 63:16]
    end else if (io_tag_wen) begin // @[Cache.scala 44:21]
      valid_63 <= _GEN_63;
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_0 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_0 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h0 == io_idx) begin // @[Cache.scala 56:16]
        dirty_0 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_1 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_1 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h1 == io_idx) begin // @[Cache.scala 56:16]
        dirty_1 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_2 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_2 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h2 == io_idx) begin // @[Cache.scala 56:16]
        dirty_2 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_3 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_3 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h3 == io_idx) begin // @[Cache.scala 56:16]
        dirty_3 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_4 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_4 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h4 == io_idx) begin // @[Cache.scala 56:16]
        dirty_4 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_5 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_5 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h5 == io_idx) begin // @[Cache.scala 56:16]
        dirty_5 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_6 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_6 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h6 == io_idx) begin // @[Cache.scala 56:16]
        dirty_6 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_7 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_7 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h7 == io_idx) begin // @[Cache.scala 56:16]
        dirty_7 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_8 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_8 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h8 == io_idx) begin // @[Cache.scala 56:16]
        dirty_8 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_9 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_9 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h9 == io_idx) begin // @[Cache.scala 56:16]
        dirty_9 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_10 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_10 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'ha == io_idx) begin // @[Cache.scala 56:16]
        dirty_10 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_11 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_11 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'hb == io_idx) begin // @[Cache.scala 56:16]
        dirty_11 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_12 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_12 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'hc == io_idx) begin // @[Cache.scala 56:16]
        dirty_12 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_13 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_13 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'hd == io_idx) begin // @[Cache.scala 56:16]
        dirty_13 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_14 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_14 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'he == io_idx) begin // @[Cache.scala 56:16]
        dirty_14 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_15 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_15 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'hf == io_idx) begin // @[Cache.scala 56:16]
        dirty_15 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_16 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_16 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h10 == io_idx) begin // @[Cache.scala 56:16]
        dirty_16 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_17 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_17 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h11 == io_idx) begin // @[Cache.scala 56:16]
        dirty_17 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_18 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_18 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h12 == io_idx) begin // @[Cache.scala 56:16]
        dirty_18 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_19 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_19 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h13 == io_idx) begin // @[Cache.scala 56:16]
        dirty_19 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_20 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_20 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h14 == io_idx) begin // @[Cache.scala 56:16]
        dirty_20 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_21 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_21 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h15 == io_idx) begin // @[Cache.scala 56:16]
        dirty_21 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_22 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_22 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h16 == io_idx) begin // @[Cache.scala 56:16]
        dirty_22 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_23 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_23 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h17 == io_idx) begin // @[Cache.scala 56:16]
        dirty_23 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_24 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_24 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h18 == io_idx) begin // @[Cache.scala 56:16]
        dirty_24 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_25 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_25 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h19 == io_idx) begin // @[Cache.scala 56:16]
        dirty_25 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_26 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_26 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h1a == io_idx) begin // @[Cache.scala 56:16]
        dirty_26 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_27 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_27 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h1b == io_idx) begin // @[Cache.scala 56:16]
        dirty_27 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_28 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_28 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h1c == io_idx) begin // @[Cache.scala 56:16]
        dirty_28 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_29 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_29 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h1d == io_idx) begin // @[Cache.scala 56:16]
        dirty_29 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_30 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_30 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h1e == io_idx) begin // @[Cache.scala 56:16]
        dirty_30 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_31 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_31 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h1f == io_idx) begin // @[Cache.scala 56:16]
        dirty_31 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_32 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_32 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h20 == io_idx) begin // @[Cache.scala 56:16]
        dirty_32 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_33 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_33 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h21 == io_idx) begin // @[Cache.scala 56:16]
        dirty_33 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_34 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_34 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h22 == io_idx) begin // @[Cache.scala 56:16]
        dirty_34 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_35 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_35 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h23 == io_idx) begin // @[Cache.scala 56:16]
        dirty_35 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_36 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_36 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h24 == io_idx) begin // @[Cache.scala 56:16]
        dirty_36 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_37 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_37 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h25 == io_idx) begin // @[Cache.scala 56:16]
        dirty_37 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_38 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_38 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h26 == io_idx) begin // @[Cache.scala 56:16]
        dirty_38 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_39 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_39 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h27 == io_idx) begin // @[Cache.scala 56:16]
        dirty_39 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_40 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_40 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h28 == io_idx) begin // @[Cache.scala 56:16]
        dirty_40 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_41 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_41 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h29 == io_idx) begin // @[Cache.scala 56:16]
        dirty_41 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_42 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_42 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h2a == io_idx) begin // @[Cache.scala 56:16]
        dirty_42 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_43 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_43 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h2b == io_idx) begin // @[Cache.scala 56:16]
        dirty_43 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_44 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_44 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h2c == io_idx) begin // @[Cache.scala 56:16]
        dirty_44 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_45 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_45 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h2d == io_idx) begin // @[Cache.scala 56:16]
        dirty_45 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_46 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_46 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h2e == io_idx) begin // @[Cache.scala 56:16]
        dirty_46 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_47 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_47 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h2f == io_idx) begin // @[Cache.scala 56:16]
        dirty_47 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_48 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_48 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h30 == io_idx) begin // @[Cache.scala 56:16]
        dirty_48 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_49 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_49 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h31 == io_idx) begin // @[Cache.scala 56:16]
        dirty_49 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_50 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_50 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h32 == io_idx) begin // @[Cache.scala 56:16]
        dirty_50 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_51 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_51 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h33 == io_idx) begin // @[Cache.scala 56:16]
        dirty_51 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_52 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_52 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h34 == io_idx) begin // @[Cache.scala 56:16]
        dirty_52 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_53 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_53 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h35 == io_idx) begin // @[Cache.scala 56:16]
        dirty_53 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_54 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_54 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h36 == io_idx) begin // @[Cache.scala 56:16]
        dirty_54 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_55 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_55 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h37 == io_idx) begin // @[Cache.scala 56:16]
        dirty_55 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_56 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_56 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h38 == io_idx) begin // @[Cache.scala 56:16]
        dirty_56 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_57 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_57 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h39 == io_idx) begin // @[Cache.scala 56:16]
        dirty_57 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_58 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_58 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h3a == io_idx) begin // @[Cache.scala 56:16]
        dirty_58 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_59 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_59 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h3b == io_idx) begin // @[Cache.scala 56:16]
        dirty_59 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_60 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_60 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h3c == io_idx) begin // @[Cache.scala 56:16]
        dirty_60 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_61 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_61 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h3d == io_idx) begin // @[Cache.scala 56:16]
        dirty_61 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_62 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_62 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h3e == io_idx) begin // @[Cache.scala 56:16]
        dirty_62 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
    if (reset) begin // @[Cache.scala 39:22]
      dirty_63 <= 1'h0; // @[Cache.scala 39:22]
    end else if (io_invalidate) begin // @[Cache.scala 60:24]
      dirty_63 <= 1'h0; // @[Cache.scala 62:16]
    end else if (io_dirty_wen) begin // @[Cache.scala 55:23]
      if (6'h3f == io_idx) begin // @[Cache.scala 56:16]
        dirty_63 <= io_dirty_w; // @[Cache.scala 56:16]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tags[initvar] = _RAND_0[20:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
//   tags_MPORT_1_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  tags_MPORT_1_addr_pipe_0 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  valid_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  valid_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  valid_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid_4 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  valid_5 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_6 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_7 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  valid_8 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_9 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid_10 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  valid_11 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  valid_12 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  valid_13 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_14 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_15 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_16 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_17 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_18 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_19 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_20 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_21 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_22 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_23 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_24 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_25 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_26 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_27 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_28 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_29 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_30 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_31 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_32 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_33 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_34 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_35 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_36 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  valid_37 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  valid_38 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  valid_39 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  valid_40 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  valid_41 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  valid_42 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  valid_43 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  valid_44 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  valid_45 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  valid_46 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  valid_47 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  valid_48 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  valid_49 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  valid_50 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  valid_51 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  valid_52 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  valid_53 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  valid_54 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  valid_55 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  valid_56 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  valid_57 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  valid_58 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  valid_59 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  valid_60 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  valid_61 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_62 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_63 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  dirty_0 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  dirty_1 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  dirty_2 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  dirty_3 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  dirty_4 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  dirty_5 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  dirty_6 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  dirty_7 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  dirty_8 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  dirty_9 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  dirty_10 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  dirty_11 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  dirty_12 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  dirty_13 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  dirty_14 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  dirty_15 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  dirty_16 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  dirty_17 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  dirty_18 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  dirty_19 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  dirty_20 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  dirty_21 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  dirty_22 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  dirty_23 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  dirty_24 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  dirty_25 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  dirty_26 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  dirty_27 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  dirty_28 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  dirty_29 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  dirty_30 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  dirty_31 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  dirty_32 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  dirty_33 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  dirty_34 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  dirty_35 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  dirty_36 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  dirty_37 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  dirty_38 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  dirty_39 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  dirty_40 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  dirty_41 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  dirty_42 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  dirty_43 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  dirty_44 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  dirty_45 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  dirty_46 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  dirty_47 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  dirty_48 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  dirty_49 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  dirty_50 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  dirty_51 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  dirty_52 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  dirty_53 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  dirty_54 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  dirty_55 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  dirty_56 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  dirty_57 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  dirty_58 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  dirty_59 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  dirty_60 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  dirty_61 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  dirty_62 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  dirty_63 = _RAND_130[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_Cache(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [67:0] io_in_req_bits_user,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output [67:0] io_in_resp_bits_user,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output        io_out_req_bits_aen,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_req_bits_wlast,
  output        io_out_req_bits_wen,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_out_resp_bits_rlast,
  input         fence_i_0,
  input         dcache_fi_complete,
  input         sq_empty_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [95:0] _RAND_205;
  reg [127:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [127:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [63:0] _RAND_215;
`endif // RANDOMIZE_REG_INIT
  wire  sram_0_clock; // @[Cache.scala 89:22]
  wire  sram_0_io_en; // @[Cache.scala 89:22]
  wire  sram_0_io_wen; // @[Cache.scala 89:22]
  wire [5:0] sram_0_io_addr; // @[Cache.scala 89:22]
  wire [127:0] sram_0_io_wdata; // @[Cache.scala 89:22]
  wire [127:0] sram_0_io_rdata; // @[Cache.scala 89:22]
  wire  sram_1_clock; // @[Cache.scala 89:22]
  wire  sram_1_io_en; // @[Cache.scala 89:22]
  wire  sram_1_io_wen; // @[Cache.scala 89:22]
  wire [5:0] sram_1_io_addr; // @[Cache.scala 89:22]
  wire [127:0] sram_1_io_wdata; // @[Cache.scala 89:22]
  wire [127:0] sram_1_io_rdata; // @[Cache.scala 89:22]
  wire  sram_2_clock; // @[Cache.scala 89:22]
  wire  sram_2_io_en; // @[Cache.scala 89:22]
  wire  sram_2_io_wen; // @[Cache.scala 89:22]
  wire [5:0] sram_2_io_addr; // @[Cache.scala 89:22]
  wire [127:0] sram_2_io_wdata; // @[Cache.scala 89:22]
  wire [127:0] sram_2_io_rdata; // @[Cache.scala 89:22]
  wire  sram_3_clock; // @[Cache.scala 89:22]
  wire  sram_3_io_en; // @[Cache.scala 89:22]
  wire  sram_3_io_wen; // @[Cache.scala 89:22]
  wire [5:0] sram_3_io_addr; // @[Cache.scala 89:22]
  wire [127:0] sram_3_io_wdata; // @[Cache.scala 89:22]
  wire [127:0] sram_3_io_rdata; // @[Cache.scala 89:22]
  wire  meta_0_clock; // @[Cache.scala 97:22]
  wire  meta_0_reset; // @[Cache.scala 97:22]
  wire [5:0] meta_0_io_idx; // @[Cache.scala 97:22]
  wire [20:0] meta_0_io_tag_r; // @[Cache.scala 97:22]
  wire [20:0] meta_0_io_tag_w; // @[Cache.scala 97:22]
  wire  meta_0_io_tag_wen; // @[Cache.scala 97:22]
  wire  meta_0_io_dirty_r_async; // @[Cache.scala 97:22]
  wire  meta_0_io_dirty_w; // @[Cache.scala 97:22]
  wire  meta_0_io_dirty_wen; // @[Cache.scala 97:22]
  wire  meta_0_io_valid_r_async; // @[Cache.scala 97:22]
  wire  meta_0_io_invalidate; // @[Cache.scala 97:22]
  wire  meta_1_clock; // @[Cache.scala 97:22]
  wire  meta_1_reset; // @[Cache.scala 97:22]
  wire [5:0] meta_1_io_idx; // @[Cache.scala 97:22]
  wire [20:0] meta_1_io_tag_r; // @[Cache.scala 97:22]
  wire [20:0] meta_1_io_tag_w; // @[Cache.scala 97:22]
  wire  meta_1_io_tag_wen; // @[Cache.scala 97:22]
  wire  meta_1_io_dirty_r_async; // @[Cache.scala 97:22]
  wire  meta_1_io_dirty_w; // @[Cache.scala 97:22]
  wire  meta_1_io_dirty_wen; // @[Cache.scala 97:22]
  wire  meta_1_io_valid_r_async; // @[Cache.scala 97:22]
  wire  meta_1_io_invalidate; // @[Cache.scala 97:22]
  wire  meta_2_clock; // @[Cache.scala 97:22]
  wire  meta_2_reset; // @[Cache.scala 97:22]
  wire [5:0] meta_2_io_idx; // @[Cache.scala 97:22]
  wire [20:0] meta_2_io_tag_r; // @[Cache.scala 97:22]
  wire [20:0] meta_2_io_tag_w; // @[Cache.scala 97:22]
  wire  meta_2_io_tag_wen; // @[Cache.scala 97:22]
  wire  meta_2_io_dirty_r_async; // @[Cache.scala 97:22]
  wire  meta_2_io_dirty_w; // @[Cache.scala 97:22]
  wire  meta_2_io_dirty_wen; // @[Cache.scala 97:22]
  wire  meta_2_io_valid_r_async; // @[Cache.scala 97:22]
  wire  meta_2_io_invalidate; // @[Cache.scala 97:22]
  wire  meta_3_clock; // @[Cache.scala 97:22]
  wire  meta_3_reset; // @[Cache.scala 97:22]
  wire [5:0] meta_3_io_idx; // @[Cache.scala 97:22]
  wire [20:0] meta_3_io_tag_r; // @[Cache.scala 97:22]
  wire [20:0] meta_3_io_tag_w; // @[Cache.scala 97:22]
  wire  meta_3_io_tag_wen; // @[Cache.scala 97:22]
  wire  meta_3_io_dirty_r_async; // @[Cache.scala 97:22]
  wire  meta_3_io_dirty_w; // @[Cache.scala 97:22]
  wire  meta_3_io_dirty_wen; // @[Cache.scala 97:22]
  wire  meta_3_io_valid_r_async; // @[Cache.scala 97:22]
  wire  meta_3_io_invalidate; // @[Cache.scala 97:22]
  reg  REG; // @[Cache.scala 123:59]
  reg  REG_1; // @[Cache.scala 123:59]
  reg  REG_2; // @[Cache.scala 123:59]
  reg  REG_3; // @[Cache.scala 123:59]
  reg  REG_4; // @[Cache.scala 124:59]
  reg  REG_5; // @[Cache.scala 124:59]
  reg  REG_6; // @[Cache.scala 124:59]
  reg  REG_7; // @[Cache.scala 124:59]
  reg  plru0_0; // @[Cache.scala 129:22]
  reg  plru0_1; // @[Cache.scala 129:22]
  reg  plru0_2; // @[Cache.scala 129:22]
  reg  plru0_3; // @[Cache.scala 129:22]
  reg  plru0_4; // @[Cache.scala 129:22]
  reg  plru0_5; // @[Cache.scala 129:22]
  reg  plru0_6; // @[Cache.scala 129:22]
  reg  plru0_7; // @[Cache.scala 129:22]
  reg  plru0_8; // @[Cache.scala 129:22]
  reg  plru0_9; // @[Cache.scala 129:22]
  reg  plru0_10; // @[Cache.scala 129:22]
  reg  plru0_11; // @[Cache.scala 129:22]
  reg  plru0_12; // @[Cache.scala 129:22]
  reg  plru0_13; // @[Cache.scala 129:22]
  reg  plru0_14; // @[Cache.scala 129:22]
  reg  plru0_15; // @[Cache.scala 129:22]
  reg  plru0_16; // @[Cache.scala 129:22]
  reg  plru0_17; // @[Cache.scala 129:22]
  reg  plru0_18; // @[Cache.scala 129:22]
  reg  plru0_19; // @[Cache.scala 129:22]
  reg  plru0_20; // @[Cache.scala 129:22]
  reg  plru0_21; // @[Cache.scala 129:22]
  reg  plru0_22; // @[Cache.scala 129:22]
  reg  plru0_23; // @[Cache.scala 129:22]
  reg  plru0_24; // @[Cache.scala 129:22]
  reg  plru0_25; // @[Cache.scala 129:22]
  reg  plru0_26; // @[Cache.scala 129:22]
  reg  plru0_27; // @[Cache.scala 129:22]
  reg  plru0_28; // @[Cache.scala 129:22]
  reg  plru0_29; // @[Cache.scala 129:22]
  reg  plru0_30; // @[Cache.scala 129:22]
  reg  plru0_31; // @[Cache.scala 129:22]
  reg  plru0_32; // @[Cache.scala 129:22]
  reg  plru0_33; // @[Cache.scala 129:22]
  reg  plru0_34; // @[Cache.scala 129:22]
  reg  plru0_35; // @[Cache.scala 129:22]
  reg  plru0_36; // @[Cache.scala 129:22]
  reg  plru0_37; // @[Cache.scala 129:22]
  reg  plru0_38; // @[Cache.scala 129:22]
  reg  plru0_39; // @[Cache.scala 129:22]
  reg  plru0_40; // @[Cache.scala 129:22]
  reg  plru0_41; // @[Cache.scala 129:22]
  reg  plru0_42; // @[Cache.scala 129:22]
  reg  plru0_43; // @[Cache.scala 129:22]
  reg  plru0_44; // @[Cache.scala 129:22]
  reg  plru0_45; // @[Cache.scala 129:22]
  reg  plru0_46; // @[Cache.scala 129:22]
  reg  plru0_47; // @[Cache.scala 129:22]
  reg  plru0_48; // @[Cache.scala 129:22]
  reg  plru0_49; // @[Cache.scala 129:22]
  reg  plru0_50; // @[Cache.scala 129:22]
  reg  plru0_51; // @[Cache.scala 129:22]
  reg  plru0_52; // @[Cache.scala 129:22]
  reg  plru0_53; // @[Cache.scala 129:22]
  reg  plru0_54; // @[Cache.scala 129:22]
  reg  plru0_55; // @[Cache.scala 129:22]
  reg  plru0_56; // @[Cache.scala 129:22]
  reg  plru0_57; // @[Cache.scala 129:22]
  reg  plru0_58; // @[Cache.scala 129:22]
  reg  plru0_59; // @[Cache.scala 129:22]
  reg  plru0_60; // @[Cache.scala 129:22]
  reg  plru0_61; // @[Cache.scala 129:22]
  reg  plru0_62; // @[Cache.scala 129:22]
  reg  plru0_63; // @[Cache.scala 129:22]
  reg  plru1_0; // @[Cache.scala 131:22]
  reg  plru1_1; // @[Cache.scala 131:22]
  reg  plru1_2; // @[Cache.scala 131:22]
  reg  plru1_3; // @[Cache.scala 131:22]
  reg  plru1_4; // @[Cache.scala 131:22]
  reg  plru1_5; // @[Cache.scala 131:22]
  reg  plru1_6; // @[Cache.scala 131:22]
  reg  plru1_7; // @[Cache.scala 131:22]
  reg  plru1_8; // @[Cache.scala 131:22]
  reg  plru1_9; // @[Cache.scala 131:22]
  reg  plru1_10; // @[Cache.scala 131:22]
  reg  plru1_11; // @[Cache.scala 131:22]
  reg  plru1_12; // @[Cache.scala 131:22]
  reg  plru1_13; // @[Cache.scala 131:22]
  reg  plru1_14; // @[Cache.scala 131:22]
  reg  plru1_15; // @[Cache.scala 131:22]
  reg  plru1_16; // @[Cache.scala 131:22]
  reg  plru1_17; // @[Cache.scala 131:22]
  reg  plru1_18; // @[Cache.scala 131:22]
  reg  plru1_19; // @[Cache.scala 131:22]
  reg  plru1_20; // @[Cache.scala 131:22]
  reg  plru1_21; // @[Cache.scala 131:22]
  reg  plru1_22; // @[Cache.scala 131:22]
  reg  plru1_23; // @[Cache.scala 131:22]
  reg  plru1_24; // @[Cache.scala 131:22]
  reg  plru1_25; // @[Cache.scala 131:22]
  reg  plru1_26; // @[Cache.scala 131:22]
  reg  plru1_27; // @[Cache.scala 131:22]
  reg  plru1_28; // @[Cache.scala 131:22]
  reg  plru1_29; // @[Cache.scala 131:22]
  reg  plru1_30; // @[Cache.scala 131:22]
  reg  plru1_31; // @[Cache.scala 131:22]
  reg  plru1_32; // @[Cache.scala 131:22]
  reg  plru1_33; // @[Cache.scala 131:22]
  reg  plru1_34; // @[Cache.scala 131:22]
  reg  plru1_35; // @[Cache.scala 131:22]
  reg  plru1_36; // @[Cache.scala 131:22]
  reg  plru1_37; // @[Cache.scala 131:22]
  reg  plru1_38; // @[Cache.scala 131:22]
  reg  plru1_39; // @[Cache.scala 131:22]
  reg  plru1_40; // @[Cache.scala 131:22]
  reg  plru1_41; // @[Cache.scala 131:22]
  reg  plru1_42; // @[Cache.scala 131:22]
  reg  plru1_43; // @[Cache.scala 131:22]
  reg  plru1_44; // @[Cache.scala 131:22]
  reg  plru1_45; // @[Cache.scala 131:22]
  reg  plru1_46; // @[Cache.scala 131:22]
  reg  plru1_47; // @[Cache.scala 131:22]
  reg  plru1_48; // @[Cache.scala 131:22]
  reg  plru1_49; // @[Cache.scala 131:22]
  reg  plru1_50; // @[Cache.scala 131:22]
  reg  plru1_51; // @[Cache.scala 131:22]
  reg  plru1_52; // @[Cache.scala 131:22]
  reg  plru1_53; // @[Cache.scala 131:22]
  reg  plru1_54; // @[Cache.scala 131:22]
  reg  plru1_55; // @[Cache.scala 131:22]
  reg  plru1_56; // @[Cache.scala 131:22]
  reg  plru1_57; // @[Cache.scala 131:22]
  reg  plru1_58; // @[Cache.scala 131:22]
  reg  plru1_59; // @[Cache.scala 131:22]
  reg  plru1_60; // @[Cache.scala 131:22]
  reg  plru1_61; // @[Cache.scala 131:22]
  reg  plru1_62; // @[Cache.scala 131:22]
  reg  plru1_63; // @[Cache.scala 131:22]
  reg  plru2_0; // @[Cache.scala 133:22]
  reg  plru2_1; // @[Cache.scala 133:22]
  reg  plru2_2; // @[Cache.scala 133:22]
  reg  plru2_3; // @[Cache.scala 133:22]
  reg  plru2_4; // @[Cache.scala 133:22]
  reg  plru2_5; // @[Cache.scala 133:22]
  reg  plru2_6; // @[Cache.scala 133:22]
  reg  plru2_7; // @[Cache.scala 133:22]
  reg  plru2_8; // @[Cache.scala 133:22]
  reg  plru2_9; // @[Cache.scala 133:22]
  reg  plru2_10; // @[Cache.scala 133:22]
  reg  plru2_11; // @[Cache.scala 133:22]
  reg  plru2_12; // @[Cache.scala 133:22]
  reg  plru2_13; // @[Cache.scala 133:22]
  reg  plru2_14; // @[Cache.scala 133:22]
  reg  plru2_15; // @[Cache.scala 133:22]
  reg  plru2_16; // @[Cache.scala 133:22]
  reg  plru2_17; // @[Cache.scala 133:22]
  reg  plru2_18; // @[Cache.scala 133:22]
  reg  plru2_19; // @[Cache.scala 133:22]
  reg  plru2_20; // @[Cache.scala 133:22]
  reg  plru2_21; // @[Cache.scala 133:22]
  reg  plru2_22; // @[Cache.scala 133:22]
  reg  plru2_23; // @[Cache.scala 133:22]
  reg  plru2_24; // @[Cache.scala 133:22]
  reg  plru2_25; // @[Cache.scala 133:22]
  reg  plru2_26; // @[Cache.scala 133:22]
  reg  plru2_27; // @[Cache.scala 133:22]
  reg  plru2_28; // @[Cache.scala 133:22]
  reg  plru2_29; // @[Cache.scala 133:22]
  reg  plru2_30; // @[Cache.scala 133:22]
  reg  plru2_31; // @[Cache.scala 133:22]
  reg  plru2_32; // @[Cache.scala 133:22]
  reg  plru2_33; // @[Cache.scala 133:22]
  reg  plru2_34; // @[Cache.scala 133:22]
  reg  plru2_35; // @[Cache.scala 133:22]
  reg  plru2_36; // @[Cache.scala 133:22]
  reg  plru2_37; // @[Cache.scala 133:22]
  reg  plru2_38; // @[Cache.scala 133:22]
  reg  plru2_39; // @[Cache.scala 133:22]
  reg  plru2_40; // @[Cache.scala 133:22]
  reg  plru2_41; // @[Cache.scala 133:22]
  reg  plru2_42; // @[Cache.scala 133:22]
  reg  plru2_43; // @[Cache.scala 133:22]
  reg  plru2_44; // @[Cache.scala 133:22]
  reg  plru2_45; // @[Cache.scala 133:22]
  reg  plru2_46; // @[Cache.scala 133:22]
  reg  plru2_47; // @[Cache.scala 133:22]
  reg  plru2_48; // @[Cache.scala 133:22]
  reg  plru2_49; // @[Cache.scala 133:22]
  reg  plru2_50; // @[Cache.scala 133:22]
  reg  plru2_51; // @[Cache.scala 133:22]
  reg  plru2_52; // @[Cache.scala 133:22]
  reg  plru2_53; // @[Cache.scala 133:22]
  reg  plru2_54; // @[Cache.scala 133:22]
  reg  plru2_55; // @[Cache.scala 133:22]
  reg  plru2_56; // @[Cache.scala 133:22]
  reg  plru2_57; // @[Cache.scala 133:22]
  reg  plru2_58; // @[Cache.scala 133:22]
  reg  plru2_59; // @[Cache.scala 133:22]
  reg  plru2_60; // @[Cache.scala 133:22]
  reg  plru2_61; // @[Cache.scala 133:22]
  reg  plru2_62; // @[Cache.scala 133:22]
  reg  plru2_63; // @[Cache.scala 133:22]
  reg  REG_9; // @[Cache.scala 275:32]
  wire [20:0] tag_out_0 = meta_0_io_tag_r;
  reg [31:0] s2_addr; // @[Cache.scala 215:25]
  wire [20:0] s2_tag = s2_addr[30:10]; // @[Cache.scala 218:25]
  wire  hit_0 = tag_out_0 == s2_tag & REG; // @[Cache.scala 230:25]
  wire [20:0] tag_out_1 = meta_1_io_tag_r;
  wire  hit_1 = tag_out_1 == s2_tag & REG_1; // @[Cache.scala 230:25]
  wire [20:0] tag_out_2 = meta_2_io_tag_r;
  wire  hit_2 = tag_out_2 == s2_tag & REG_2; // @[Cache.scala 230:25]
  wire [20:0] tag_out_3 = meta_3_io_tag_r;
  wire  hit_3 = tag_out_3 == s2_tag & REG_3; // @[Cache.scala 230:25]
  wire [3:0] _T_8 = {hit_0,hit_1,hit_2,hit_3}; // @[Cat.scala 30:58]
  wire  s2_hit = |_T_8; // @[Cache.scala 232:25]
  reg  s2_reg_hit; // @[Cache.scala 239:27]
  wire  s2_hit_real = REG_9 ? s2_hit : s2_reg_hit; // @[Cache.scala 275:24]
  reg [3:0] state; // @[Cache.scala 213:22]
  wire  _T_18 = state == 4'h7; // @[Cache.scala 277:37]
  wire  _T_19 = state == 4'h0; // @[Cache.scala 277:59]
  wire  hit_ready = s2_hit_real & _T_19; // @[Cache.scala 276:31]
  wire  invalid_ready = state == 4'h8; // @[Cache.scala 279:30]
  wire  pipeline_ready = (hit_ready | _T_18) & io_in_resp_ready | invalid_ready; // @[Cache.scala 282:66]
  reg  fi_valid; // @[Utils.scala 34:20]
  wire  _GEN_0 = fence_i_0 | fi_valid; // @[Utils.scala 34:20 40:{20,24}]
  wire  fi_ready = pipeline_ready & sq_empty_0; // @[Cache.scala 163:33]
  wire  fi_fire = fi_valid & fi_ready; // @[Cache.scala 164:26]
  wire [5:0] s1_idx = io_in_req_bits_addr[9:4]; // @[Cache.scala 170:25]
  wire [5:0] _GEN_3 = pipeline_ready ? s1_idx : 6'h0; // @[Cache.scala 109:15 187:24 190:17]
  wire  s2_offs = s2_addr[3]; // @[Cache.scala 216:25]
  wire [5:0] s2_idx = s2_addr[9:4]; // @[Cache.scala 217:25]
  reg [67:0] s2_user; // @[Cache.scala 222:25]
  wire [3:0] _T_9 = {hit_3,hit_2,hit_1,hit_0}; // @[OneHot.scala 22:45]
  wire [1:0] hi_2 = _T_9[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] lo_2 = _T_9[1:0]; // @[OneHot.scala 31:18]
  wire  _T_10 = |hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _T_11 = hi_2 | lo_2; // @[OneHot.scala 32:28]
  wire [1:0] s2_way = {_T_10,_T_11[1]}; // @[Cat.scala 30:58]
  reg [127:0] s2_reg_rdata; // @[Cache.scala 241:29]
  reg  s2_reg_dirty; // @[Cache.scala 242:29]
  reg [20:0] s2_reg_tag_r; // @[Cache.scala 243:29]
  reg [127:0] s2_reg_dat_w; // @[Cache.scala 244:29]
  reg  REG_8; // @[Cache.scala 256:41]
  wire [127:0] sram_out_0 = sram_0_io_rdata;
  wire [127:0] sram_out_1 = sram_1_io_rdata;
  wire [127:0] _GEN_5 = 2'h1 == s2_way ? sram_out_1 : sram_out_0; // @[Cache.scala 261:{18,18}]
  wire [127:0] sram_out_2 = sram_2_io_rdata;
  wire [127:0] _GEN_6 = 2'h2 == s2_way ? sram_out_2 : _GEN_5; // @[Cache.scala 261:{18,18}]
  wire [127:0] sram_out_3 = sram_3_io_rdata;
  wire [127:0] _GEN_7 = 2'h3 == s2_way ? sram_out_3 : _GEN_6; // @[Cache.scala 261:{18,18}]
  wire  _GEN_39 = 6'h1 == s2_idx ? plru0_1 : plru0_0; // @[Cache.scala 268:{40,40}]
  wire  _GEN_40 = 6'h2 == s2_idx ? plru0_2 : _GEN_39; // @[Cache.scala 268:{40,40}]
  wire  _GEN_41 = 6'h3 == s2_idx ? plru0_3 : _GEN_40; // @[Cache.scala 268:{40,40}]
  wire  _GEN_42 = 6'h4 == s2_idx ? plru0_4 : _GEN_41; // @[Cache.scala 268:{40,40}]
  wire  _GEN_43 = 6'h5 == s2_idx ? plru0_5 : _GEN_42; // @[Cache.scala 268:{40,40}]
  wire  _GEN_44 = 6'h6 == s2_idx ? plru0_6 : _GEN_43; // @[Cache.scala 268:{40,40}]
  wire  _GEN_45 = 6'h7 == s2_idx ? plru0_7 : _GEN_44; // @[Cache.scala 268:{40,40}]
  wire  _GEN_46 = 6'h8 == s2_idx ? plru0_8 : _GEN_45; // @[Cache.scala 268:{40,40}]
  wire  _GEN_47 = 6'h9 == s2_idx ? plru0_9 : _GEN_46; // @[Cache.scala 268:{40,40}]
  wire  _GEN_48 = 6'ha == s2_idx ? plru0_10 : _GEN_47; // @[Cache.scala 268:{40,40}]
  wire  _GEN_49 = 6'hb == s2_idx ? plru0_11 : _GEN_48; // @[Cache.scala 268:{40,40}]
  wire  _GEN_50 = 6'hc == s2_idx ? plru0_12 : _GEN_49; // @[Cache.scala 268:{40,40}]
  wire  _GEN_51 = 6'hd == s2_idx ? plru0_13 : _GEN_50; // @[Cache.scala 268:{40,40}]
  wire  _GEN_52 = 6'he == s2_idx ? plru0_14 : _GEN_51; // @[Cache.scala 268:{40,40}]
  wire  _GEN_53 = 6'hf == s2_idx ? plru0_15 : _GEN_52; // @[Cache.scala 268:{40,40}]
  wire  _GEN_54 = 6'h10 == s2_idx ? plru0_16 : _GEN_53; // @[Cache.scala 268:{40,40}]
  wire  _GEN_55 = 6'h11 == s2_idx ? plru0_17 : _GEN_54; // @[Cache.scala 268:{40,40}]
  wire  _GEN_56 = 6'h12 == s2_idx ? plru0_18 : _GEN_55; // @[Cache.scala 268:{40,40}]
  wire  _GEN_57 = 6'h13 == s2_idx ? plru0_19 : _GEN_56; // @[Cache.scala 268:{40,40}]
  wire  _GEN_58 = 6'h14 == s2_idx ? plru0_20 : _GEN_57; // @[Cache.scala 268:{40,40}]
  wire  _GEN_59 = 6'h15 == s2_idx ? plru0_21 : _GEN_58; // @[Cache.scala 268:{40,40}]
  wire  _GEN_60 = 6'h16 == s2_idx ? plru0_22 : _GEN_59; // @[Cache.scala 268:{40,40}]
  wire  _GEN_61 = 6'h17 == s2_idx ? plru0_23 : _GEN_60; // @[Cache.scala 268:{40,40}]
  wire  _GEN_62 = 6'h18 == s2_idx ? plru0_24 : _GEN_61; // @[Cache.scala 268:{40,40}]
  wire  _GEN_63 = 6'h19 == s2_idx ? plru0_25 : _GEN_62; // @[Cache.scala 268:{40,40}]
  wire  _GEN_64 = 6'h1a == s2_idx ? plru0_26 : _GEN_63; // @[Cache.scala 268:{40,40}]
  wire  _GEN_65 = 6'h1b == s2_idx ? plru0_27 : _GEN_64; // @[Cache.scala 268:{40,40}]
  wire  _GEN_66 = 6'h1c == s2_idx ? plru0_28 : _GEN_65; // @[Cache.scala 268:{40,40}]
  wire  _GEN_67 = 6'h1d == s2_idx ? plru0_29 : _GEN_66; // @[Cache.scala 268:{40,40}]
  wire  _GEN_68 = 6'h1e == s2_idx ? plru0_30 : _GEN_67; // @[Cache.scala 268:{40,40}]
  wire  _GEN_69 = 6'h1f == s2_idx ? plru0_31 : _GEN_68; // @[Cache.scala 268:{40,40}]
  wire  _GEN_70 = 6'h20 == s2_idx ? plru0_32 : _GEN_69; // @[Cache.scala 268:{40,40}]
  wire  _GEN_71 = 6'h21 == s2_idx ? plru0_33 : _GEN_70; // @[Cache.scala 268:{40,40}]
  wire  _GEN_72 = 6'h22 == s2_idx ? plru0_34 : _GEN_71; // @[Cache.scala 268:{40,40}]
  wire  _GEN_73 = 6'h23 == s2_idx ? plru0_35 : _GEN_72; // @[Cache.scala 268:{40,40}]
  wire  _GEN_74 = 6'h24 == s2_idx ? plru0_36 : _GEN_73; // @[Cache.scala 268:{40,40}]
  wire  _GEN_75 = 6'h25 == s2_idx ? plru0_37 : _GEN_74; // @[Cache.scala 268:{40,40}]
  wire  _GEN_76 = 6'h26 == s2_idx ? plru0_38 : _GEN_75; // @[Cache.scala 268:{40,40}]
  wire  _GEN_77 = 6'h27 == s2_idx ? plru0_39 : _GEN_76; // @[Cache.scala 268:{40,40}]
  wire  _GEN_78 = 6'h28 == s2_idx ? plru0_40 : _GEN_77; // @[Cache.scala 268:{40,40}]
  wire  _GEN_79 = 6'h29 == s2_idx ? plru0_41 : _GEN_78; // @[Cache.scala 268:{40,40}]
  wire  _GEN_80 = 6'h2a == s2_idx ? plru0_42 : _GEN_79; // @[Cache.scala 268:{40,40}]
  wire  _GEN_81 = 6'h2b == s2_idx ? plru0_43 : _GEN_80; // @[Cache.scala 268:{40,40}]
  wire  _GEN_82 = 6'h2c == s2_idx ? plru0_44 : _GEN_81; // @[Cache.scala 268:{40,40}]
  wire  _GEN_83 = 6'h2d == s2_idx ? plru0_45 : _GEN_82; // @[Cache.scala 268:{40,40}]
  wire  _GEN_84 = 6'h2e == s2_idx ? plru0_46 : _GEN_83; // @[Cache.scala 268:{40,40}]
  wire  _GEN_85 = 6'h2f == s2_idx ? plru0_47 : _GEN_84; // @[Cache.scala 268:{40,40}]
  wire  _GEN_86 = 6'h30 == s2_idx ? plru0_48 : _GEN_85; // @[Cache.scala 268:{40,40}]
  wire  _GEN_87 = 6'h31 == s2_idx ? plru0_49 : _GEN_86; // @[Cache.scala 268:{40,40}]
  wire  _GEN_88 = 6'h32 == s2_idx ? plru0_50 : _GEN_87; // @[Cache.scala 268:{40,40}]
  wire  _GEN_89 = 6'h33 == s2_idx ? plru0_51 : _GEN_88; // @[Cache.scala 268:{40,40}]
  wire  _GEN_90 = 6'h34 == s2_idx ? plru0_52 : _GEN_89; // @[Cache.scala 268:{40,40}]
  wire  _GEN_91 = 6'h35 == s2_idx ? plru0_53 : _GEN_90; // @[Cache.scala 268:{40,40}]
  wire  _GEN_92 = 6'h36 == s2_idx ? plru0_54 : _GEN_91; // @[Cache.scala 268:{40,40}]
  wire  _GEN_93 = 6'h37 == s2_idx ? plru0_55 : _GEN_92; // @[Cache.scala 268:{40,40}]
  wire  _GEN_94 = 6'h38 == s2_idx ? plru0_56 : _GEN_93; // @[Cache.scala 268:{40,40}]
  wire  _GEN_95 = 6'h39 == s2_idx ? plru0_57 : _GEN_94; // @[Cache.scala 268:{40,40}]
  wire  _GEN_96 = 6'h3a == s2_idx ? plru0_58 : _GEN_95; // @[Cache.scala 268:{40,40}]
  wire  _GEN_97 = 6'h3b == s2_idx ? plru0_59 : _GEN_96; // @[Cache.scala 268:{40,40}]
  wire  _GEN_98 = 6'h3c == s2_idx ? plru0_60 : _GEN_97; // @[Cache.scala 268:{40,40}]
  wire  _GEN_99 = 6'h3d == s2_idx ? plru0_61 : _GEN_98; // @[Cache.scala 268:{40,40}]
  wire  _GEN_100 = 6'h3e == s2_idx ? plru0_62 : _GEN_99; // @[Cache.scala 268:{40,40}]
  wire  _GEN_101 = 6'h3f == s2_idx ? plru0_63 : _GEN_100; // @[Cache.scala 268:{40,40}]
  wire  _GEN_103 = 6'h1 == s2_idx ? plru1_1 : plru1_0; // @[Cache.scala 268:{25,25}]
  wire  _GEN_104 = 6'h2 == s2_idx ? plru1_2 : _GEN_103; // @[Cache.scala 268:{25,25}]
  wire  _GEN_105 = 6'h3 == s2_idx ? plru1_3 : _GEN_104; // @[Cache.scala 268:{25,25}]
  wire  _GEN_106 = 6'h4 == s2_idx ? plru1_4 : _GEN_105; // @[Cache.scala 268:{25,25}]
  wire  _GEN_107 = 6'h5 == s2_idx ? plru1_5 : _GEN_106; // @[Cache.scala 268:{25,25}]
  wire  _GEN_108 = 6'h6 == s2_idx ? plru1_6 : _GEN_107; // @[Cache.scala 268:{25,25}]
  wire  _GEN_109 = 6'h7 == s2_idx ? plru1_7 : _GEN_108; // @[Cache.scala 268:{25,25}]
  wire  _GEN_110 = 6'h8 == s2_idx ? plru1_8 : _GEN_109; // @[Cache.scala 268:{25,25}]
  wire  _GEN_111 = 6'h9 == s2_idx ? plru1_9 : _GEN_110; // @[Cache.scala 268:{25,25}]
  wire  _GEN_112 = 6'ha == s2_idx ? plru1_10 : _GEN_111; // @[Cache.scala 268:{25,25}]
  wire  _GEN_113 = 6'hb == s2_idx ? plru1_11 : _GEN_112; // @[Cache.scala 268:{25,25}]
  wire  _GEN_114 = 6'hc == s2_idx ? plru1_12 : _GEN_113; // @[Cache.scala 268:{25,25}]
  wire  _GEN_115 = 6'hd == s2_idx ? plru1_13 : _GEN_114; // @[Cache.scala 268:{25,25}]
  wire  _GEN_116 = 6'he == s2_idx ? plru1_14 : _GEN_115; // @[Cache.scala 268:{25,25}]
  wire  _GEN_117 = 6'hf == s2_idx ? plru1_15 : _GEN_116; // @[Cache.scala 268:{25,25}]
  wire  _GEN_118 = 6'h10 == s2_idx ? plru1_16 : _GEN_117; // @[Cache.scala 268:{25,25}]
  wire  _GEN_119 = 6'h11 == s2_idx ? plru1_17 : _GEN_118; // @[Cache.scala 268:{25,25}]
  wire  _GEN_120 = 6'h12 == s2_idx ? plru1_18 : _GEN_119; // @[Cache.scala 268:{25,25}]
  wire  _GEN_121 = 6'h13 == s2_idx ? plru1_19 : _GEN_120; // @[Cache.scala 268:{25,25}]
  wire  _GEN_122 = 6'h14 == s2_idx ? plru1_20 : _GEN_121; // @[Cache.scala 268:{25,25}]
  wire  _GEN_123 = 6'h15 == s2_idx ? plru1_21 : _GEN_122; // @[Cache.scala 268:{25,25}]
  wire  _GEN_124 = 6'h16 == s2_idx ? plru1_22 : _GEN_123; // @[Cache.scala 268:{25,25}]
  wire  _GEN_125 = 6'h17 == s2_idx ? plru1_23 : _GEN_124; // @[Cache.scala 268:{25,25}]
  wire  _GEN_126 = 6'h18 == s2_idx ? plru1_24 : _GEN_125; // @[Cache.scala 268:{25,25}]
  wire  _GEN_127 = 6'h19 == s2_idx ? plru1_25 : _GEN_126; // @[Cache.scala 268:{25,25}]
  wire  _GEN_128 = 6'h1a == s2_idx ? plru1_26 : _GEN_127; // @[Cache.scala 268:{25,25}]
  wire  _GEN_129 = 6'h1b == s2_idx ? plru1_27 : _GEN_128; // @[Cache.scala 268:{25,25}]
  wire  _GEN_130 = 6'h1c == s2_idx ? plru1_28 : _GEN_129; // @[Cache.scala 268:{25,25}]
  wire  _GEN_131 = 6'h1d == s2_idx ? plru1_29 : _GEN_130; // @[Cache.scala 268:{25,25}]
  wire  _GEN_132 = 6'h1e == s2_idx ? plru1_30 : _GEN_131; // @[Cache.scala 268:{25,25}]
  wire  _GEN_133 = 6'h1f == s2_idx ? plru1_31 : _GEN_132; // @[Cache.scala 268:{25,25}]
  wire  _GEN_134 = 6'h20 == s2_idx ? plru1_32 : _GEN_133; // @[Cache.scala 268:{25,25}]
  wire  _GEN_135 = 6'h21 == s2_idx ? plru1_33 : _GEN_134; // @[Cache.scala 268:{25,25}]
  wire  _GEN_136 = 6'h22 == s2_idx ? plru1_34 : _GEN_135; // @[Cache.scala 268:{25,25}]
  wire  _GEN_137 = 6'h23 == s2_idx ? plru1_35 : _GEN_136; // @[Cache.scala 268:{25,25}]
  wire  _GEN_138 = 6'h24 == s2_idx ? plru1_36 : _GEN_137; // @[Cache.scala 268:{25,25}]
  wire  _GEN_139 = 6'h25 == s2_idx ? plru1_37 : _GEN_138; // @[Cache.scala 268:{25,25}]
  wire  _GEN_140 = 6'h26 == s2_idx ? plru1_38 : _GEN_139; // @[Cache.scala 268:{25,25}]
  wire  _GEN_141 = 6'h27 == s2_idx ? plru1_39 : _GEN_140; // @[Cache.scala 268:{25,25}]
  wire  _GEN_142 = 6'h28 == s2_idx ? plru1_40 : _GEN_141; // @[Cache.scala 268:{25,25}]
  wire  _GEN_143 = 6'h29 == s2_idx ? plru1_41 : _GEN_142; // @[Cache.scala 268:{25,25}]
  wire  _GEN_144 = 6'h2a == s2_idx ? plru1_42 : _GEN_143; // @[Cache.scala 268:{25,25}]
  wire  _GEN_145 = 6'h2b == s2_idx ? plru1_43 : _GEN_144; // @[Cache.scala 268:{25,25}]
  wire  _GEN_146 = 6'h2c == s2_idx ? plru1_44 : _GEN_145; // @[Cache.scala 268:{25,25}]
  wire  _GEN_147 = 6'h2d == s2_idx ? plru1_45 : _GEN_146; // @[Cache.scala 268:{25,25}]
  wire  _GEN_148 = 6'h2e == s2_idx ? plru1_46 : _GEN_147; // @[Cache.scala 268:{25,25}]
  wire  _GEN_149 = 6'h2f == s2_idx ? plru1_47 : _GEN_148; // @[Cache.scala 268:{25,25}]
  wire  _GEN_150 = 6'h30 == s2_idx ? plru1_48 : _GEN_149; // @[Cache.scala 268:{25,25}]
  wire  _GEN_151 = 6'h31 == s2_idx ? plru1_49 : _GEN_150; // @[Cache.scala 268:{25,25}]
  wire  _GEN_152 = 6'h32 == s2_idx ? plru1_50 : _GEN_151; // @[Cache.scala 268:{25,25}]
  wire  _GEN_153 = 6'h33 == s2_idx ? plru1_51 : _GEN_152; // @[Cache.scala 268:{25,25}]
  wire  _GEN_154 = 6'h34 == s2_idx ? plru1_52 : _GEN_153; // @[Cache.scala 268:{25,25}]
  wire  _GEN_155 = 6'h35 == s2_idx ? plru1_53 : _GEN_154; // @[Cache.scala 268:{25,25}]
  wire  _GEN_156 = 6'h36 == s2_idx ? plru1_54 : _GEN_155; // @[Cache.scala 268:{25,25}]
  wire  _GEN_157 = 6'h37 == s2_idx ? plru1_55 : _GEN_156; // @[Cache.scala 268:{25,25}]
  wire  _GEN_158 = 6'h38 == s2_idx ? plru1_56 : _GEN_157; // @[Cache.scala 268:{25,25}]
  wire  _GEN_159 = 6'h39 == s2_idx ? plru1_57 : _GEN_158; // @[Cache.scala 268:{25,25}]
  wire  _GEN_160 = 6'h3a == s2_idx ? plru1_58 : _GEN_159; // @[Cache.scala 268:{25,25}]
  wire  _GEN_161 = 6'h3b == s2_idx ? plru1_59 : _GEN_160; // @[Cache.scala 268:{25,25}]
  wire  _GEN_162 = 6'h3c == s2_idx ? plru1_60 : _GEN_161; // @[Cache.scala 268:{25,25}]
  wire  _GEN_163 = 6'h3d == s2_idx ? plru1_61 : _GEN_162; // @[Cache.scala 268:{25,25}]
  wire  _GEN_164 = 6'h3e == s2_idx ? plru1_62 : _GEN_163; // @[Cache.scala 268:{25,25}]
  wire  _GEN_165 = 6'h3f == s2_idx ? plru1_63 : _GEN_164; // @[Cache.scala 268:{25,25}]
  wire  _GEN_167 = 6'h1 == s2_idx ? plru2_1 : plru2_0; // @[Cache.scala 268:{25,25}]
  wire  _GEN_168 = 6'h2 == s2_idx ? plru2_2 : _GEN_167; // @[Cache.scala 268:{25,25}]
  wire  _GEN_169 = 6'h3 == s2_idx ? plru2_3 : _GEN_168; // @[Cache.scala 268:{25,25}]
  wire  _GEN_170 = 6'h4 == s2_idx ? plru2_4 : _GEN_169; // @[Cache.scala 268:{25,25}]
  wire  _GEN_171 = 6'h5 == s2_idx ? plru2_5 : _GEN_170; // @[Cache.scala 268:{25,25}]
  wire  _GEN_172 = 6'h6 == s2_idx ? plru2_6 : _GEN_171; // @[Cache.scala 268:{25,25}]
  wire  _GEN_173 = 6'h7 == s2_idx ? plru2_7 : _GEN_172; // @[Cache.scala 268:{25,25}]
  wire  _GEN_174 = 6'h8 == s2_idx ? plru2_8 : _GEN_173; // @[Cache.scala 268:{25,25}]
  wire  _GEN_175 = 6'h9 == s2_idx ? plru2_9 : _GEN_174; // @[Cache.scala 268:{25,25}]
  wire  _GEN_176 = 6'ha == s2_idx ? plru2_10 : _GEN_175; // @[Cache.scala 268:{25,25}]
  wire  _GEN_177 = 6'hb == s2_idx ? plru2_11 : _GEN_176; // @[Cache.scala 268:{25,25}]
  wire  _GEN_178 = 6'hc == s2_idx ? plru2_12 : _GEN_177; // @[Cache.scala 268:{25,25}]
  wire  _GEN_179 = 6'hd == s2_idx ? plru2_13 : _GEN_178; // @[Cache.scala 268:{25,25}]
  wire  _GEN_180 = 6'he == s2_idx ? plru2_14 : _GEN_179; // @[Cache.scala 268:{25,25}]
  wire  _GEN_181 = 6'hf == s2_idx ? plru2_15 : _GEN_180; // @[Cache.scala 268:{25,25}]
  wire  _GEN_182 = 6'h10 == s2_idx ? plru2_16 : _GEN_181; // @[Cache.scala 268:{25,25}]
  wire  _GEN_183 = 6'h11 == s2_idx ? plru2_17 : _GEN_182; // @[Cache.scala 268:{25,25}]
  wire  _GEN_184 = 6'h12 == s2_idx ? plru2_18 : _GEN_183; // @[Cache.scala 268:{25,25}]
  wire  _GEN_185 = 6'h13 == s2_idx ? plru2_19 : _GEN_184; // @[Cache.scala 268:{25,25}]
  wire  _GEN_186 = 6'h14 == s2_idx ? plru2_20 : _GEN_185; // @[Cache.scala 268:{25,25}]
  wire  _GEN_187 = 6'h15 == s2_idx ? plru2_21 : _GEN_186; // @[Cache.scala 268:{25,25}]
  wire  _GEN_188 = 6'h16 == s2_idx ? plru2_22 : _GEN_187; // @[Cache.scala 268:{25,25}]
  wire  _GEN_189 = 6'h17 == s2_idx ? plru2_23 : _GEN_188; // @[Cache.scala 268:{25,25}]
  wire  _GEN_190 = 6'h18 == s2_idx ? plru2_24 : _GEN_189; // @[Cache.scala 268:{25,25}]
  wire  _GEN_191 = 6'h19 == s2_idx ? plru2_25 : _GEN_190; // @[Cache.scala 268:{25,25}]
  wire  _GEN_192 = 6'h1a == s2_idx ? plru2_26 : _GEN_191; // @[Cache.scala 268:{25,25}]
  wire  _GEN_193 = 6'h1b == s2_idx ? plru2_27 : _GEN_192; // @[Cache.scala 268:{25,25}]
  wire  _GEN_194 = 6'h1c == s2_idx ? plru2_28 : _GEN_193; // @[Cache.scala 268:{25,25}]
  wire  _GEN_195 = 6'h1d == s2_idx ? plru2_29 : _GEN_194; // @[Cache.scala 268:{25,25}]
  wire  _GEN_196 = 6'h1e == s2_idx ? plru2_30 : _GEN_195; // @[Cache.scala 268:{25,25}]
  wire  _GEN_197 = 6'h1f == s2_idx ? plru2_31 : _GEN_196; // @[Cache.scala 268:{25,25}]
  wire  _GEN_198 = 6'h20 == s2_idx ? plru2_32 : _GEN_197; // @[Cache.scala 268:{25,25}]
  wire  _GEN_199 = 6'h21 == s2_idx ? plru2_33 : _GEN_198; // @[Cache.scala 268:{25,25}]
  wire  _GEN_200 = 6'h22 == s2_idx ? plru2_34 : _GEN_199; // @[Cache.scala 268:{25,25}]
  wire  _GEN_201 = 6'h23 == s2_idx ? plru2_35 : _GEN_200; // @[Cache.scala 268:{25,25}]
  wire  _GEN_202 = 6'h24 == s2_idx ? plru2_36 : _GEN_201; // @[Cache.scala 268:{25,25}]
  wire  _GEN_203 = 6'h25 == s2_idx ? plru2_37 : _GEN_202; // @[Cache.scala 268:{25,25}]
  wire  _GEN_204 = 6'h26 == s2_idx ? plru2_38 : _GEN_203; // @[Cache.scala 268:{25,25}]
  wire  _GEN_205 = 6'h27 == s2_idx ? plru2_39 : _GEN_204; // @[Cache.scala 268:{25,25}]
  wire  _GEN_206 = 6'h28 == s2_idx ? plru2_40 : _GEN_205; // @[Cache.scala 268:{25,25}]
  wire  _GEN_207 = 6'h29 == s2_idx ? plru2_41 : _GEN_206; // @[Cache.scala 268:{25,25}]
  wire  _GEN_208 = 6'h2a == s2_idx ? plru2_42 : _GEN_207; // @[Cache.scala 268:{25,25}]
  wire  _GEN_209 = 6'h2b == s2_idx ? plru2_43 : _GEN_208; // @[Cache.scala 268:{25,25}]
  wire  _GEN_210 = 6'h2c == s2_idx ? plru2_44 : _GEN_209; // @[Cache.scala 268:{25,25}]
  wire  _GEN_211 = 6'h2d == s2_idx ? plru2_45 : _GEN_210; // @[Cache.scala 268:{25,25}]
  wire  _GEN_212 = 6'h2e == s2_idx ? plru2_46 : _GEN_211; // @[Cache.scala 268:{25,25}]
  wire  _GEN_213 = 6'h2f == s2_idx ? plru2_47 : _GEN_212; // @[Cache.scala 268:{25,25}]
  wire  _GEN_214 = 6'h30 == s2_idx ? plru2_48 : _GEN_213; // @[Cache.scala 268:{25,25}]
  wire  _GEN_215 = 6'h31 == s2_idx ? plru2_49 : _GEN_214; // @[Cache.scala 268:{25,25}]
  wire  _GEN_216 = 6'h32 == s2_idx ? plru2_50 : _GEN_215; // @[Cache.scala 268:{25,25}]
  wire  _GEN_217 = 6'h33 == s2_idx ? plru2_51 : _GEN_216; // @[Cache.scala 268:{25,25}]
  wire  _GEN_218 = 6'h34 == s2_idx ? plru2_52 : _GEN_217; // @[Cache.scala 268:{25,25}]
  wire  _GEN_219 = 6'h35 == s2_idx ? plru2_53 : _GEN_218; // @[Cache.scala 268:{25,25}]
  wire  _GEN_220 = 6'h36 == s2_idx ? plru2_54 : _GEN_219; // @[Cache.scala 268:{25,25}]
  wire  _GEN_221 = 6'h37 == s2_idx ? plru2_55 : _GEN_220; // @[Cache.scala 268:{25,25}]
  wire  _GEN_222 = 6'h38 == s2_idx ? plru2_56 : _GEN_221; // @[Cache.scala 268:{25,25}]
  wire  _GEN_223 = 6'h39 == s2_idx ? plru2_57 : _GEN_222; // @[Cache.scala 268:{25,25}]
  wire  _GEN_224 = 6'h3a == s2_idx ? plru2_58 : _GEN_223; // @[Cache.scala 268:{25,25}]
  wire  _GEN_225 = 6'h3b == s2_idx ? plru2_59 : _GEN_224; // @[Cache.scala 268:{25,25}]
  wire  _GEN_226 = 6'h3c == s2_idx ? plru2_60 : _GEN_225; // @[Cache.scala 268:{25,25}]
  wire  _GEN_227 = 6'h3d == s2_idx ? plru2_61 : _GEN_226; // @[Cache.scala 268:{25,25}]
  wire  _GEN_228 = 6'h3e == s2_idx ? plru2_62 : _GEN_227; // @[Cache.scala 268:{25,25}]
  wire  _GEN_229 = 6'h3f == s2_idx ? plru2_63 : _GEN_228; // @[Cache.scala 268:{25,25}]
  wire  _T_16 = ~_GEN_101 ? _GEN_165 : _GEN_229; // @[Cache.scala 268:25]
  wire [1:0] replace_way = {_GEN_101,_T_16}; // @[Cat.scala 30:58]
  wire  _GEN_9 = 2'h1 == replace_way ? REG_5 : REG_4; // @[Cache.scala 262:{18,18}]
  wire  _GEN_10 = 2'h2 == replace_way ? REG_6 : _GEN_9; // @[Cache.scala 262:{18,18}]
  wire [20:0] _GEN_13 = 2'h1 == replace_way ? tag_out_1 : tag_out_0; // @[Cache.scala 263:{18,18}]
  wire [20:0] _GEN_14 = 2'h2 == replace_way ? tag_out_2 : _GEN_13; // @[Cache.scala 263:{18,18}]
  wire [127:0] _GEN_17 = 2'h1 == replace_way ? sram_out_1 : sram_out_0; // @[Cache.scala 264:{18,18}]
  wire [127:0] _GEN_18 = 2'h2 == replace_way ? sram_out_2 : _GEN_17; // @[Cache.scala 264:{18,18}]
  reg [63:0] wdata1; // @[Cache.scala 270:23]
  reg [63:0] wdata2; // @[Cache.scala 271:23]
  reg  REG_10; // @[Cache.scala 320:20]
  wire [63:0] _T_36 = s2_offs ? _GEN_7[127:64] : _GEN_7[63:0]; // @[Cache.scala 321:34]
  wire [63:0] _T_40 = s2_offs ? s2_reg_rdata[127:64] : s2_reg_rdata[63:0]; // @[Cache.scala 323:34]
  wire [63:0] _GEN_230 = REG_10 ? _T_36 : _T_40; // @[Cache.scala 320:37 321:28 323:28]
  reg  REG_11; // @[Cache.scala 325:20]
  wire  _T_42 = ~s2_way[1]; // @[Cache.scala 136:19]
  wire  _GEN_231 = 6'h0 == s2_idx ? ~s2_way[1] : plru0_0; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_232 = 6'h1 == s2_idx ? ~s2_way[1] : plru0_1; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_233 = 6'h2 == s2_idx ? ~s2_way[1] : plru0_2; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_234 = 6'h3 == s2_idx ? ~s2_way[1] : plru0_3; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_235 = 6'h4 == s2_idx ? ~s2_way[1] : plru0_4; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_236 = 6'h5 == s2_idx ? ~s2_way[1] : plru0_5; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_237 = 6'h6 == s2_idx ? ~s2_way[1] : plru0_6; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_238 = 6'h7 == s2_idx ? ~s2_way[1] : plru0_7; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_239 = 6'h8 == s2_idx ? ~s2_way[1] : plru0_8; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_240 = 6'h9 == s2_idx ? ~s2_way[1] : plru0_9; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_241 = 6'ha == s2_idx ? ~s2_way[1] : plru0_10; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_242 = 6'hb == s2_idx ? ~s2_way[1] : plru0_11; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_243 = 6'hc == s2_idx ? ~s2_way[1] : plru0_12; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_244 = 6'hd == s2_idx ? ~s2_way[1] : plru0_13; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_245 = 6'he == s2_idx ? ~s2_way[1] : plru0_14; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_246 = 6'hf == s2_idx ? ~s2_way[1] : plru0_15; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_247 = 6'h10 == s2_idx ? ~s2_way[1] : plru0_16; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_248 = 6'h11 == s2_idx ? ~s2_way[1] : plru0_17; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_249 = 6'h12 == s2_idx ? ~s2_way[1] : plru0_18; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_250 = 6'h13 == s2_idx ? ~s2_way[1] : plru0_19; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_251 = 6'h14 == s2_idx ? ~s2_way[1] : plru0_20; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_252 = 6'h15 == s2_idx ? ~s2_way[1] : plru0_21; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_253 = 6'h16 == s2_idx ? ~s2_way[1] : plru0_22; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_254 = 6'h17 == s2_idx ? ~s2_way[1] : plru0_23; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_255 = 6'h18 == s2_idx ? ~s2_way[1] : plru0_24; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_256 = 6'h19 == s2_idx ? ~s2_way[1] : plru0_25; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_257 = 6'h1a == s2_idx ? ~s2_way[1] : plru0_26; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_258 = 6'h1b == s2_idx ? ~s2_way[1] : plru0_27; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_259 = 6'h1c == s2_idx ? ~s2_way[1] : plru0_28; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_260 = 6'h1d == s2_idx ? ~s2_way[1] : plru0_29; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_261 = 6'h1e == s2_idx ? ~s2_way[1] : plru0_30; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_262 = 6'h1f == s2_idx ? ~s2_way[1] : plru0_31; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_263 = 6'h20 == s2_idx ? ~s2_way[1] : plru0_32; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_264 = 6'h21 == s2_idx ? ~s2_way[1] : plru0_33; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_265 = 6'h22 == s2_idx ? ~s2_way[1] : plru0_34; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_266 = 6'h23 == s2_idx ? ~s2_way[1] : plru0_35; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_267 = 6'h24 == s2_idx ? ~s2_way[1] : plru0_36; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_268 = 6'h25 == s2_idx ? ~s2_way[1] : plru0_37; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_269 = 6'h26 == s2_idx ? ~s2_way[1] : plru0_38; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_270 = 6'h27 == s2_idx ? ~s2_way[1] : plru0_39; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_271 = 6'h28 == s2_idx ? ~s2_way[1] : plru0_40; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_272 = 6'h29 == s2_idx ? ~s2_way[1] : plru0_41; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_273 = 6'h2a == s2_idx ? ~s2_way[1] : plru0_42; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_274 = 6'h2b == s2_idx ? ~s2_way[1] : plru0_43; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_275 = 6'h2c == s2_idx ? ~s2_way[1] : plru0_44; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_276 = 6'h2d == s2_idx ? ~s2_way[1] : plru0_45; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_277 = 6'h2e == s2_idx ? ~s2_way[1] : plru0_46; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_278 = 6'h2f == s2_idx ? ~s2_way[1] : plru0_47; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_279 = 6'h30 == s2_idx ? ~s2_way[1] : plru0_48; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_280 = 6'h31 == s2_idx ? ~s2_way[1] : plru0_49; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_281 = 6'h32 == s2_idx ? ~s2_way[1] : plru0_50; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_282 = 6'h33 == s2_idx ? ~s2_way[1] : plru0_51; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_283 = 6'h34 == s2_idx ? ~s2_way[1] : plru0_52; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_284 = 6'h35 == s2_idx ? ~s2_way[1] : plru0_53; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_285 = 6'h36 == s2_idx ? ~s2_way[1] : plru0_54; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_286 = 6'h37 == s2_idx ? ~s2_way[1] : plru0_55; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_287 = 6'h38 == s2_idx ? ~s2_way[1] : plru0_56; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_288 = 6'h39 == s2_idx ? ~s2_way[1] : plru0_57; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_289 = 6'h3a == s2_idx ? ~s2_way[1] : plru0_58; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_290 = 6'h3b == s2_idx ? ~s2_way[1] : plru0_59; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_291 = 6'h3c == s2_idx ? ~s2_way[1] : plru0_60; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_292 = 6'h3d == s2_idx ? ~s2_way[1] : plru0_61; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_293 = 6'h3e == s2_idx ? ~s2_way[1] : plru0_62; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_294 = 6'h3f == s2_idx ? ~s2_way[1] : plru0_63; // @[Cache.scala 136:{16,16} 129:22]
  wire  _T_46 = ~s2_way[0]; // @[Cache.scala 138:21]
  wire  _GEN_295 = 6'h0 == s2_idx ? ~s2_way[0] : plru1_0; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_296 = 6'h1 == s2_idx ? ~s2_way[0] : plru1_1; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_297 = 6'h2 == s2_idx ? ~s2_way[0] : plru1_2; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_298 = 6'h3 == s2_idx ? ~s2_way[0] : plru1_3; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_299 = 6'h4 == s2_idx ? ~s2_way[0] : plru1_4; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_300 = 6'h5 == s2_idx ? ~s2_way[0] : plru1_5; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_301 = 6'h6 == s2_idx ? ~s2_way[0] : plru1_6; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_302 = 6'h7 == s2_idx ? ~s2_way[0] : plru1_7; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_303 = 6'h8 == s2_idx ? ~s2_way[0] : plru1_8; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_304 = 6'h9 == s2_idx ? ~s2_way[0] : plru1_9; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_305 = 6'ha == s2_idx ? ~s2_way[0] : plru1_10; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_306 = 6'hb == s2_idx ? ~s2_way[0] : plru1_11; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_307 = 6'hc == s2_idx ? ~s2_way[0] : plru1_12; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_308 = 6'hd == s2_idx ? ~s2_way[0] : plru1_13; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_309 = 6'he == s2_idx ? ~s2_way[0] : plru1_14; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_310 = 6'hf == s2_idx ? ~s2_way[0] : plru1_15; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_311 = 6'h10 == s2_idx ? ~s2_way[0] : plru1_16; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_312 = 6'h11 == s2_idx ? ~s2_way[0] : plru1_17; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_313 = 6'h12 == s2_idx ? ~s2_way[0] : plru1_18; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_314 = 6'h13 == s2_idx ? ~s2_way[0] : plru1_19; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_315 = 6'h14 == s2_idx ? ~s2_way[0] : plru1_20; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_316 = 6'h15 == s2_idx ? ~s2_way[0] : plru1_21; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_317 = 6'h16 == s2_idx ? ~s2_way[0] : plru1_22; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_318 = 6'h17 == s2_idx ? ~s2_way[0] : plru1_23; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_319 = 6'h18 == s2_idx ? ~s2_way[0] : plru1_24; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_320 = 6'h19 == s2_idx ? ~s2_way[0] : plru1_25; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_321 = 6'h1a == s2_idx ? ~s2_way[0] : plru1_26; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_322 = 6'h1b == s2_idx ? ~s2_way[0] : plru1_27; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_323 = 6'h1c == s2_idx ? ~s2_way[0] : plru1_28; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_324 = 6'h1d == s2_idx ? ~s2_way[0] : plru1_29; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_325 = 6'h1e == s2_idx ? ~s2_way[0] : plru1_30; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_326 = 6'h1f == s2_idx ? ~s2_way[0] : plru1_31; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_327 = 6'h20 == s2_idx ? ~s2_way[0] : plru1_32; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_328 = 6'h21 == s2_idx ? ~s2_way[0] : plru1_33; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_329 = 6'h22 == s2_idx ? ~s2_way[0] : plru1_34; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_330 = 6'h23 == s2_idx ? ~s2_way[0] : plru1_35; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_331 = 6'h24 == s2_idx ? ~s2_way[0] : plru1_36; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_332 = 6'h25 == s2_idx ? ~s2_way[0] : plru1_37; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_333 = 6'h26 == s2_idx ? ~s2_way[0] : plru1_38; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_334 = 6'h27 == s2_idx ? ~s2_way[0] : plru1_39; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_335 = 6'h28 == s2_idx ? ~s2_way[0] : plru1_40; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_336 = 6'h29 == s2_idx ? ~s2_way[0] : plru1_41; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_337 = 6'h2a == s2_idx ? ~s2_way[0] : plru1_42; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_338 = 6'h2b == s2_idx ? ~s2_way[0] : plru1_43; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_339 = 6'h2c == s2_idx ? ~s2_way[0] : plru1_44; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_340 = 6'h2d == s2_idx ? ~s2_way[0] : plru1_45; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_341 = 6'h2e == s2_idx ? ~s2_way[0] : plru1_46; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_342 = 6'h2f == s2_idx ? ~s2_way[0] : plru1_47; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_343 = 6'h30 == s2_idx ? ~s2_way[0] : plru1_48; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_344 = 6'h31 == s2_idx ? ~s2_way[0] : plru1_49; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_345 = 6'h32 == s2_idx ? ~s2_way[0] : plru1_50; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_346 = 6'h33 == s2_idx ? ~s2_way[0] : plru1_51; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_347 = 6'h34 == s2_idx ? ~s2_way[0] : plru1_52; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_348 = 6'h35 == s2_idx ? ~s2_way[0] : plru1_53; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_349 = 6'h36 == s2_idx ? ~s2_way[0] : plru1_54; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_350 = 6'h37 == s2_idx ? ~s2_way[0] : plru1_55; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_351 = 6'h38 == s2_idx ? ~s2_way[0] : plru1_56; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_352 = 6'h39 == s2_idx ? ~s2_way[0] : plru1_57; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_353 = 6'h3a == s2_idx ? ~s2_way[0] : plru1_58; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_354 = 6'h3b == s2_idx ? ~s2_way[0] : plru1_59; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_355 = 6'h3c == s2_idx ? ~s2_way[0] : plru1_60; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_356 = 6'h3d == s2_idx ? ~s2_way[0] : plru1_61; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_357 = 6'h3e == s2_idx ? ~s2_way[0] : plru1_62; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_358 = 6'h3f == s2_idx ? ~s2_way[0] : plru1_63; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_359 = 6'h0 == s2_idx ? _T_46 : plru2_0; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_360 = 6'h1 == s2_idx ? _T_46 : plru2_1; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_361 = 6'h2 == s2_idx ? _T_46 : plru2_2; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_362 = 6'h3 == s2_idx ? _T_46 : plru2_3; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_363 = 6'h4 == s2_idx ? _T_46 : plru2_4; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_364 = 6'h5 == s2_idx ? _T_46 : plru2_5; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_365 = 6'h6 == s2_idx ? _T_46 : plru2_6; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_366 = 6'h7 == s2_idx ? _T_46 : plru2_7; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_367 = 6'h8 == s2_idx ? _T_46 : plru2_8; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_368 = 6'h9 == s2_idx ? _T_46 : plru2_9; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_369 = 6'ha == s2_idx ? _T_46 : plru2_10; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_370 = 6'hb == s2_idx ? _T_46 : plru2_11; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_371 = 6'hc == s2_idx ? _T_46 : plru2_12; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_372 = 6'hd == s2_idx ? _T_46 : plru2_13; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_373 = 6'he == s2_idx ? _T_46 : plru2_14; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_374 = 6'hf == s2_idx ? _T_46 : plru2_15; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_375 = 6'h10 == s2_idx ? _T_46 : plru2_16; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_376 = 6'h11 == s2_idx ? _T_46 : plru2_17; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_377 = 6'h12 == s2_idx ? _T_46 : plru2_18; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_378 = 6'h13 == s2_idx ? _T_46 : plru2_19; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_379 = 6'h14 == s2_idx ? _T_46 : plru2_20; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_380 = 6'h15 == s2_idx ? _T_46 : plru2_21; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_381 = 6'h16 == s2_idx ? _T_46 : plru2_22; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_382 = 6'h17 == s2_idx ? _T_46 : plru2_23; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_383 = 6'h18 == s2_idx ? _T_46 : plru2_24; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_384 = 6'h19 == s2_idx ? _T_46 : plru2_25; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_385 = 6'h1a == s2_idx ? _T_46 : plru2_26; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_386 = 6'h1b == s2_idx ? _T_46 : plru2_27; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_387 = 6'h1c == s2_idx ? _T_46 : plru2_28; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_388 = 6'h1d == s2_idx ? _T_46 : plru2_29; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_389 = 6'h1e == s2_idx ? _T_46 : plru2_30; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_390 = 6'h1f == s2_idx ? _T_46 : plru2_31; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_391 = 6'h20 == s2_idx ? _T_46 : plru2_32; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_392 = 6'h21 == s2_idx ? _T_46 : plru2_33; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_393 = 6'h22 == s2_idx ? _T_46 : plru2_34; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_394 = 6'h23 == s2_idx ? _T_46 : plru2_35; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_395 = 6'h24 == s2_idx ? _T_46 : plru2_36; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_396 = 6'h25 == s2_idx ? _T_46 : plru2_37; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_397 = 6'h26 == s2_idx ? _T_46 : plru2_38; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_398 = 6'h27 == s2_idx ? _T_46 : plru2_39; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_399 = 6'h28 == s2_idx ? _T_46 : plru2_40; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_400 = 6'h29 == s2_idx ? _T_46 : plru2_41; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_401 = 6'h2a == s2_idx ? _T_46 : plru2_42; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_402 = 6'h2b == s2_idx ? _T_46 : plru2_43; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_403 = 6'h2c == s2_idx ? _T_46 : plru2_44; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_404 = 6'h2d == s2_idx ? _T_46 : plru2_45; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_405 = 6'h2e == s2_idx ? _T_46 : plru2_46; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_406 = 6'h2f == s2_idx ? _T_46 : plru2_47; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_407 = 6'h30 == s2_idx ? _T_46 : plru2_48; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_408 = 6'h31 == s2_idx ? _T_46 : plru2_49; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_409 = 6'h32 == s2_idx ? _T_46 : plru2_50; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_410 = 6'h33 == s2_idx ? _T_46 : plru2_51; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_411 = 6'h34 == s2_idx ? _T_46 : plru2_52; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_412 = 6'h35 == s2_idx ? _T_46 : plru2_53; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_413 = 6'h36 == s2_idx ? _T_46 : plru2_54; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_414 = 6'h37 == s2_idx ? _T_46 : plru2_55; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_415 = 6'h38 == s2_idx ? _T_46 : plru2_56; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_416 = 6'h39 == s2_idx ? _T_46 : plru2_57; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_417 = 6'h3a == s2_idx ? _T_46 : plru2_58; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_418 = 6'h3b == s2_idx ? _T_46 : plru2_59; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_419 = 6'h3c == s2_idx ? _T_46 : plru2_60; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_420 = 6'h3d == s2_idx ? _T_46 : plru2_61; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_421 = 6'h3e == s2_idx ? _T_46 : plru2_62; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_422 = 6'h3f == s2_idx ? _T_46 : plru2_63; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_423 = _T_42 ? _GEN_295 : plru1_0; // @[Cache.scala 131:22 137:27]
  wire  _GEN_424 = _T_42 ? _GEN_296 : plru1_1; // @[Cache.scala 131:22 137:27]
  wire  _GEN_425 = _T_42 ? _GEN_297 : plru1_2; // @[Cache.scala 131:22 137:27]
  wire  _GEN_426 = _T_42 ? _GEN_298 : plru1_3; // @[Cache.scala 131:22 137:27]
  wire  _GEN_427 = _T_42 ? _GEN_299 : plru1_4; // @[Cache.scala 131:22 137:27]
  wire  _GEN_428 = _T_42 ? _GEN_300 : plru1_5; // @[Cache.scala 131:22 137:27]
  wire  _GEN_429 = _T_42 ? _GEN_301 : plru1_6; // @[Cache.scala 131:22 137:27]
  wire  _GEN_430 = _T_42 ? _GEN_302 : plru1_7; // @[Cache.scala 131:22 137:27]
  wire  _GEN_431 = _T_42 ? _GEN_303 : plru1_8; // @[Cache.scala 131:22 137:27]
  wire  _GEN_432 = _T_42 ? _GEN_304 : plru1_9; // @[Cache.scala 131:22 137:27]
  wire  _GEN_433 = _T_42 ? _GEN_305 : plru1_10; // @[Cache.scala 131:22 137:27]
  wire  _GEN_434 = _T_42 ? _GEN_306 : plru1_11; // @[Cache.scala 131:22 137:27]
  wire  _GEN_435 = _T_42 ? _GEN_307 : plru1_12; // @[Cache.scala 131:22 137:27]
  wire  _GEN_436 = _T_42 ? _GEN_308 : plru1_13; // @[Cache.scala 131:22 137:27]
  wire  _GEN_437 = _T_42 ? _GEN_309 : plru1_14; // @[Cache.scala 131:22 137:27]
  wire  _GEN_438 = _T_42 ? _GEN_310 : plru1_15; // @[Cache.scala 131:22 137:27]
  wire  _GEN_439 = _T_42 ? _GEN_311 : plru1_16; // @[Cache.scala 131:22 137:27]
  wire  _GEN_440 = _T_42 ? _GEN_312 : plru1_17; // @[Cache.scala 131:22 137:27]
  wire  _GEN_441 = _T_42 ? _GEN_313 : plru1_18; // @[Cache.scala 131:22 137:27]
  wire  _GEN_442 = _T_42 ? _GEN_314 : plru1_19; // @[Cache.scala 131:22 137:27]
  wire  _GEN_443 = _T_42 ? _GEN_315 : plru1_20; // @[Cache.scala 131:22 137:27]
  wire  _GEN_444 = _T_42 ? _GEN_316 : plru1_21; // @[Cache.scala 131:22 137:27]
  wire  _GEN_445 = _T_42 ? _GEN_317 : plru1_22; // @[Cache.scala 131:22 137:27]
  wire  _GEN_446 = _T_42 ? _GEN_318 : plru1_23; // @[Cache.scala 131:22 137:27]
  wire  _GEN_447 = _T_42 ? _GEN_319 : plru1_24; // @[Cache.scala 131:22 137:27]
  wire  _GEN_448 = _T_42 ? _GEN_320 : plru1_25; // @[Cache.scala 131:22 137:27]
  wire  _GEN_449 = _T_42 ? _GEN_321 : plru1_26; // @[Cache.scala 131:22 137:27]
  wire  _GEN_450 = _T_42 ? _GEN_322 : plru1_27; // @[Cache.scala 131:22 137:27]
  wire  _GEN_451 = _T_42 ? _GEN_323 : plru1_28; // @[Cache.scala 131:22 137:27]
  wire  _GEN_452 = _T_42 ? _GEN_324 : plru1_29; // @[Cache.scala 131:22 137:27]
  wire  _GEN_453 = _T_42 ? _GEN_325 : plru1_30; // @[Cache.scala 131:22 137:27]
  wire  _GEN_454 = _T_42 ? _GEN_326 : plru1_31; // @[Cache.scala 131:22 137:27]
  wire  _GEN_455 = _T_42 ? _GEN_327 : plru1_32; // @[Cache.scala 131:22 137:27]
  wire  _GEN_456 = _T_42 ? _GEN_328 : plru1_33; // @[Cache.scala 131:22 137:27]
  wire  _GEN_457 = _T_42 ? _GEN_329 : plru1_34; // @[Cache.scala 131:22 137:27]
  wire  _GEN_458 = _T_42 ? _GEN_330 : plru1_35; // @[Cache.scala 131:22 137:27]
  wire  _GEN_459 = _T_42 ? _GEN_331 : plru1_36; // @[Cache.scala 131:22 137:27]
  wire  _GEN_460 = _T_42 ? _GEN_332 : plru1_37; // @[Cache.scala 131:22 137:27]
  wire  _GEN_461 = _T_42 ? _GEN_333 : plru1_38; // @[Cache.scala 131:22 137:27]
  wire  _GEN_462 = _T_42 ? _GEN_334 : plru1_39; // @[Cache.scala 131:22 137:27]
  wire  _GEN_463 = _T_42 ? _GEN_335 : plru1_40; // @[Cache.scala 131:22 137:27]
  wire  _GEN_464 = _T_42 ? _GEN_336 : plru1_41; // @[Cache.scala 131:22 137:27]
  wire  _GEN_465 = _T_42 ? _GEN_337 : plru1_42; // @[Cache.scala 131:22 137:27]
  wire  _GEN_466 = _T_42 ? _GEN_338 : plru1_43; // @[Cache.scala 131:22 137:27]
  wire  _GEN_467 = _T_42 ? _GEN_339 : plru1_44; // @[Cache.scala 131:22 137:27]
  wire  _GEN_468 = _T_42 ? _GEN_340 : plru1_45; // @[Cache.scala 131:22 137:27]
  wire  _GEN_469 = _T_42 ? _GEN_341 : plru1_46; // @[Cache.scala 131:22 137:27]
  wire  _GEN_470 = _T_42 ? _GEN_342 : plru1_47; // @[Cache.scala 131:22 137:27]
  wire  _GEN_471 = _T_42 ? _GEN_343 : plru1_48; // @[Cache.scala 131:22 137:27]
  wire  _GEN_472 = _T_42 ? _GEN_344 : plru1_49; // @[Cache.scala 131:22 137:27]
  wire  _GEN_473 = _T_42 ? _GEN_345 : plru1_50; // @[Cache.scala 131:22 137:27]
  wire  _GEN_474 = _T_42 ? _GEN_346 : plru1_51; // @[Cache.scala 131:22 137:27]
  wire  _GEN_475 = _T_42 ? _GEN_347 : plru1_52; // @[Cache.scala 131:22 137:27]
  wire  _GEN_476 = _T_42 ? _GEN_348 : plru1_53; // @[Cache.scala 131:22 137:27]
  wire  _GEN_477 = _T_42 ? _GEN_349 : plru1_54; // @[Cache.scala 131:22 137:27]
  wire  _GEN_478 = _T_42 ? _GEN_350 : plru1_55; // @[Cache.scala 131:22 137:27]
  wire  _GEN_479 = _T_42 ? _GEN_351 : plru1_56; // @[Cache.scala 131:22 137:27]
  wire  _GEN_480 = _T_42 ? _GEN_352 : plru1_57; // @[Cache.scala 131:22 137:27]
  wire  _GEN_481 = _T_42 ? _GEN_353 : plru1_58; // @[Cache.scala 131:22 137:27]
  wire  _GEN_482 = _T_42 ? _GEN_354 : plru1_59; // @[Cache.scala 131:22 137:27]
  wire  _GEN_483 = _T_42 ? _GEN_355 : plru1_60; // @[Cache.scala 131:22 137:27]
  wire  _GEN_484 = _T_42 ? _GEN_356 : plru1_61; // @[Cache.scala 131:22 137:27]
  wire  _GEN_485 = _T_42 ? _GEN_357 : plru1_62; // @[Cache.scala 131:22 137:27]
  wire  _GEN_486 = _T_42 ? _GEN_358 : plru1_63; // @[Cache.scala 131:22 137:27]
  wire  _GEN_487 = _T_42 ? plru2_0 : _GEN_359; // @[Cache.scala 133:22 137:27]
  wire  _GEN_488 = _T_42 ? plru2_1 : _GEN_360; // @[Cache.scala 133:22 137:27]
  wire  _GEN_489 = _T_42 ? plru2_2 : _GEN_361; // @[Cache.scala 133:22 137:27]
  wire  _GEN_490 = _T_42 ? plru2_3 : _GEN_362; // @[Cache.scala 133:22 137:27]
  wire  _GEN_491 = _T_42 ? plru2_4 : _GEN_363; // @[Cache.scala 133:22 137:27]
  wire  _GEN_492 = _T_42 ? plru2_5 : _GEN_364; // @[Cache.scala 133:22 137:27]
  wire  _GEN_493 = _T_42 ? plru2_6 : _GEN_365; // @[Cache.scala 133:22 137:27]
  wire  _GEN_494 = _T_42 ? plru2_7 : _GEN_366; // @[Cache.scala 133:22 137:27]
  wire  _GEN_495 = _T_42 ? plru2_8 : _GEN_367; // @[Cache.scala 133:22 137:27]
  wire  _GEN_496 = _T_42 ? plru2_9 : _GEN_368; // @[Cache.scala 133:22 137:27]
  wire  _GEN_497 = _T_42 ? plru2_10 : _GEN_369; // @[Cache.scala 133:22 137:27]
  wire  _GEN_498 = _T_42 ? plru2_11 : _GEN_370; // @[Cache.scala 133:22 137:27]
  wire  _GEN_499 = _T_42 ? plru2_12 : _GEN_371; // @[Cache.scala 133:22 137:27]
  wire  _GEN_500 = _T_42 ? plru2_13 : _GEN_372; // @[Cache.scala 133:22 137:27]
  wire  _GEN_501 = _T_42 ? plru2_14 : _GEN_373; // @[Cache.scala 133:22 137:27]
  wire  _GEN_502 = _T_42 ? plru2_15 : _GEN_374; // @[Cache.scala 133:22 137:27]
  wire  _GEN_503 = _T_42 ? plru2_16 : _GEN_375; // @[Cache.scala 133:22 137:27]
  wire  _GEN_504 = _T_42 ? plru2_17 : _GEN_376; // @[Cache.scala 133:22 137:27]
  wire  _GEN_505 = _T_42 ? plru2_18 : _GEN_377; // @[Cache.scala 133:22 137:27]
  wire  _GEN_506 = _T_42 ? plru2_19 : _GEN_378; // @[Cache.scala 133:22 137:27]
  wire  _GEN_507 = _T_42 ? plru2_20 : _GEN_379; // @[Cache.scala 133:22 137:27]
  wire  _GEN_508 = _T_42 ? plru2_21 : _GEN_380; // @[Cache.scala 133:22 137:27]
  wire  _GEN_509 = _T_42 ? plru2_22 : _GEN_381; // @[Cache.scala 133:22 137:27]
  wire  _GEN_510 = _T_42 ? plru2_23 : _GEN_382; // @[Cache.scala 133:22 137:27]
  wire  _GEN_511 = _T_42 ? plru2_24 : _GEN_383; // @[Cache.scala 133:22 137:27]
  wire  _GEN_512 = _T_42 ? plru2_25 : _GEN_384; // @[Cache.scala 133:22 137:27]
  wire  _GEN_513 = _T_42 ? plru2_26 : _GEN_385; // @[Cache.scala 133:22 137:27]
  wire  _GEN_514 = _T_42 ? plru2_27 : _GEN_386; // @[Cache.scala 133:22 137:27]
  wire  _GEN_515 = _T_42 ? plru2_28 : _GEN_387; // @[Cache.scala 133:22 137:27]
  wire  _GEN_516 = _T_42 ? plru2_29 : _GEN_388; // @[Cache.scala 133:22 137:27]
  wire  _GEN_517 = _T_42 ? plru2_30 : _GEN_389; // @[Cache.scala 133:22 137:27]
  wire  _GEN_518 = _T_42 ? plru2_31 : _GEN_390; // @[Cache.scala 133:22 137:27]
  wire  _GEN_519 = _T_42 ? plru2_32 : _GEN_391; // @[Cache.scala 133:22 137:27]
  wire  _GEN_520 = _T_42 ? plru2_33 : _GEN_392; // @[Cache.scala 133:22 137:27]
  wire  _GEN_521 = _T_42 ? plru2_34 : _GEN_393; // @[Cache.scala 133:22 137:27]
  wire  _GEN_522 = _T_42 ? plru2_35 : _GEN_394; // @[Cache.scala 133:22 137:27]
  wire  _GEN_523 = _T_42 ? plru2_36 : _GEN_395; // @[Cache.scala 133:22 137:27]
  wire  _GEN_524 = _T_42 ? plru2_37 : _GEN_396; // @[Cache.scala 133:22 137:27]
  wire  _GEN_525 = _T_42 ? plru2_38 : _GEN_397; // @[Cache.scala 133:22 137:27]
  wire  _GEN_526 = _T_42 ? plru2_39 : _GEN_398; // @[Cache.scala 133:22 137:27]
  wire  _GEN_527 = _T_42 ? plru2_40 : _GEN_399; // @[Cache.scala 133:22 137:27]
  wire  _GEN_528 = _T_42 ? plru2_41 : _GEN_400; // @[Cache.scala 133:22 137:27]
  wire  _GEN_529 = _T_42 ? plru2_42 : _GEN_401; // @[Cache.scala 133:22 137:27]
  wire  _GEN_530 = _T_42 ? plru2_43 : _GEN_402; // @[Cache.scala 133:22 137:27]
  wire  _GEN_531 = _T_42 ? plru2_44 : _GEN_403; // @[Cache.scala 133:22 137:27]
  wire  _GEN_532 = _T_42 ? plru2_45 : _GEN_404; // @[Cache.scala 133:22 137:27]
  wire  _GEN_533 = _T_42 ? plru2_46 : _GEN_405; // @[Cache.scala 133:22 137:27]
  wire  _GEN_534 = _T_42 ? plru2_47 : _GEN_406; // @[Cache.scala 133:22 137:27]
  wire  _GEN_535 = _T_42 ? plru2_48 : _GEN_407; // @[Cache.scala 133:22 137:27]
  wire  _GEN_536 = _T_42 ? plru2_49 : _GEN_408; // @[Cache.scala 133:22 137:27]
  wire  _GEN_537 = _T_42 ? plru2_50 : _GEN_409; // @[Cache.scala 133:22 137:27]
  wire  _GEN_538 = _T_42 ? plru2_51 : _GEN_410; // @[Cache.scala 133:22 137:27]
  wire  _GEN_539 = _T_42 ? plru2_52 : _GEN_411; // @[Cache.scala 133:22 137:27]
  wire  _GEN_540 = _T_42 ? plru2_53 : _GEN_412; // @[Cache.scala 133:22 137:27]
  wire  _GEN_541 = _T_42 ? plru2_54 : _GEN_413; // @[Cache.scala 133:22 137:27]
  wire  _GEN_542 = _T_42 ? plru2_55 : _GEN_414; // @[Cache.scala 133:22 137:27]
  wire  _GEN_543 = _T_42 ? plru2_56 : _GEN_415; // @[Cache.scala 133:22 137:27]
  wire  _GEN_544 = _T_42 ? plru2_57 : _GEN_416; // @[Cache.scala 133:22 137:27]
  wire  _GEN_545 = _T_42 ? plru2_58 : _GEN_417; // @[Cache.scala 133:22 137:27]
  wire  _GEN_546 = _T_42 ? plru2_59 : _GEN_418; // @[Cache.scala 133:22 137:27]
  wire  _GEN_547 = _T_42 ? plru2_60 : _GEN_419; // @[Cache.scala 133:22 137:27]
  wire  _GEN_548 = _T_42 ? plru2_61 : _GEN_420; // @[Cache.scala 133:22 137:27]
  wire  _GEN_549 = _T_42 ? plru2_62 : _GEN_421; // @[Cache.scala 133:22 137:27]
  wire  _GEN_550 = _T_42 ? plru2_63 : _GEN_422; // @[Cache.scala 133:22 137:27]
  wire [3:0] _GEN_759 = ~s2_hit ? 4'h1 : state; // @[Cache.scala 344:31 345:17 213:22]
  wire [3:0] _GEN_985 = REG_11 ? _GEN_759 : state; // @[Cache.scala 213:22 325:37]
  wire  _T_320 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_986 = _T_320 ? 4'h2 : state; // @[Cache.scala 350:29 351:15 213:22]
  wire  _T_322 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_987 = ~io_out_resp_bits_rlast ? io_out_resp_bits_rdata : wdata1; // @[Cache.scala 356:37 357:18 270:23]
  wire [63:0] _GEN_988 = ~io_out_resp_bits_rlast ? wdata2 : io_out_resp_bits_rdata; // @[Cache.scala 271:23 356:37 359:18]
  wire [3:0] _GEN_989 = ~io_out_resp_bits_rlast ? state : 4'h3; // @[Cache.scala 213:22 356:37 360:17]
  wire [63:0] _GEN_990 = _T_322 ? _GEN_987 : wdata1; // @[Cache.scala 270:23 355:30]
  wire [63:0] _GEN_991 = _T_322 ? _GEN_988 : wdata2; // @[Cache.scala 271:23 355:30]
  wire [3:0] _GEN_992 = _T_322 ? _GEN_989 : state; // @[Cache.scala 213:22 355:30]
  wire  _T_325 = replace_way == 2'h0; // @[Cache.scala 366:27]
  wire [127:0] _T_356 = {wdata2,wdata1}; // @[Cat.scala 30:58]
  wire  _GEN_994 = replace_way == 2'h0 | pipeline_ready; // @[Cache.scala 366:36 367:25]
  wire [5:0] _GEN_996 = replace_way == 2'h0 ? s2_idx : _GEN_3; // @[Cache.scala 366:36 369:27]
  wire [127:0] _GEN_997 = replace_way == 2'h0 ? _T_356 : 128'h0; // @[Cache.scala 110:16 366:36]
  wire [20:0] _GEN_998 = replace_way == 2'h0 ? s2_tag : 21'h0; // @[Cache.scala 114:16 366:36 380:28]
  wire  _T_389 = replace_way == 2'h1; // @[Cache.scala 366:27]
  wire  _GEN_1001 = replace_way == 2'h1 | pipeline_ready; // @[Cache.scala 366:36 367:25]
  wire [5:0] _GEN_1003 = replace_way == 2'h1 ? s2_idx : _GEN_3; // @[Cache.scala 366:36 369:27]
  wire [127:0] _GEN_1004 = replace_way == 2'h1 ? _T_356 : 128'h0; // @[Cache.scala 110:16 366:36]
  wire [20:0] _GEN_1005 = replace_way == 2'h1 ? s2_tag : 21'h0; // @[Cache.scala 114:16 366:36 380:28]
  wire  _T_453 = replace_way == 2'h2; // @[Cache.scala 366:27]
  wire  _GEN_1008 = replace_way == 2'h2 | pipeline_ready; // @[Cache.scala 366:36 367:25]
  wire [5:0] _GEN_1010 = replace_way == 2'h2 ? s2_idx : _GEN_3; // @[Cache.scala 366:36 369:27]
  wire [127:0] _GEN_1011 = replace_way == 2'h2 ? _T_356 : 128'h0; // @[Cache.scala 110:16 366:36]
  wire [20:0] _GEN_1012 = replace_way == 2'h2 ? s2_tag : 21'h0; // @[Cache.scala 114:16 366:36 380:28]
  wire  _T_517 = replace_way == 2'h3; // @[Cache.scala 366:27]
  wire  _GEN_1015 = replace_way == 2'h3 | pipeline_ready; // @[Cache.scala 366:36 367:25]
  wire [5:0] _GEN_1017 = replace_way == 2'h3 ? s2_idx : _GEN_3; // @[Cache.scala 366:36 369:27]
  wire [127:0] _GEN_1018 = replace_way == 2'h3 ? _T_356 : 128'h0; // @[Cache.scala 110:16 366:36]
  wire [20:0] _GEN_1019 = replace_way == 2'h3 ? s2_tag : 21'h0; // @[Cache.scala 114:16 366:36 380:28]
  wire  _T_582 = ~replace_way[1]; // @[Cache.scala 136:19]
  wire  _GEN_1021 = 6'h0 == s2_idx ? ~replace_way[1] : plru0_0; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1022 = 6'h1 == s2_idx ? ~replace_way[1] : plru0_1; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1023 = 6'h2 == s2_idx ? ~replace_way[1] : plru0_2; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1024 = 6'h3 == s2_idx ? ~replace_way[1] : plru0_3; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1025 = 6'h4 == s2_idx ? ~replace_way[1] : plru0_4; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1026 = 6'h5 == s2_idx ? ~replace_way[1] : plru0_5; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1027 = 6'h6 == s2_idx ? ~replace_way[1] : plru0_6; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1028 = 6'h7 == s2_idx ? ~replace_way[1] : plru0_7; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1029 = 6'h8 == s2_idx ? ~replace_way[1] : plru0_8; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1030 = 6'h9 == s2_idx ? ~replace_way[1] : plru0_9; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1031 = 6'ha == s2_idx ? ~replace_way[1] : plru0_10; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1032 = 6'hb == s2_idx ? ~replace_way[1] : plru0_11; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1033 = 6'hc == s2_idx ? ~replace_way[1] : plru0_12; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1034 = 6'hd == s2_idx ? ~replace_way[1] : plru0_13; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1035 = 6'he == s2_idx ? ~replace_way[1] : plru0_14; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1036 = 6'hf == s2_idx ? ~replace_way[1] : plru0_15; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1037 = 6'h10 == s2_idx ? ~replace_way[1] : plru0_16; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1038 = 6'h11 == s2_idx ? ~replace_way[1] : plru0_17; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1039 = 6'h12 == s2_idx ? ~replace_way[1] : plru0_18; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1040 = 6'h13 == s2_idx ? ~replace_way[1] : plru0_19; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1041 = 6'h14 == s2_idx ? ~replace_way[1] : plru0_20; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1042 = 6'h15 == s2_idx ? ~replace_way[1] : plru0_21; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1043 = 6'h16 == s2_idx ? ~replace_way[1] : plru0_22; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1044 = 6'h17 == s2_idx ? ~replace_way[1] : plru0_23; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1045 = 6'h18 == s2_idx ? ~replace_way[1] : plru0_24; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1046 = 6'h19 == s2_idx ? ~replace_way[1] : plru0_25; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1047 = 6'h1a == s2_idx ? ~replace_way[1] : plru0_26; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1048 = 6'h1b == s2_idx ? ~replace_way[1] : plru0_27; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1049 = 6'h1c == s2_idx ? ~replace_way[1] : plru0_28; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1050 = 6'h1d == s2_idx ? ~replace_way[1] : plru0_29; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1051 = 6'h1e == s2_idx ? ~replace_way[1] : plru0_30; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1052 = 6'h1f == s2_idx ? ~replace_way[1] : plru0_31; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1053 = 6'h20 == s2_idx ? ~replace_way[1] : plru0_32; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1054 = 6'h21 == s2_idx ? ~replace_way[1] : plru0_33; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1055 = 6'h22 == s2_idx ? ~replace_way[1] : plru0_34; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1056 = 6'h23 == s2_idx ? ~replace_way[1] : plru0_35; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1057 = 6'h24 == s2_idx ? ~replace_way[1] : plru0_36; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1058 = 6'h25 == s2_idx ? ~replace_way[1] : plru0_37; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1059 = 6'h26 == s2_idx ? ~replace_way[1] : plru0_38; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1060 = 6'h27 == s2_idx ? ~replace_way[1] : plru0_39; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1061 = 6'h28 == s2_idx ? ~replace_way[1] : plru0_40; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1062 = 6'h29 == s2_idx ? ~replace_way[1] : plru0_41; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1063 = 6'h2a == s2_idx ? ~replace_way[1] : plru0_42; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1064 = 6'h2b == s2_idx ? ~replace_way[1] : plru0_43; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1065 = 6'h2c == s2_idx ? ~replace_way[1] : plru0_44; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1066 = 6'h2d == s2_idx ? ~replace_way[1] : plru0_45; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1067 = 6'h2e == s2_idx ? ~replace_way[1] : plru0_46; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1068 = 6'h2f == s2_idx ? ~replace_way[1] : plru0_47; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1069 = 6'h30 == s2_idx ? ~replace_way[1] : plru0_48; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1070 = 6'h31 == s2_idx ? ~replace_way[1] : plru0_49; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1071 = 6'h32 == s2_idx ? ~replace_way[1] : plru0_50; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1072 = 6'h33 == s2_idx ? ~replace_way[1] : plru0_51; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1073 = 6'h34 == s2_idx ? ~replace_way[1] : plru0_52; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1074 = 6'h35 == s2_idx ? ~replace_way[1] : plru0_53; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1075 = 6'h36 == s2_idx ? ~replace_way[1] : plru0_54; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1076 = 6'h37 == s2_idx ? ~replace_way[1] : plru0_55; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1077 = 6'h38 == s2_idx ? ~replace_way[1] : plru0_56; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1078 = 6'h39 == s2_idx ? ~replace_way[1] : plru0_57; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1079 = 6'h3a == s2_idx ? ~replace_way[1] : plru0_58; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1080 = 6'h3b == s2_idx ? ~replace_way[1] : plru0_59; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1081 = 6'h3c == s2_idx ? ~replace_way[1] : plru0_60; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1082 = 6'h3d == s2_idx ? ~replace_way[1] : plru0_61; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1083 = 6'h3e == s2_idx ? ~replace_way[1] : plru0_62; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1084 = 6'h3f == s2_idx ? ~replace_way[1] : plru0_63; // @[Cache.scala 136:{16,16} 129:22]
  wire  _T_586 = ~replace_way[0]; // @[Cache.scala 138:21]
  wire  _GEN_1085 = 6'h0 == s2_idx ? ~replace_way[0] : plru1_0; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1086 = 6'h1 == s2_idx ? ~replace_way[0] : plru1_1; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1087 = 6'h2 == s2_idx ? ~replace_way[0] : plru1_2; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1088 = 6'h3 == s2_idx ? ~replace_way[0] : plru1_3; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1089 = 6'h4 == s2_idx ? ~replace_way[0] : plru1_4; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1090 = 6'h5 == s2_idx ? ~replace_way[0] : plru1_5; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1091 = 6'h6 == s2_idx ? ~replace_way[0] : plru1_6; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1092 = 6'h7 == s2_idx ? ~replace_way[0] : plru1_7; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1093 = 6'h8 == s2_idx ? ~replace_way[0] : plru1_8; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1094 = 6'h9 == s2_idx ? ~replace_way[0] : plru1_9; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1095 = 6'ha == s2_idx ? ~replace_way[0] : plru1_10; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1096 = 6'hb == s2_idx ? ~replace_way[0] : plru1_11; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1097 = 6'hc == s2_idx ? ~replace_way[0] : plru1_12; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1098 = 6'hd == s2_idx ? ~replace_way[0] : plru1_13; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1099 = 6'he == s2_idx ? ~replace_way[0] : plru1_14; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1100 = 6'hf == s2_idx ? ~replace_way[0] : plru1_15; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1101 = 6'h10 == s2_idx ? ~replace_way[0] : plru1_16; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1102 = 6'h11 == s2_idx ? ~replace_way[0] : plru1_17; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1103 = 6'h12 == s2_idx ? ~replace_way[0] : plru1_18; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1104 = 6'h13 == s2_idx ? ~replace_way[0] : plru1_19; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1105 = 6'h14 == s2_idx ? ~replace_way[0] : plru1_20; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1106 = 6'h15 == s2_idx ? ~replace_way[0] : plru1_21; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1107 = 6'h16 == s2_idx ? ~replace_way[0] : plru1_22; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1108 = 6'h17 == s2_idx ? ~replace_way[0] : plru1_23; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1109 = 6'h18 == s2_idx ? ~replace_way[0] : plru1_24; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1110 = 6'h19 == s2_idx ? ~replace_way[0] : plru1_25; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1111 = 6'h1a == s2_idx ? ~replace_way[0] : plru1_26; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1112 = 6'h1b == s2_idx ? ~replace_way[0] : plru1_27; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1113 = 6'h1c == s2_idx ? ~replace_way[0] : plru1_28; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1114 = 6'h1d == s2_idx ? ~replace_way[0] : plru1_29; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1115 = 6'h1e == s2_idx ? ~replace_way[0] : plru1_30; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1116 = 6'h1f == s2_idx ? ~replace_way[0] : plru1_31; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1117 = 6'h20 == s2_idx ? ~replace_way[0] : plru1_32; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1118 = 6'h21 == s2_idx ? ~replace_way[0] : plru1_33; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1119 = 6'h22 == s2_idx ? ~replace_way[0] : plru1_34; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1120 = 6'h23 == s2_idx ? ~replace_way[0] : plru1_35; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1121 = 6'h24 == s2_idx ? ~replace_way[0] : plru1_36; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1122 = 6'h25 == s2_idx ? ~replace_way[0] : plru1_37; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1123 = 6'h26 == s2_idx ? ~replace_way[0] : plru1_38; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1124 = 6'h27 == s2_idx ? ~replace_way[0] : plru1_39; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1125 = 6'h28 == s2_idx ? ~replace_way[0] : plru1_40; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1126 = 6'h29 == s2_idx ? ~replace_way[0] : plru1_41; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1127 = 6'h2a == s2_idx ? ~replace_way[0] : plru1_42; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1128 = 6'h2b == s2_idx ? ~replace_way[0] : plru1_43; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1129 = 6'h2c == s2_idx ? ~replace_way[0] : plru1_44; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1130 = 6'h2d == s2_idx ? ~replace_way[0] : plru1_45; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1131 = 6'h2e == s2_idx ? ~replace_way[0] : plru1_46; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1132 = 6'h2f == s2_idx ? ~replace_way[0] : plru1_47; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1133 = 6'h30 == s2_idx ? ~replace_way[0] : plru1_48; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1134 = 6'h31 == s2_idx ? ~replace_way[0] : plru1_49; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1135 = 6'h32 == s2_idx ? ~replace_way[0] : plru1_50; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1136 = 6'h33 == s2_idx ? ~replace_way[0] : plru1_51; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1137 = 6'h34 == s2_idx ? ~replace_way[0] : plru1_52; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1138 = 6'h35 == s2_idx ? ~replace_way[0] : plru1_53; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1139 = 6'h36 == s2_idx ? ~replace_way[0] : plru1_54; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1140 = 6'h37 == s2_idx ? ~replace_way[0] : plru1_55; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1141 = 6'h38 == s2_idx ? ~replace_way[0] : plru1_56; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1142 = 6'h39 == s2_idx ? ~replace_way[0] : plru1_57; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1143 = 6'h3a == s2_idx ? ~replace_way[0] : plru1_58; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1144 = 6'h3b == s2_idx ? ~replace_way[0] : plru1_59; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1145 = 6'h3c == s2_idx ? ~replace_way[0] : plru1_60; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1146 = 6'h3d == s2_idx ? ~replace_way[0] : plru1_61; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1147 = 6'h3e == s2_idx ? ~replace_way[0] : plru1_62; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1148 = 6'h3f == s2_idx ? ~replace_way[0] : plru1_63; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1149 = 6'h0 == s2_idx ? _T_586 : plru2_0; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1150 = 6'h1 == s2_idx ? _T_586 : plru2_1; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1151 = 6'h2 == s2_idx ? _T_586 : plru2_2; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1152 = 6'h3 == s2_idx ? _T_586 : plru2_3; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1153 = 6'h4 == s2_idx ? _T_586 : plru2_4; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1154 = 6'h5 == s2_idx ? _T_586 : plru2_5; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1155 = 6'h6 == s2_idx ? _T_586 : plru2_6; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1156 = 6'h7 == s2_idx ? _T_586 : plru2_7; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1157 = 6'h8 == s2_idx ? _T_586 : plru2_8; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1158 = 6'h9 == s2_idx ? _T_586 : plru2_9; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1159 = 6'ha == s2_idx ? _T_586 : plru2_10; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1160 = 6'hb == s2_idx ? _T_586 : plru2_11; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1161 = 6'hc == s2_idx ? _T_586 : plru2_12; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1162 = 6'hd == s2_idx ? _T_586 : plru2_13; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1163 = 6'he == s2_idx ? _T_586 : plru2_14; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1164 = 6'hf == s2_idx ? _T_586 : plru2_15; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1165 = 6'h10 == s2_idx ? _T_586 : plru2_16; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1166 = 6'h11 == s2_idx ? _T_586 : plru2_17; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1167 = 6'h12 == s2_idx ? _T_586 : plru2_18; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1168 = 6'h13 == s2_idx ? _T_586 : plru2_19; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1169 = 6'h14 == s2_idx ? _T_586 : plru2_20; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1170 = 6'h15 == s2_idx ? _T_586 : plru2_21; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1171 = 6'h16 == s2_idx ? _T_586 : plru2_22; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1172 = 6'h17 == s2_idx ? _T_586 : plru2_23; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1173 = 6'h18 == s2_idx ? _T_586 : plru2_24; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1174 = 6'h19 == s2_idx ? _T_586 : plru2_25; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1175 = 6'h1a == s2_idx ? _T_586 : plru2_26; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1176 = 6'h1b == s2_idx ? _T_586 : plru2_27; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1177 = 6'h1c == s2_idx ? _T_586 : plru2_28; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1178 = 6'h1d == s2_idx ? _T_586 : plru2_29; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1179 = 6'h1e == s2_idx ? _T_586 : plru2_30; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1180 = 6'h1f == s2_idx ? _T_586 : plru2_31; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1181 = 6'h20 == s2_idx ? _T_586 : plru2_32; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1182 = 6'h21 == s2_idx ? _T_586 : plru2_33; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1183 = 6'h22 == s2_idx ? _T_586 : plru2_34; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1184 = 6'h23 == s2_idx ? _T_586 : plru2_35; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1185 = 6'h24 == s2_idx ? _T_586 : plru2_36; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1186 = 6'h25 == s2_idx ? _T_586 : plru2_37; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1187 = 6'h26 == s2_idx ? _T_586 : plru2_38; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1188 = 6'h27 == s2_idx ? _T_586 : plru2_39; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1189 = 6'h28 == s2_idx ? _T_586 : plru2_40; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1190 = 6'h29 == s2_idx ? _T_586 : plru2_41; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1191 = 6'h2a == s2_idx ? _T_586 : plru2_42; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1192 = 6'h2b == s2_idx ? _T_586 : plru2_43; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1193 = 6'h2c == s2_idx ? _T_586 : plru2_44; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1194 = 6'h2d == s2_idx ? _T_586 : plru2_45; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1195 = 6'h2e == s2_idx ? _T_586 : plru2_46; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1196 = 6'h2f == s2_idx ? _T_586 : plru2_47; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1197 = 6'h30 == s2_idx ? _T_586 : plru2_48; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1198 = 6'h31 == s2_idx ? _T_586 : plru2_49; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1199 = 6'h32 == s2_idx ? _T_586 : plru2_50; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1200 = 6'h33 == s2_idx ? _T_586 : plru2_51; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1201 = 6'h34 == s2_idx ? _T_586 : plru2_52; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1202 = 6'h35 == s2_idx ? _T_586 : plru2_53; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1203 = 6'h36 == s2_idx ? _T_586 : plru2_54; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1204 = 6'h37 == s2_idx ? _T_586 : plru2_55; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1205 = 6'h38 == s2_idx ? _T_586 : plru2_56; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1206 = 6'h39 == s2_idx ? _T_586 : plru2_57; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1207 = 6'h3a == s2_idx ? _T_586 : plru2_58; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1208 = 6'h3b == s2_idx ? _T_586 : plru2_59; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1209 = 6'h3c == s2_idx ? _T_586 : plru2_60; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1210 = 6'h3d == s2_idx ? _T_586 : plru2_61; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1211 = 6'h3e == s2_idx ? _T_586 : plru2_62; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1212 = 6'h3f == s2_idx ? _T_586 : plru2_63; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1213 = _T_582 ? _GEN_1085 : plru1_0; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1214 = _T_582 ? _GEN_1086 : plru1_1; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1215 = _T_582 ? _GEN_1087 : plru1_2; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1216 = _T_582 ? _GEN_1088 : plru1_3; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1217 = _T_582 ? _GEN_1089 : plru1_4; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1218 = _T_582 ? _GEN_1090 : plru1_5; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1219 = _T_582 ? _GEN_1091 : plru1_6; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1220 = _T_582 ? _GEN_1092 : plru1_7; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1221 = _T_582 ? _GEN_1093 : plru1_8; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1222 = _T_582 ? _GEN_1094 : plru1_9; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1223 = _T_582 ? _GEN_1095 : plru1_10; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1224 = _T_582 ? _GEN_1096 : plru1_11; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1225 = _T_582 ? _GEN_1097 : plru1_12; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1226 = _T_582 ? _GEN_1098 : plru1_13; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1227 = _T_582 ? _GEN_1099 : plru1_14; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1228 = _T_582 ? _GEN_1100 : plru1_15; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1229 = _T_582 ? _GEN_1101 : plru1_16; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1230 = _T_582 ? _GEN_1102 : plru1_17; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1231 = _T_582 ? _GEN_1103 : plru1_18; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1232 = _T_582 ? _GEN_1104 : plru1_19; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1233 = _T_582 ? _GEN_1105 : plru1_20; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1234 = _T_582 ? _GEN_1106 : plru1_21; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1235 = _T_582 ? _GEN_1107 : plru1_22; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1236 = _T_582 ? _GEN_1108 : plru1_23; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1237 = _T_582 ? _GEN_1109 : plru1_24; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1238 = _T_582 ? _GEN_1110 : plru1_25; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1239 = _T_582 ? _GEN_1111 : plru1_26; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1240 = _T_582 ? _GEN_1112 : plru1_27; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1241 = _T_582 ? _GEN_1113 : plru1_28; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1242 = _T_582 ? _GEN_1114 : plru1_29; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1243 = _T_582 ? _GEN_1115 : plru1_30; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1244 = _T_582 ? _GEN_1116 : plru1_31; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1245 = _T_582 ? _GEN_1117 : plru1_32; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1246 = _T_582 ? _GEN_1118 : plru1_33; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1247 = _T_582 ? _GEN_1119 : plru1_34; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1248 = _T_582 ? _GEN_1120 : plru1_35; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1249 = _T_582 ? _GEN_1121 : plru1_36; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1250 = _T_582 ? _GEN_1122 : plru1_37; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1251 = _T_582 ? _GEN_1123 : plru1_38; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1252 = _T_582 ? _GEN_1124 : plru1_39; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1253 = _T_582 ? _GEN_1125 : plru1_40; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1254 = _T_582 ? _GEN_1126 : plru1_41; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1255 = _T_582 ? _GEN_1127 : plru1_42; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1256 = _T_582 ? _GEN_1128 : plru1_43; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1257 = _T_582 ? _GEN_1129 : plru1_44; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1258 = _T_582 ? _GEN_1130 : plru1_45; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1259 = _T_582 ? _GEN_1131 : plru1_46; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1260 = _T_582 ? _GEN_1132 : plru1_47; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1261 = _T_582 ? _GEN_1133 : plru1_48; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1262 = _T_582 ? _GEN_1134 : plru1_49; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1263 = _T_582 ? _GEN_1135 : plru1_50; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1264 = _T_582 ? _GEN_1136 : plru1_51; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1265 = _T_582 ? _GEN_1137 : plru1_52; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1266 = _T_582 ? _GEN_1138 : plru1_53; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1267 = _T_582 ? _GEN_1139 : plru1_54; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1268 = _T_582 ? _GEN_1140 : plru1_55; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1269 = _T_582 ? _GEN_1141 : plru1_56; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1270 = _T_582 ? _GEN_1142 : plru1_57; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1271 = _T_582 ? _GEN_1143 : plru1_58; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1272 = _T_582 ? _GEN_1144 : plru1_59; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1273 = _T_582 ? _GEN_1145 : plru1_60; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1274 = _T_582 ? _GEN_1146 : plru1_61; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1275 = _T_582 ? _GEN_1147 : plru1_62; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1276 = _T_582 ? _GEN_1148 : plru1_63; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1277 = _T_582 ? plru2_0 : _GEN_1149; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1278 = _T_582 ? plru2_1 : _GEN_1150; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1279 = _T_582 ? plru2_2 : _GEN_1151; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1280 = _T_582 ? plru2_3 : _GEN_1152; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1281 = _T_582 ? plru2_4 : _GEN_1153; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1282 = _T_582 ? plru2_5 : _GEN_1154; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1283 = _T_582 ? plru2_6 : _GEN_1155; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1284 = _T_582 ? plru2_7 : _GEN_1156; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1285 = _T_582 ? plru2_8 : _GEN_1157; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1286 = _T_582 ? plru2_9 : _GEN_1158; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1287 = _T_582 ? plru2_10 : _GEN_1159; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1288 = _T_582 ? plru2_11 : _GEN_1160; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1289 = _T_582 ? plru2_12 : _GEN_1161; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1290 = _T_582 ? plru2_13 : _GEN_1162; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1291 = _T_582 ? plru2_14 : _GEN_1163; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1292 = _T_582 ? plru2_15 : _GEN_1164; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1293 = _T_582 ? plru2_16 : _GEN_1165; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1294 = _T_582 ? plru2_17 : _GEN_1166; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1295 = _T_582 ? plru2_18 : _GEN_1167; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1296 = _T_582 ? plru2_19 : _GEN_1168; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1297 = _T_582 ? plru2_20 : _GEN_1169; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1298 = _T_582 ? plru2_21 : _GEN_1170; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1299 = _T_582 ? plru2_22 : _GEN_1171; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1300 = _T_582 ? plru2_23 : _GEN_1172; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1301 = _T_582 ? plru2_24 : _GEN_1173; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1302 = _T_582 ? plru2_25 : _GEN_1174; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1303 = _T_582 ? plru2_26 : _GEN_1175; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1304 = _T_582 ? plru2_27 : _GEN_1176; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1305 = _T_582 ? plru2_28 : _GEN_1177; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1306 = _T_582 ? plru2_29 : _GEN_1178; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1307 = _T_582 ? plru2_30 : _GEN_1179; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1308 = _T_582 ? plru2_31 : _GEN_1180; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1309 = _T_582 ? plru2_32 : _GEN_1181; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1310 = _T_582 ? plru2_33 : _GEN_1182; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1311 = _T_582 ? plru2_34 : _GEN_1183; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1312 = _T_582 ? plru2_35 : _GEN_1184; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1313 = _T_582 ? plru2_36 : _GEN_1185; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1314 = _T_582 ? plru2_37 : _GEN_1186; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1315 = _T_582 ? plru2_38 : _GEN_1187; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1316 = _T_582 ? plru2_39 : _GEN_1188; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1317 = _T_582 ? plru2_40 : _GEN_1189; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1318 = _T_582 ? plru2_41 : _GEN_1190; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1319 = _T_582 ? plru2_42 : _GEN_1191; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1320 = _T_582 ? plru2_43 : _GEN_1192; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1321 = _T_582 ? plru2_44 : _GEN_1193; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1322 = _T_582 ? plru2_45 : _GEN_1194; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1323 = _T_582 ? plru2_46 : _GEN_1195; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1324 = _T_582 ? plru2_47 : _GEN_1196; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1325 = _T_582 ? plru2_48 : _GEN_1197; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1326 = _T_582 ? plru2_49 : _GEN_1198; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1327 = _T_582 ? plru2_50 : _GEN_1199; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1328 = _T_582 ? plru2_51 : _GEN_1200; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1329 = _T_582 ? plru2_52 : _GEN_1201; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1330 = _T_582 ? plru2_53 : _GEN_1202; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1331 = _T_582 ? plru2_54 : _GEN_1203; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1332 = _T_582 ? plru2_55 : _GEN_1204; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1333 = _T_582 ? plru2_56 : _GEN_1205; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1334 = _T_582 ? plru2_57 : _GEN_1206; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1335 = _T_582 ? plru2_58 : _GEN_1207; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1336 = _T_582 ? plru2_59 : _GEN_1208; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1337 = _T_582 ? plru2_60 : _GEN_1209; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1338 = _T_582 ? plru2_61 : _GEN_1210; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1339 = _T_582 ? plru2_62 : _GEN_1211; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1340 = _T_582 ? plru2_63 : _GEN_1212; // @[Cache.scala 133:22 137:27]
  wire [3:0] _GEN_1341 = s2_reg_dirty ? 4'h4 : 4'h7; // @[Cache.scala 385:27 386:15 389:15]
  wire  _GEN_1342 = s2_reg_dirty ? plru0_0 : _GEN_1021; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1343 = s2_reg_dirty ? plru0_1 : _GEN_1022; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1344 = s2_reg_dirty ? plru0_2 : _GEN_1023; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1345 = s2_reg_dirty ? plru0_3 : _GEN_1024; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1346 = s2_reg_dirty ? plru0_4 : _GEN_1025; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1347 = s2_reg_dirty ? plru0_5 : _GEN_1026; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1348 = s2_reg_dirty ? plru0_6 : _GEN_1027; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1349 = s2_reg_dirty ? plru0_7 : _GEN_1028; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1350 = s2_reg_dirty ? plru0_8 : _GEN_1029; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1351 = s2_reg_dirty ? plru0_9 : _GEN_1030; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1352 = s2_reg_dirty ? plru0_10 : _GEN_1031; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1353 = s2_reg_dirty ? plru0_11 : _GEN_1032; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1354 = s2_reg_dirty ? plru0_12 : _GEN_1033; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1355 = s2_reg_dirty ? plru0_13 : _GEN_1034; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1356 = s2_reg_dirty ? plru0_14 : _GEN_1035; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1357 = s2_reg_dirty ? plru0_15 : _GEN_1036; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1358 = s2_reg_dirty ? plru0_16 : _GEN_1037; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1359 = s2_reg_dirty ? plru0_17 : _GEN_1038; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1360 = s2_reg_dirty ? plru0_18 : _GEN_1039; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1361 = s2_reg_dirty ? plru0_19 : _GEN_1040; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1362 = s2_reg_dirty ? plru0_20 : _GEN_1041; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1363 = s2_reg_dirty ? plru0_21 : _GEN_1042; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1364 = s2_reg_dirty ? plru0_22 : _GEN_1043; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1365 = s2_reg_dirty ? plru0_23 : _GEN_1044; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1366 = s2_reg_dirty ? plru0_24 : _GEN_1045; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1367 = s2_reg_dirty ? plru0_25 : _GEN_1046; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1368 = s2_reg_dirty ? plru0_26 : _GEN_1047; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1369 = s2_reg_dirty ? plru0_27 : _GEN_1048; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1370 = s2_reg_dirty ? plru0_28 : _GEN_1049; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1371 = s2_reg_dirty ? plru0_29 : _GEN_1050; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1372 = s2_reg_dirty ? plru0_30 : _GEN_1051; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1373 = s2_reg_dirty ? plru0_31 : _GEN_1052; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1374 = s2_reg_dirty ? plru0_32 : _GEN_1053; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1375 = s2_reg_dirty ? plru0_33 : _GEN_1054; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1376 = s2_reg_dirty ? plru0_34 : _GEN_1055; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1377 = s2_reg_dirty ? plru0_35 : _GEN_1056; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1378 = s2_reg_dirty ? plru0_36 : _GEN_1057; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1379 = s2_reg_dirty ? plru0_37 : _GEN_1058; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1380 = s2_reg_dirty ? plru0_38 : _GEN_1059; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1381 = s2_reg_dirty ? plru0_39 : _GEN_1060; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1382 = s2_reg_dirty ? plru0_40 : _GEN_1061; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1383 = s2_reg_dirty ? plru0_41 : _GEN_1062; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1384 = s2_reg_dirty ? plru0_42 : _GEN_1063; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1385 = s2_reg_dirty ? plru0_43 : _GEN_1064; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1386 = s2_reg_dirty ? plru0_44 : _GEN_1065; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1387 = s2_reg_dirty ? plru0_45 : _GEN_1066; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1388 = s2_reg_dirty ? plru0_46 : _GEN_1067; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1389 = s2_reg_dirty ? plru0_47 : _GEN_1068; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1390 = s2_reg_dirty ? plru0_48 : _GEN_1069; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1391 = s2_reg_dirty ? plru0_49 : _GEN_1070; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1392 = s2_reg_dirty ? plru0_50 : _GEN_1071; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1393 = s2_reg_dirty ? plru0_51 : _GEN_1072; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1394 = s2_reg_dirty ? plru0_52 : _GEN_1073; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1395 = s2_reg_dirty ? plru0_53 : _GEN_1074; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1396 = s2_reg_dirty ? plru0_54 : _GEN_1075; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1397 = s2_reg_dirty ? plru0_55 : _GEN_1076; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1398 = s2_reg_dirty ? plru0_56 : _GEN_1077; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1399 = s2_reg_dirty ? plru0_57 : _GEN_1078; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1400 = s2_reg_dirty ? plru0_58 : _GEN_1079; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1401 = s2_reg_dirty ? plru0_59 : _GEN_1080; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1402 = s2_reg_dirty ? plru0_60 : _GEN_1081; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1403 = s2_reg_dirty ? plru0_61 : _GEN_1082; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1404 = s2_reg_dirty ? plru0_62 : _GEN_1083; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1405 = s2_reg_dirty ? plru0_63 : _GEN_1084; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1406 = s2_reg_dirty ? plru1_0 : _GEN_1213; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1407 = s2_reg_dirty ? plru1_1 : _GEN_1214; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1408 = s2_reg_dirty ? plru1_2 : _GEN_1215; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1409 = s2_reg_dirty ? plru1_3 : _GEN_1216; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1410 = s2_reg_dirty ? plru1_4 : _GEN_1217; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1411 = s2_reg_dirty ? plru1_5 : _GEN_1218; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1412 = s2_reg_dirty ? plru1_6 : _GEN_1219; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1413 = s2_reg_dirty ? plru1_7 : _GEN_1220; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1414 = s2_reg_dirty ? plru1_8 : _GEN_1221; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1415 = s2_reg_dirty ? plru1_9 : _GEN_1222; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1416 = s2_reg_dirty ? plru1_10 : _GEN_1223; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1417 = s2_reg_dirty ? plru1_11 : _GEN_1224; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1418 = s2_reg_dirty ? plru1_12 : _GEN_1225; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1419 = s2_reg_dirty ? plru1_13 : _GEN_1226; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1420 = s2_reg_dirty ? plru1_14 : _GEN_1227; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1421 = s2_reg_dirty ? plru1_15 : _GEN_1228; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1422 = s2_reg_dirty ? plru1_16 : _GEN_1229; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1423 = s2_reg_dirty ? plru1_17 : _GEN_1230; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1424 = s2_reg_dirty ? plru1_18 : _GEN_1231; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1425 = s2_reg_dirty ? plru1_19 : _GEN_1232; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1426 = s2_reg_dirty ? plru1_20 : _GEN_1233; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1427 = s2_reg_dirty ? plru1_21 : _GEN_1234; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1428 = s2_reg_dirty ? plru1_22 : _GEN_1235; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1429 = s2_reg_dirty ? plru1_23 : _GEN_1236; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1430 = s2_reg_dirty ? plru1_24 : _GEN_1237; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1431 = s2_reg_dirty ? plru1_25 : _GEN_1238; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1432 = s2_reg_dirty ? plru1_26 : _GEN_1239; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1433 = s2_reg_dirty ? plru1_27 : _GEN_1240; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1434 = s2_reg_dirty ? plru1_28 : _GEN_1241; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1435 = s2_reg_dirty ? plru1_29 : _GEN_1242; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1436 = s2_reg_dirty ? plru1_30 : _GEN_1243; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1437 = s2_reg_dirty ? plru1_31 : _GEN_1244; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1438 = s2_reg_dirty ? plru1_32 : _GEN_1245; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1439 = s2_reg_dirty ? plru1_33 : _GEN_1246; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1440 = s2_reg_dirty ? plru1_34 : _GEN_1247; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1441 = s2_reg_dirty ? plru1_35 : _GEN_1248; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1442 = s2_reg_dirty ? plru1_36 : _GEN_1249; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1443 = s2_reg_dirty ? plru1_37 : _GEN_1250; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1444 = s2_reg_dirty ? plru1_38 : _GEN_1251; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1445 = s2_reg_dirty ? plru1_39 : _GEN_1252; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1446 = s2_reg_dirty ? plru1_40 : _GEN_1253; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1447 = s2_reg_dirty ? plru1_41 : _GEN_1254; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1448 = s2_reg_dirty ? plru1_42 : _GEN_1255; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1449 = s2_reg_dirty ? plru1_43 : _GEN_1256; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1450 = s2_reg_dirty ? plru1_44 : _GEN_1257; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1451 = s2_reg_dirty ? plru1_45 : _GEN_1258; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1452 = s2_reg_dirty ? plru1_46 : _GEN_1259; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1453 = s2_reg_dirty ? plru1_47 : _GEN_1260; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1454 = s2_reg_dirty ? plru1_48 : _GEN_1261; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1455 = s2_reg_dirty ? plru1_49 : _GEN_1262; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1456 = s2_reg_dirty ? plru1_50 : _GEN_1263; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1457 = s2_reg_dirty ? plru1_51 : _GEN_1264; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1458 = s2_reg_dirty ? plru1_52 : _GEN_1265; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1459 = s2_reg_dirty ? plru1_53 : _GEN_1266; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1460 = s2_reg_dirty ? plru1_54 : _GEN_1267; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1461 = s2_reg_dirty ? plru1_55 : _GEN_1268; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1462 = s2_reg_dirty ? plru1_56 : _GEN_1269; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1463 = s2_reg_dirty ? plru1_57 : _GEN_1270; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1464 = s2_reg_dirty ? plru1_58 : _GEN_1271; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1465 = s2_reg_dirty ? plru1_59 : _GEN_1272; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1466 = s2_reg_dirty ? plru1_60 : _GEN_1273; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1467 = s2_reg_dirty ? plru1_61 : _GEN_1274; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1468 = s2_reg_dirty ? plru1_62 : _GEN_1275; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1469 = s2_reg_dirty ? plru1_63 : _GEN_1276; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1470 = s2_reg_dirty ? plru2_0 : _GEN_1277; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1471 = s2_reg_dirty ? plru2_1 : _GEN_1278; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1472 = s2_reg_dirty ? plru2_2 : _GEN_1279; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1473 = s2_reg_dirty ? plru2_3 : _GEN_1280; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1474 = s2_reg_dirty ? plru2_4 : _GEN_1281; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1475 = s2_reg_dirty ? plru2_5 : _GEN_1282; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1476 = s2_reg_dirty ? plru2_6 : _GEN_1283; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1477 = s2_reg_dirty ? plru2_7 : _GEN_1284; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1478 = s2_reg_dirty ? plru2_8 : _GEN_1285; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1479 = s2_reg_dirty ? plru2_9 : _GEN_1286; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1480 = s2_reg_dirty ? plru2_10 : _GEN_1287; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1481 = s2_reg_dirty ? plru2_11 : _GEN_1288; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1482 = s2_reg_dirty ? plru2_12 : _GEN_1289; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1483 = s2_reg_dirty ? plru2_13 : _GEN_1290; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1484 = s2_reg_dirty ? plru2_14 : _GEN_1291; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1485 = s2_reg_dirty ? plru2_15 : _GEN_1292; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1486 = s2_reg_dirty ? plru2_16 : _GEN_1293; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1487 = s2_reg_dirty ? plru2_17 : _GEN_1294; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1488 = s2_reg_dirty ? plru2_18 : _GEN_1295; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1489 = s2_reg_dirty ? plru2_19 : _GEN_1296; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1490 = s2_reg_dirty ? plru2_20 : _GEN_1297; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1491 = s2_reg_dirty ? plru2_21 : _GEN_1298; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1492 = s2_reg_dirty ? plru2_22 : _GEN_1299; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1493 = s2_reg_dirty ? plru2_23 : _GEN_1300; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1494 = s2_reg_dirty ? plru2_24 : _GEN_1301; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1495 = s2_reg_dirty ? plru2_25 : _GEN_1302; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1496 = s2_reg_dirty ? plru2_26 : _GEN_1303; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1497 = s2_reg_dirty ? plru2_27 : _GEN_1304; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1498 = s2_reg_dirty ? plru2_28 : _GEN_1305; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1499 = s2_reg_dirty ? plru2_29 : _GEN_1306; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1500 = s2_reg_dirty ? plru2_30 : _GEN_1307; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1501 = s2_reg_dirty ? plru2_31 : _GEN_1308; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1502 = s2_reg_dirty ? plru2_32 : _GEN_1309; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1503 = s2_reg_dirty ? plru2_33 : _GEN_1310; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1504 = s2_reg_dirty ? plru2_34 : _GEN_1311; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1505 = s2_reg_dirty ? plru2_35 : _GEN_1312; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1506 = s2_reg_dirty ? plru2_36 : _GEN_1313; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1507 = s2_reg_dirty ? plru2_37 : _GEN_1314; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1508 = s2_reg_dirty ? plru2_38 : _GEN_1315; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1509 = s2_reg_dirty ? plru2_39 : _GEN_1316; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1510 = s2_reg_dirty ? plru2_40 : _GEN_1317; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1511 = s2_reg_dirty ? plru2_41 : _GEN_1318; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1512 = s2_reg_dirty ? plru2_42 : _GEN_1319; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1513 = s2_reg_dirty ? plru2_43 : _GEN_1320; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1514 = s2_reg_dirty ? plru2_44 : _GEN_1321; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1515 = s2_reg_dirty ? plru2_45 : _GEN_1322; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1516 = s2_reg_dirty ? plru2_46 : _GEN_1323; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1517 = s2_reg_dirty ? plru2_47 : _GEN_1324; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1518 = s2_reg_dirty ? plru2_48 : _GEN_1325; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1519 = s2_reg_dirty ? plru2_49 : _GEN_1326; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1520 = s2_reg_dirty ? plru2_50 : _GEN_1327; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1521 = s2_reg_dirty ? plru2_51 : _GEN_1328; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1522 = s2_reg_dirty ? plru2_52 : _GEN_1329; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1523 = s2_reg_dirty ? plru2_53 : _GEN_1330; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1524 = s2_reg_dirty ? plru2_54 : _GEN_1331; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1525 = s2_reg_dirty ? plru2_55 : _GEN_1332; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1526 = s2_reg_dirty ? plru2_56 : _GEN_1333; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1527 = s2_reg_dirty ? plru2_57 : _GEN_1334; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1528 = s2_reg_dirty ? plru2_58 : _GEN_1335; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1529 = s2_reg_dirty ? plru2_59 : _GEN_1336; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1530 = s2_reg_dirty ? plru2_60 : _GEN_1337; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1531 = s2_reg_dirty ? plru2_61 : _GEN_1338; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1532 = s2_reg_dirty ? plru2_62 : _GEN_1339; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1533 = s2_reg_dirty ? plru2_63 : _GEN_1340; // @[Cache.scala 133:22 385:27]
  wire [3:0] _GEN_1534 = _T_320 ? 4'h5 : state; // @[Cache.scala 393:29 394:15 213:22]
  wire [3:0] _GEN_1535 = _T_320 ? 4'h6 : state; // @[Cache.scala 398:29 399:15 213:22]
  wire  _GEN_1856 = _T_322 ? _GEN_1021 : plru0_0; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1857 = _T_322 ? _GEN_1022 : plru0_1; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1858 = _T_322 ? _GEN_1023 : plru0_2; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1859 = _T_322 ? _GEN_1024 : plru0_3; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1860 = _T_322 ? _GEN_1025 : plru0_4; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1861 = _T_322 ? _GEN_1026 : plru0_5; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1862 = _T_322 ? _GEN_1027 : plru0_6; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1863 = _T_322 ? _GEN_1028 : plru0_7; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1864 = _T_322 ? _GEN_1029 : plru0_8; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1865 = _T_322 ? _GEN_1030 : plru0_9; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1866 = _T_322 ? _GEN_1031 : plru0_10; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1867 = _T_322 ? _GEN_1032 : plru0_11; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1868 = _T_322 ? _GEN_1033 : plru0_12; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1869 = _T_322 ? _GEN_1034 : plru0_13; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1870 = _T_322 ? _GEN_1035 : plru0_14; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1871 = _T_322 ? _GEN_1036 : plru0_15; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1872 = _T_322 ? _GEN_1037 : plru0_16; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1873 = _T_322 ? _GEN_1038 : plru0_17; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1874 = _T_322 ? _GEN_1039 : plru0_18; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1875 = _T_322 ? _GEN_1040 : plru0_19; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1876 = _T_322 ? _GEN_1041 : plru0_20; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1877 = _T_322 ? _GEN_1042 : plru0_21; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1878 = _T_322 ? _GEN_1043 : plru0_22; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1879 = _T_322 ? _GEN_1044 : plru0_23; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1880 = _T_322 ? _GEN_1045 : plru0_24; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1881 = _T_322 ? _GEN_1046 : plru0_25; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1882 = _T_322 ? _GEN_1047 : plru0_26; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1883 = _T_322 ? _GEN_1048 : plru0_27; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1884 = _T_322 ? _GEN_1049 : plru0_28; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1885 = _T_322 ? _GEN_1050 : plru0_29; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1886 = _T_322 ? _GEN_1051 : plru0_30; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1887 = _T_322 ? _GEN_1052 : plru0_31; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1888 = _T_322 ? _GEN_1053 : plru0_32; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1889 = _T_322 ? _GEN_1054 : plru0_33; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1890 = _T_322 ? _GEN_1055 : plru0_34; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1891 = _T_322 ? _GEN_1056 : plru0_35; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1892 = _T_322 ? _GEN_1057 : plru0_36; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1893 = _T_322 ? _GEN_1058 : plru0_37; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1894 = _T_322 ? _GEN_1059 : plru0_38; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1895 = _T_322 ? _GEN_1060 : plru0_39; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1896 = _T_322 ? _GEN_1061 : plru0_40; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1897 = _T_322 ? _GEN_1062 : plru0_41; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1898 = _T_322 ? _GEN_1063 : plru0_42; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1899 = _T_322 ? _GEN_1064 : plru0_43; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1900 = _T_322 ? _GEN_1065 : plru0_44; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1901 = _T_322 ? _GEN_1066 : plru0_45; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1902 = _T_322 ? _GEN_1067 : plru0_46; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1903 = _T_322 ? _GEN_1068 : plru0_47; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1904 = _T_322 ? _GEN_1069 : plru0_48; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1905 = _T_322 ? _GEN_1070 : plru0_49; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1906 = _T_322 ? _GEN_1071 : plru0_50; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1907 = _T_322 ? _GEN_1072 : plru0_51; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1908 = _T_322 ? _GEN_1073 : plru0_52; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1909 = _T_322 ? _GEN_1074 : plru0_53; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1910 = _T_322 ? _GEN_1075 : plru0_54; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1911 = _T_322 ? _GEN_1076 : plru0_55; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1912 = _T_322 ? _GEN_1077 : plru0_56; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1913 = _T_322 ? _GEN_1078 : plru0_57; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1914 = _T_322 ? _GEN_1079 : plru0_58; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1915 = _T_322 ? _GEN_1080 : plru0_59; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1916 = _T_322 ? _GEN_1081 : plru0_60; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1917 = _T_322 ? _GEN_1082 : plru0_61; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1918 = _T_322 ? _GEN_1083 : plru0_62; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1919 = _T_322 ? _GEN_1084 : plru0_63; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1920 = _T_322 ? _GEN_1213 : plru1_0; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1921 = _T_322 ? _GEN_1214 : plru1_1; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1922 = _T_322 ? _GEN_1215 : plru1_2; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1923 = _T_322 ? _GEN_1216 : plru1_3; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1924 = _T_322 ? _GEN_1217 : plru1_4; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1925 = _T_322 ? _GEN_1218 : plru1_5; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1926 = _T_322 ? _GEN_1219 : plru1_6; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1927 = _T_322 ? _GEN_1220 : plru1_7; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1928 = _T_322 ? _GEN_1221 : plru1_8; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1929 = _T_322 ? _GEN_1222 : plru1_9; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1930 = _T_322 ? _GEN_1223 : plru1_10; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1931 = _T_322 ? _GEN_1224 : plru1_11; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1932 = _T_322 ? _GEN_1225 : plru1_12; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1933 = _T_322 ? _GEN_1226 : plru1_13; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1934 = _T_322 ? _GEN_1227 : plru1_14; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1935 = _T_322 ? _GEN_1228 : plru1_15; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1936 = _T_322 ? _GEN_1229 : plru1_16; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1937 = _T_322 ? _GEN_1230 : plru1_17; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1938 = _T_322 ? _GEN_1231 : plru1_18; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1939 = _T_322 ? _GEN_1232 : plru1_19; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1940 = _T_322 ? _GEN_1233 : plru1_20; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1941 = _T_322 ? _GEN_1234 : plru1_21; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1942 = _T_322 ? _GEN_1235 : plru1_22; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1943 = _T_322 ? _GEN_1236 : plru1_23; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1944 = _T_322 ? _GEN_1237 : plru1_24; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1945 = _T_322 ? _GEN_1238 : plru1_25; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1946 = _T_322 ? _GEN_1239 : plru1_26; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1947 = _T_322 ? _GEN_1240 : plru1_27; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1948 = _T_322 ? _GEN_1241 : plru1_28; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1949 = _T_322 ? _GEN_1242 : plru1_29; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1950 = _T_322 ? _GEN_1243 : plru1_30; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1951 = _T_322 ? _GEN_1244 : plru1_31; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1952 = _T_322 ? _GEN_1245 : plru1_32; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1953 = _T_322 ? _GEN_1246 : plru1_33; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1954 = _T_322 ? _GEN_1247 : plru1_34; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1955 = _T_322 ? _GEN_1248 : plru1_35; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1956 = _T_322 ? _GEN_1249 : plru1_36; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1957 = _T_322 ? _GEN_1250 : plru1_37; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1958 = _T_322 ? _GEN_1251 : plru1_38; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1959 = _T_322 ? _GEN_1252 : plru1_39; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1960 = _T_322 ? _GEN_1253 : plru1_40; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1961 = _T_322 ? _GEN_1254 : plru1_41; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1962 = _T_322 ? _GEN_1255 : plru1_42; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1963 = _T_322 ? _GEN_1256 : plru1_43; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1964 = _T_322 ? _GEN_1257 : plru1_44; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1965 = _T_322 ? _GEN_1258 : plru1_45; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1966 = _T_322 ? _GEN_1259 : plru1_46; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1967 = _T_322 ? _GEN_1260 : plru1_47; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1968 = _T_322 ? _GEN_1261 : plru1_48; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1969 = _T_322 ? _GEN_1262 : plru1_49; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1970 = _T_322 ? _GEN_1263 : plru1_50; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1971 = _T_322 ? _GEN_1264 : plru1_51; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1972 = _T_322 ? _GEN_1265 : plru1_52; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1973 = _T_322 ? _GEN_1266 : plru1_53; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1974 = _T_322 ? _GEN_1267 : plru1_54; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1975 = _T_322 ? _GEN_1268 : plru1_55; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1976 = _T_322 ? _GEN_1269 : plru1_56; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1977 = _T_322 ? _GEN_1270 : plru1_57; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1978 = _T_322 ? _GEN_1271 : plru1_58; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1979 = _T_322 ? _GEN_1272 : plru1_59; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1980 = _T_322 ? _GEN_1273 : plru1_60; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1981 = _T_322 ? _GEN_1274 : plru1_61; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1982 = _T_322 ? _GEN_1275 : plru1_62; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1983 = _T_322 ? _GEN_1276 : plru1_63; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1984 = _T_322 ? _GEN_1277 : plru2_0; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1985 = _T_322 ? _GEN_1278 : plru2_1; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1986 = _T_322 ? _GEN_1279 : plru2_2; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1987 = _T_322 ? _GEN_1280 : plru2_3; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1988 = _T_322 ? _GEN_1281 : plru2_4; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1989 = _T_322 ? _GEN_1282 : plru2_5; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1990 = _T_322 ? _GEN_1283 : plru2_6; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1991 = _T_322 ? _GEN_1284 : plru2_7; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1992 = _T_322 ? _GEN_1285 : plru2_8; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1993 = _T_322 ? _GEN_1286 : plru2_9; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1994 = _T_322 ? _GEN_1287 : plru2_10; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1995 = _T_322 ? _GEN_1288 : plru2_11; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1996 = _T_322 ? _GEN_1289 : plru2_12; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1997 = _T_322 ? _GEN_1290 : plru2_13; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1998 = _T_322 ? _GEN_1291 : plru2_14; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1999 = _T_322 ? _GEN_1292 : plru2_15; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2000 = _T_322 ? _GEN_1293 : plru2_16; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2001 = _T_322 ? _GEN_1294 : plru2_17; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2002 = _T_322 ? _GEN_1295 : plru2_18; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2003 = _T_322 ? _GEN_1296 : plru2_19; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2004 = _T_322 ? _GEN_1297 : plru2_20; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2005 = _T_322 ? _GEN_1298 : plru2_21; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2006 = _T_322 ? _GEN_1299 : plru2_22; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2007 = _T_322 ? _GEN_1300 : plru2_23; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2008 = _T_322 ? _GEN_1301 : plru2_24; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2009 = _T_322 ? _GEN_1302 : plru2_25; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2010 = _T_322 ? _GEN_1303 : plru2_26; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2011 = _T_322 ? _GEN_1304 : plru2_27; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2012 = _T_322 ? _GEN_1305 : plru2_28; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2013 = _T_322 ? _GEN_1306 : plru2_29; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2014 = _T_322 ? _GEN_1307 : plru2_30; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2015 = _T_322 ? _GEN_1308 : plru2_31; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2016 = _T_322 ? _GEN_1309 : plru2_32; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2017 = _T_322 ? _GEN_1310 : plru2_33; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2018 = _T_322 ? _GEN_1311 : plru2_34; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2019 = _T_322 ? _GEN_1312 : plru2_35; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2020 = _T_322 ? _GEN_1313 : plru2_36; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2021 = _T_322 ? _GEN_1314 : plru2_37; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2022 = _T_322 ? _GEN_1315 : plru2_38; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2023 = _T_322 ? _GEN_1316 : plru2_39; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2024 = _T_322 ? _GEN_1317 : plru2_40; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2025 = _T_322 ? _GEN_1318 : plru2_41; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2026 = _T_322 ? _GEN_1319 : plru2_42; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2027 = _T_322 ? _GEN_1320 : plru2_43; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2028 = _T_322 ? _GEN_1321 : plru2_44; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2029 = _T_322 ? _GEN_1322 : plru2_45; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2030 = _T_322 ? _GEN_1323 : plru2_46; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2031 = _T_322 ? _GEN_1324 : plru2_47; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2032 = _T_322 ? _GEN_1325 : plru2_48; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2033 = _T_322 ? _GEN_1326 : plru2_49; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2034 = _T_322 ? _GEN_1327 : plru2_50; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2035 = _T_322 ? _GEN_1328 : plru2_51; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2036 = _T_322 ? _GEN_1329 : plru2_52; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2037 = _T_322 ? _GEN_1330 : plru2_53; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2038 = _T_322 ? _GEN_1331 : plru2_54; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2039 = _T_322 ? _GEN_1332 : plru2_55; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2040 = _T_322 ? _GEN_1333 : plru2_56; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2041 = _T_322 ? _GEN_1334 : plru2_57; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2042 = _T_322 ? _GEN_1335 : plru2_58; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2043 = _T_322 ? _GEN_1336 : plru2_59; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2044 = _T_322 ? _GEN_1337 : plru2_60; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2045 = _T_322 ? _GEN_1338 : plru2_61; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2046 = _T_322 ? _GEN_1339 : plru2_62; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2047 = _T_322 ? _GEN_1340 : plru2_63; // @[Cache.scala 133:22 404:30]
  wire [3:0] _GEN_2048 = _T_322 ? 4'h7 : state; // @[Cache.scala 404:30 406:15 213:22]
  reg [63:0] REG_12; // @[Cache.scala 410:36]
  wire  _T_606 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_2049 = _T_606 ? 4'h8 : state; // @[Cache.scala 411:29 412:15 213:22]
  wire [63:0] _GEN_2050 = 4'h7 == state ? REG_12 : 64'h0; // @[Cache.scala 318:18 289:22 410:26]
  wire [3:0] _GEN_2051 = 4'h7 == state ? _GEN_2049 : state; // @[Cache.scala 318:18 213:22]
  wire  _GEN_2053 = 4'h6 == state ? _GEN_1856 : plru0_0; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2054 = 4'h6 == state ? _GEN_1857 : plru0_1; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2055 = 4'h6 == state ? _GEN_1858 : plru0_2; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2056 = 4'h6 == state ? _GEN_1859 : plru0_3; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2057 = 4'h6 == state ? _GEN_1860 : plru0_4; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2058 = 4'h6 == state ? _GEN_1861 : plru0_5; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2059 = 4'h6 == state ? _GEN_1862 : plru0_6; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2060 = 4'h6 == state ? _GEN_1863 : plru0_7; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2061 = 4'h6 == state ? _GEN_1864 : plru0_8; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2062 = 4'h6 == state ? _GEN_1865 : plru0_9; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2063 = 4'h6 == state ? _GEN_1866 : plru0_10; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2064 = 4'h6 == state ? _GEN_1867 : plru0_11; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2065 = 4'h6 == state ? _GEN_1868 : plru0_12; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2066 = 4'h6 == state ? _GEN_1869 : plru0_13; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2067 = 4'h6 == state ? _GEN_1870 : plru0_14; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2068 = 4'h6 == state ? _GEN_1871 : plru0_15; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2069 = 4'h6 == state ? _GEN_1872 : plru0_16; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2070 = 4'h6 == state ? _GEN_1873 : plru0_17; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2071 = 4'h6 == state ? _GEN_1874 : plru0_18; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2072 = 4'h6 == state ? _GEN_1875 : plru0_19; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2073 = 4'h6 == state ? _GEN_1876 : plru0_20; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2074 = 4'h6 == state ? _GEN_1877 : plru0_21; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2075 = 4'h6 == state ? _GEN_1878 : plru0_22; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2076 = 4'h6 == state ? _GEN_1879 : plru0_23; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2077 = 4'h6 == state ? _GEN_1880 : plru0_24; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2078 = 4'h6 == state ? _GEN_1881 : plru0_25; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2079 = 4'h6 == state ? _GEN_1882 : plru0_26; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2080 = 4'h6 == state ? _GEN_1883 : plru0_27; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2081 = 4'h6 == state ? _GEN_1884 : plru0_28; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2082 = 4'h6 == state ? _GEN_1885 : plru0_29; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2083 = 4'h6 == state ? _GEN_1886 : plru0_30; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2084 = 4'h6 == state ? _GEN_1887 : plru0_31; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2085 = 4'h6 == state ? _GEN_1888 : plru0_32; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2086 = 4'h6 == state ? _GEN_1889 : plru0_33; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2087 = 4'h6 == state ? _GEN_1890 : plru0_34; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2088 = 4'h6 == state ? _GEN_1891 : plru0_35; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2089 = 4'h6 == state ? _GEN_1892 : plru0_36; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2090 = 4'h6 == state ? _GEN_1893 : plru0_37; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2091 = 4'h6 == state ? _GEN_1894 : plru0_38; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2092 = 4'h6 == state ? _GEN_1895 : plru0_39; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2093 = 4'h6 == state ? _GEN_1896 : plru0_40; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2094 = 4'h6 == state ? _GEN_1897 : plru0_41; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2095 = 4'h6 == state ? _GEN_1898 : plru0_42; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2096 = 4'h6 == state ? _GEN_1899 : plru0_43; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2097 = 4'h6 == state ? _GEN_1900 : plru0_44; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2098 = 4'h6 == state ? _GEN_1901 : plru0_45; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2099 = 4'h6 == state ? _GEN_1902 : plru0_46; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2100 = 4'h6 == state ? _GEN_1903 : plru0_47; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2101 = 4'h6 == state ? _GEN_1904 : plru0_48; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2102 = 4'h6 == state ? _GEN_1905 : plru0_49; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2103 = 4'h6 == state ? _GEN_1906 : plru0_50; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2104 = 4'h6 == state ? _GEN_1907 : plru0_51; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2105 = 4'h6 == state ? _GEN_1908 : plru0_52; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2106 = 4'h6 == state ? _GEN_1909 : plru0_53; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2107 = 4'h6 == state ? _GEN_1910 : plru0_54; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2108 = 4'h6 == state ? _GEN_1911 : plru0_55; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2109 = 4'h6 == state ? _GEN_1912 : plru0_56; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2110 = 4'h6 == state ? _GEN_1913 : plru0_57; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2111 = 4'h6 == state ? _GEN_1914 : plru0_58; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2112 = 4'h6 == state ? _GEN_1915 : plru0_59; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2113 = 4'h6 == state ? _GEN_1916 : plru0_60; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2114 = 4'h6 == state ? _GEN_1917 : plru0_61; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2115 = 4'h6 == state ? _GEN_1918 : plru0_62; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2116 = 4'h6 == state ? _GEN_1919 : plru0_63; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2117 = 4'h6 == state ? _GEN_1920 : plru1_0; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2118 = 4'h6 == state ? _GEN_1921 : plru1_1; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2119 = 4'h6 == state ? _GEN_1922 : plru1_2; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2120 = 4'h6 == state ? _GEN_1923 : plru1_3; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2121 = 4'h6 == state ? _GEN_1924 : plru1_4; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2122 = 4'h6 == state ? _GEN_1925 : plru1_5; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2123 = 4'h6 == state ? _GEN_1926 : plru1_6; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2124 = 4'h6 == state ? _GEN_1927 : plru1_7; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2125 = 4'h6 == state ? _GEN_1928 : plru1_8; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2126 = 4'h6 == state ? _GEN_1929 : plru1_9; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2127 = 4'h6 == state ? _GEN_1930 : plru1_10; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2128 = 4'h6 == state ? _GEN_1931 : plru1_11; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2129 = 4'h6 == state ? _GEN_1932 : plru1_12; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2130 = 4'h6 == state ? _GEN_1933 : plru1_13; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2131 = 4'h6 == state ? _GEN_1934 : plru1_14; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2132 = 4'h6 == state ? _GEN_1935 : plru1_15; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2133 = 4'h6 == state ? _GEN_1936 : plru1_16; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2134 = 4'h6 == state ? _GEN_1937 : plru1_17; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2135 = 4'h6 == state ? _GEN_1938 : plru1_18; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2136 = 4'h6 == state ? _GEN_1939 : plru1_19; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2137 = 4'h6 == state ? _GEN_1940 : plru1_20; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2138 = 4'h6 == state ? _GEN_1941 : plru1_21; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2139 = 4'h6 == state ? _GEN_1942 : plru1_22; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2140 = 4'h6 == state ? _GEN_1943 : plru1_23; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2141 = 4'h6 == state ? _GEN_1944 : plru1_24; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2142 = 4'h6 == state ? _GEN_1945 : plru1_25; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2143 = 4'h6 == state ? _GEN_1946 : plru1_26; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2144 = 4'h6 == state ? _GEN_1947 : plru1_27; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2145 = 4'h6 == state ? _GEN_1948 : plru1_28; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2146 = 4'h6 == state ? _GEN_1949 : plru1_29; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2147 = 4'h6 == state ? _GEN_1950 : plru1_30; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2148 = 4'h6 == state ? _GEN_1951 : plru1_31; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2149 = 4'h6 == state ? _GEN_1952 : plru1_32; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2150 = 4'h6 == state ? _GEN_1953 : plru1_33; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2151 = 4'h6 == state ? _GEN_1954 : plru1_34; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2152 = 4'h6 == state ? _GEN_1955 : plru1_35; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2153 = 4'h6 == state ? _GEN_1956 : plru1_36; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2154 = 4'h6 == state ? _GEN_1957 : plru1_37; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2155 = 4'h6 == state ? _GEN_1958 : plru1_38; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2156 = 4'h6 == state ? _GEN_1959 : plru1_39; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2157 = 4'h6 == state ? _GEN_1960 : plru1_40; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2158 = 4'h6 == state ? _GEN_1961 : plru1_41; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2159 = 4'h6 == state ? _GEN_1962 : plru1_42; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2160 = 4'h6 == state ? _GEN_1963 : plru1_43; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2161 = 4'h6 == state ? _GEN_1964 : plru1_44; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2162 = 4'h6 == state ? _GEN_1965 : plru1_45; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2163 = 4'h6 == state ? _GEN_1966 : plru1_46; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2164 = 4'h6 == state ? _GEN_1967 : plru1_47; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2165 = 4'h6 == state ? _GEN_1968 : plru1_48; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2166 = 4'h6 == state ? _GEN_1969 : plru1_49; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2167 = 4'h6 == state ? _GEN_1970 : plru1_50; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2168 = 4'h6 == state ? _GEN_1971 : plru1_51; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2169 = 4'h6 == state ? _GEN_1972 : plru1_52; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2170 = 4'h6 == state ? _GEN_1973 : plru1_53; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2171 = 4'h6 == state ? _GEN_1974 : plru1_54; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2172 = 4'h6 == state ? _GEN_1975 : plru1_55; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2173 = 4'h6 == state ? _GEN_1976 : plru1_56; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2174 = 4'h6 == state ? _GEN_1977 : plru1_57; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2175 = 4'h6 == state ? _GEN_1978 : plru1_58; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2176 = 4'h6 == state ? _GEN_1979 : plru1_59; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2177 = 4'h6 == state ? _GEN_1980 : plru1_60; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2178 = 4'h6 == state ? _GEN_1981 : plru1_61; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2179 = 4'h6 == state ? _GEN_1982 : plru1_62; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2180 = 4'h6 == state ? _GEN_1983 : plru1_63; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2181 = 4'h6 == state ? _GEN_1984 : plru2_0; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2182 = 4'h6 == state ? _GEN_1985 : plru2_1; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2183 = 4'h6 == state ? _GEN_1986 : plru2_2; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2184 = 4'h6 == state ? _GEN_1987 : plru2_3; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2185 = 4'h6 == state ? _GEN_1988 : plru2_4; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2186 = 4'h6 == state ? _GEN_1989 : plru2_5; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2187 = 4'h6 == state ? _GEN_1990 : plru2_6; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2188 = 4'h6 == state ? _GEN_1991 : plru2_7; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2189 = 4'h6 == state ? _GEN_1992 : plru2_8; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2190 = 4'h6 == state ? _GEN_1993 : plru2_9; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2191 = 4'h6 == state ? _GEN_1994 : plru2_10; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2192 = 4'h6 == state ? _GEN_1995 : plru2_11; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2193 = 4'h6 == state ? _GEN_1996 : plru2_12; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2194 = 4'h6 == state ? _GEN_1997 : plru2_13; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2195 = 4'h6 == state ? _GEN_1998 : plru2_14; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2196 = 4'h6 == state ? _GEN_1999 : plru2_15; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2197 = 4'h6 == state ? _GEN_2000 : plru2_16; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2198 = 4'h6 == state ? _GEN_2001 : plru2_17; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2199 = 4'h6 == state ? _GEN_2002 : plru2_18; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2200 = 4'h6 == state ? _GEN_2003 : plru2_19; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2201 = 4'h6 == state ? _GEN_2004 : plru2_20; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2202 = 4'h6 == state ? _GEN_2005 : plru2_21; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2203 = 4'h6 == state ? _GEN_2006 : plru2_22; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2204 = 4'h6 == state ? _GEN_2007 : plru2_23; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2205 = 4'h6 == state ? _GEN_2008 : plru2_24; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2206 = 4'h6 == state ? _GEN_2009 : plru2_25; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2207 = 4'h6 == state ? _GEN_2010 : plru2_26; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2208 = 4'h6 == state ? _GEN_2011 : plru2_27; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2209 = 4'h6 == state ? _GEN_2012 : plru2_28; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2210 = 4'h6 == state ? _GEN_2013 : plru2_29; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2211 = 4'h6 == state ? _GEN_2014 : plru2_30; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2212 = 4'h6 == state ? _GEN_2015 : plru2_31; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2213 = 4'h6 == state ? _GEN_2016 : plru2_32; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2214 = 4'h6 == state ? _GEN_2017 : plru2_33; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2215 = 4'h6 == state ? _GEN_2018 : plru2_34; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2216 = 4'h6 == state ? _GEN_2019 : plru2_35; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2217 = 4'h6 == state ? _GEN_2020 : plru2_36; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2218 = 4'h6 == state ? _GEN_2021 : plru2_37; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2219 = 4'h6 == state ? _GEN_2022 : plru2_38; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2220 = 4'h6 == state ? _GEN_2023 : plru2_39; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2221 = 4'h6 == state ? _GEN_2024 : plru2_40; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2222 = 4'h6 == state ? _GEN_2025 : plru2_41; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2223 = 4'h6 == state ? _GEN_2026 : plru2_42; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2224 = 4'h6 == state ? _GEN_2027 : plru2_43; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2225 = 4'h6 == state ? _GEN_2028 : plru2_44; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2226 = 4'h6 == state ? _GEN_2029 : plru2_45; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2227 = 4'h6 == state ? _GEN_2030 : plru2_46; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2228 = 4'h6 == state ? _GEN_2031 : plru2_47; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2229 = 4'h6 == state ? _GEN_2032 : plru2_48; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2230 = 4'h6 == state ? _GEN_2033 : plru2_49; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2231 = 4'h6 == state ? _GEN_2034 : plru2_50; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2232 = 4'h6 == state ? _GEN_2035 : plru2_51; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2233 = 4'h6 == state ? _GEN_2036 : plru2_52; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2234 = 4'h6 == state ? _GEN_2037 : plru2_53; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2235 = 4'h6 == state ? _GEN_2038 : plru2_54; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2236 = 4'h6 == state ? _GEN_2039 : plru2_55; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2237 = 4'h6 == state ? _GEN_2040 : plru2_56; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2238 = 4'h6 == state ? _GEN_2041 : plru2_57; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2239 = 4'h6 == state ? _GEN_2042 : plru2_58; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2240 = 4'h6 == state ? _GEN_2043 : plru2_59; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2241 = 4'h6 == state ? _GEN_2044 : plru2_60; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2242 = 4'h6 == state ? _GEN_2045 : plru2_61; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2243 = 4'h6 == state ? _GEN_2046 : plru2_62; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2244 = 4'h6 == state ? _GEN_2047 : plru2_63; // @[Cache.scala 318:18 133:22]
  wire [3:0] _GEN_2245 = 4'h6 == state ? _GEN_2048 : _GEN_2051; // @[Cache.scala 318:18]
  wire [63:0] _GEN_2246 = 4'h6 == state ? 64'h0 : _GEN_2050; // @[Cache.scala 318:18 289:22]
  wire [3:0] _GEN_2247 = 4'h5 == state ? _GEN_1535 : _GEN_2245; // @[Cache.scala 318:18]
  wire  _GEN_2249 = 4'h5 == state ? plru0_0 : _GEN_2053; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2250 = 4'h5 == state ? plru0_1 : _GEN_2054; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2251 = 4'h5 == state ? plru0_2 : _GEN_2055; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2252 = 4'h5 == state ? plru0_3 : _GEN_2056; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2253 = 4'h5 == state ? plru0_4 : _GEN_2057; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2254 = 4'h5 == state ? plru0_5 : _GEN_2058; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2255 = 4'h5 == state ? plru0_6 : _GEN_2059; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2256 = 4'h5 == state ? plru0_7 : _GEN_2060; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2257 = 4'h5 == state ? plru0_8 : _GEN_2061; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2258 = 4'h5 == state ? plru0_9 : _GEN_2062; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2259 = 4'h5 == state ? plru0_10 : _GEN_2063; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2260 = 4'h5 == state ? plru0_11 : _GEN_2064; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2261 = 4'h5 == state ? plru0_12 : _GEN_2065; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2262 = 4'h5 == state ? plru0_13 : _GEN_2066; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2263 = 4'h5 == state ? plru0_14 : _GEN_2067; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2264 = 4'h5 == state ? plru0_15 : _GEN_2068; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2265 = 4'h5 == state ? plru0_16 : _GEN_2069; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2266 = 4'h5 == state ? plru0_17 : _GEN_2070; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2267 = 4'h5 == state ? plru0_18 : _GEN_2071; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2268 = 4'h5 == state ? plru0_19 : _GEN_2072; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2269 = 4'h5 == state ? plru0_20 : _GEN_2073; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2270 = 4'h5 == state ? plru0_21 : _GEN_2074; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2271 = 4'h5 == state ? plru0_22 : _GEN_2075; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2272 = 4'h5 == state ? plru0_23 : _GEN_2076; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2273 = 4'h5 == state ? plru0_24 : _GEN_2077; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2274 = 4'h5 == state ? plru0_25 : _GEN_2078; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2275 = 4'h5 == state ? plru0_26 : _GEN_2079; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2276 = 4'h5 == state ? plru0_27 : _GEN_2080; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2277 = 4'h5 == state ? plru0_28 : _GEN_2081; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2278 = 4'h5 == state ? plru0_29 : _GEN_2082; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2279 = 4'h5 == state ? plru0_30 : _GEN_2083; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2280 = 4'h5 == state ? plru0_31 : _GEN_2084; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2281 = 4'h5 == state ? plru0_32 : _GEN_2085; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2282 = 4'h5 == state ? plru0_33 : _GEN_2086; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2283 = 4'h5 == state ? plru0_34 : _GEN_2087; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2284 = 4'h5 == state ? plru0_35 : _GEN_2088; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2285 = 4'h5 == state ? plru0_36 : _GEN_2089; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2286 = 4'h5 == state ? plru0_37 : _GEN_2090; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2287 = 4'h5 == state ? plru0_38 : _GEN_2091; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2288 = 4'h5 == state ? plru0_39 : _GEN_2092; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2289 = 4'h5 == state ? plru0_40 : _GEN_2093; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2290 = 4'h5 == state ? plru0_41 : _GEN_2094; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2291 = 4'h5 == state ? plru0_42 : _GEN_2095; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2292 = 4'h5 == state ? plru0_43 : _GEN_2096; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2293 = 4'h5 == state ? plru0_44 : _GEN_2097; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2294 = 4'h5 == state ? plru0_45 : _GEN_2098; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2295 = 4'h5 == state ? plru0_46 : _GEN_2099; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2296 = 4'h5 == state ? plru0_47 : _GEN_2100; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2297 = 4'h5 == state ? plru0_48 : _GEN_2101; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2298 = 4'h5 == state ? plru0_49 : _GEN_2102; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2299 = 4'h5 == state ? plru0_50 : _GEN_2103; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2300 = 4'h5 == state ? plru0_51 : _GEN_2104; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2301 = 4'h5 == state ? plru0_52 : _GEN_2105; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2302 = 4'h5 == state ? plru0_53 : _GEN_2106; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2303 = 4'h5 == state ? plru0_54 : _GEN_2107; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2304 = 4'h5 == state ? plru0_55 : _GEN_2108; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2305 = 4'h5 == state ? plru0_56 : _GEN_2109; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2306 = 4'h5 == state ? plru0_57 : _GEN_2110; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2307 = 4'h5 == state ? plru0_58 : _GEN_2111; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2308 = 4'h5 == state ? plru0_59 : _GEN_2112; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2309 = 4'h5 == state ? plru0_60 : _GEN_2113; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2310 = 4'h5 == state ? plru0_61 : _GEN_2114; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2311 = 4'h5 == state ? plru0_62 : _GEN_2115; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2312 = 4'h5 == state ? plru0_63 : _GEN_2116; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2313 = 4'h5 == state ? plru1_0 : _GEN_2117; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2314 = 4'h5 == state ? plru1_1 : _GEN_2118; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2315 = 4'h5 == state ? plru1_2 : _GEN_2119; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2316 = 4'h5 == state ? plru1_3 : _GEN_2120; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2317 = 4'h5 == state ? plru1_4 : _GEN_2121; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2318 = 4'h5 == state ? plru1_5 : _GEN_2122; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2319 = 4'h5 == state ? plru1_6 : _GEN_2123; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2320 = 4'h5 == state ? plru1_7 : _GEN_2124; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2321 = 4'h5 == state ? plru1_8 : _GEN_2125; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2322 = 4'h5 == state ? plru1_9 : _GEN_2126; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2323 = 4'h5 == state ? plru1_10 : _GEN_2127; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2324 = 4'h5 == state ? plru1_11 : _GEN_2128; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2325 = 4'h5 == state ? plru1_12 : _GEN_2129; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2326 = 4'h5 == state ? plru1_13 : _GEN_2130; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2327 = 4'h5 == state ? plru1_14 : _GEN_2131; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2328 = 4'h5 == state ? plru1_15 : _GEN_2132; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2329 = 4'h5 == state ? plru1_16 : _GEN_2133; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2330 = 4'h5 == state ? plru1_17 : _GEN_2134; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2331 = 4'h5 == state ? plru1_18 : _GEN_2135; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2332 = 4'h5 == state ? plru1_19 : _GEN_2136; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2333 = 4'h5 == state ? plru1_20 : _GEN_2137; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2334 = 4'h5 == state ? plru1_21 : _GEN_2138; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2335 = 4'h5 == state ? plru1_22 : _GEN_2139; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2336 = 4'h5 == state ? plru1_23 : _GEN_2140; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2337 = 4'h5 == state ? plru1_24 : _GEN_2141; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2338 = 4'h5 == state ? plru1_25 : _GEN_2142; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2339 = 4'h5 == state ? plru1_26 : _GEN_2143; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2340 = 4'h5 == state ? plru1_27 : _GEN_2144; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2341 = 4'h5 == state ? plru1_28 : _GEN_2145; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2342 = 4'h5 == state ? plru1_29 : _GEN_2146; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2343 = 4'h5 == state ? plru1_30 : _GEN_2147; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2344 = 4'h5 == state ? plru1_31 : _GEN_2148; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2345 = 4'h5 == state ? plru1_32 : _GEN_2149; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2346 = 4'h5 == state ? plru1_33 : _GEN_2150; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2347 = 4'h5 == state ? plru1_34 : _GEN_2151; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2348 = 4'h5 == state ? plru1_35 : _GEN_2152; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2349 = 4'h5 == state ? plru1_36 : _GEN_2153; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2350 = 4'h5 == state ? plru1_37 : _GEN_2154; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2351 = 4'h5 == state ? plru1_38 : _GEN_2155; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2352 = 4'h5 == state ? plru1_39 : _GEN_2156; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2353 = 4'h5 == state ? plru1_40 : _GEN_2157; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2354 = 4'h5 == state ? plru1_41 : _GEN_2158; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2355 = 4'h5 == state ? plru1_42 : _GEN_2159; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2356 = 4'h5 == state ? plru1_43 : _GEN_2160; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2357 = 4'h5 == state ? plru1_44 : _GEN_2161; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2358 = 4'h5 == state ? plru1_45 : _GEN_2162; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2359 = 4'h5 == state ? plru1_46 : _GEN_2163; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2360 = 4'h5 == state ? plru1_47 : _GEN_2164; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2361 = 4'h5 == state ? plru1_48 : _GEN_2165; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2362 = 4'h5 == state ? plru1_49 : _GEN_2166; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2363 = 4'h5 == state ? plru1_50 : _GEN_2167; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2364 = 4'h5 == state ? plru1_51 : _GEN_2168; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2365 = 4'h5 == state ? plru1_52 : _GEN_2169; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2366 = 4'h5 == state ? plru1_53 : _GEN_2170; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2367 = 4'h5 == state ? plru1_54 : _GEN_2171; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2368 = 4'h5 == state ? plru1_55 : _GEN_2172; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2369 = 4'h5 == state ? plru1_56 : _GEN_2173; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2370 = 4'h5 == state ? plru1_57 : _GEN_2174; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2371 = 4'h5 == state ? plru1_58 : _GEN_2175; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2372 = 4'h5 == state ? plru1_59 : _GEN_2176; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2373 = 4'h5 == state ? plru1_60 : _GEN_2177; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2374 = 4'h5 == state ? plru1_61 : _GEN_2178; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2375 = 4'h5 == state ? plru1_62 : _GEN_2179; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2376 = 4'h5 == state ? plru1_63 : _GEN_2180; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2377 = 4'h5 == state ? plru2_0 : _GEN_2181; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2378 = 4'h5 == state ? plru2_1 : _GEN_2182; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2379 = 4'h5 == state ? plru2_2 : _GEN_2183; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2380 = 4'h5 == state ? plru2_3 : _GEN_2184; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2381 = 4'h5 == state ? plru2_4 : _GEN_2185; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2382 = 4'h5 == state ? plru2_5 : _GEN_2186; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2383 = 4'h5 == state ? plru2_6 : _GEN_2187; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2384 = 4'h5 == state ? plru2_7 : _GEN_2188; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2385 = 4'h5 == state ? plru2_8 : _GEN_2189; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2386 = 4'h5 == state ? plru2_9 : _GEN_2190; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2387 = 4'h5 == state ? plru2_10 : _GEN_2191; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2388 = 4'h5 == state ? plru2_11 : _GEN_2192; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2389 = 4'h5 == state ? plru2_12 : _GEN_2193; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2390 = 4'h5 == state ? plru2_13 : _GEN_2194; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2391 = 4'h5 == state ? plru2_14 : _GEN_2195; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2392 = 4'h5 == state ? plru2_15 : _GEN_2196; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2393 = 4'h5 == state ? plru2_16 : _GEN_2197; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2394 = 4'h5 == state ? plru2_17 : _GEN_2198; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2395 = 4'h5 == state ? plru2_18 : _GEN_2199; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2396 = 4'h5 == state ? plru2_19 : _GEN_2200; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2397 = 4'h5 == state ? plru2_20 : _GEN_2201; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2398 = 4'h5 == state ? plru2_21 : _GEN_2202; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2399 = 4'h5 == state ? plru2_22 : _GEN_2203; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2400 = 4'h5 == state ? plru2_23 : _GEN_2204; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2401 = 4'h5 == state ? plru2_24 : _GEN_2205; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2402 = 4'h5 == state ? plru2_25 : _GEN_2206; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2403 = 4'h5 == state ? plru2_26 : _GEN_2207; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2404 = 4'h5 == state ? plru2_27 : _GEN_2208; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2405 = 4'h5 == state ? plru2_28 : _GEN_2209; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2406 = 4'h5 == state ? plru2_29 : _GEN_2210; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2407 = 4'h5 == state ? plru2_30 : _GEN_2211; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2408 = 4'h5 == state ? plru2_31 : _GEN_2212; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2409 = 4'h5 == state ? plru2_32 : _GEN_2213; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2410 = 4'h5 == state ? plru2_33 : _GEN_2214; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2411 = 4'h5 == state ? plru2_34 : _GEN_2215; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2412 = 4'h5 == state ? plru2_35 : _GEN_2216; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2413 = 4'h5 == state ? plru2_36 : _GEN_2217; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2414 = 4'h5 == state ? plru2_37 : _GEN_2218; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2415 = 4'h5 == state ? plru2_38 : _GEN_2219; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2416 = 4'h5 == state ? plru2_39 : _GEN_2220; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2417 = 4'h5 == state ? plru2_40 : _GEN_2221; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2418 = 4'h5 == state ? plru2_41 : _GEN_2222; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2419 = 4'h5 == state ? plru2_42 : _GEN_2223; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2420 = 4'h5 == state ? plru2_43 : _GEN_2224; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2421 = 4'h5 == state ? plru2_44 : _GEN_2225; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2422 = 4'h5 == state ? plru2_45 : _GEN_2226; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2423 = 4'h5 == state ? plru2_46 : _GEN_2227; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2424 = 4'h5 == state ? plru2_47 : _GEN_2228; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2425 = 4'h5 == state ? plru2_48 : _GEN_2229; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2426 = 4'h5 == state ? plru2_49 : _GEN_2230; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2427 = 4'h5 == state ? plru2_50 : _GEN_2231; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2428 = 4'h5 == state ? plru2_51 : _GEN_2232; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2429 = 4'h5 == state ? plru2_52 : _GEN_2233; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2430 = 4'h5 == state ? plru2_53 : _GEN_2234; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2431 = 4'h5 == state ? plru2_54 : _GEN_2235; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2432 = 4'h5 == state ? plru2_55 : _GEN_2236; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2433 = 4'h5 == state ? plru2_56 : _GEN_2237; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2434 = 4'h5 == state ? plru2_57 : _GEN_2238; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2435 = 4'h5 == state ? plru2_58 : _GEN_2239; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2436 = 4'h5 == state ? plru2_59 : _GEN_2240; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2437 = 4'h5 == state ? plru2_60 : _GEN_2241; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2438 = 4'h5 == state ? plru2_61 : _GEN_2242; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2439 = 4'h5 == state ? plru2_62 : _GEN_2243; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2440 = 4'h5 == state ? plru2_63 : _GEN_2244; // @[Cache.scala 318:18 133:22]
  wire [63:0] _GEN_2441 = 4'h5 == state ? 64'h0 : _GEN_2246; // @[Cache.scala 318:18 289:22]
  wire [3:0] _GEN_2442 = 4'h4 == state ? _GEN_1534 : _GEN_2247; // @[Cache.scala 318:18]
  wire  _GEN_2444 = 4'h4 == state ? plru0_0 : _GEN_2249; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2445 = 4'h4 == state ? plru0_1 : _GEN_2250; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2446 = 4'h4 == state ? plru0_2 : _GEN_2251; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2447 = 4'h4 == state ? plru0_3 : _GEN_2252; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2448 = 4'h4 == state ? plru0_4 : _GEN_2253; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2449 = 4'h4 == state ? plru0_5 : _GEN_2254; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2450 = 4'h4 == state ? plru0_6 : _GEN_2255; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2451 = 4'h4 == state ? plru0_7 : _GEN_2256; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2452 = 4'h4 == state ? plru0_8 : _GEN_2257; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2453 = 4'h4 == state ? plru0_9 : _GEN_2258; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2454 = 4'h4 == state ? plru0_10 : _GEN_2259; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2455 = 4'h4 == state ? plru0_11 : _GEN_2260; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2456 = 4'h4 == state ? plru0_12 : _GEN_2261; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2457 = 4'h4 == state ? plru0_13 : _GEN_2262; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2458 = 4'h4 == state ? plru0_14 : _GEN_2263; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2459 = 4'h4 == state ? plru0_15 : _GEN_2264; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2460 = 4'h4 == state ? plru0_16 : _GEN_2265; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2461 = 4'h4 == state ? plru0_17 : _GEN_2266; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2462 = 4'h4 == state ? plru0_18 : _GEN_2267; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2463 = 4'h4 == state ? plru0_19 : _GEN_2268; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2464 = 4'h4 == state ? plru0_20 : _GEN_2269; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2465 = 4'h4 == state ? plru0_21 : _GEN_2270; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2466 = 4'h4 == state ? plru0_22 : _GEN_2271; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2467 = 4'h4 == state ? plru0_23 : _GEN_2272; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2468 = 4'h4 == state ? plru0_24 : _GEN_2273; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2469 = 4'h4 == state ? plru0_25 : _GEN_2274; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2470 = 4'h4 == state ? plru0_26 : _GEN_2275; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2471 = 4'h4 == state ? plru0_27 : _GEN_2276; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2472 = 4'h4 == state ? plru0_28 : _GEN_2277; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2473 = 4'h4 == state ? plru0_29 : _GEN_2278; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2474 = 4'h4 == state ? plru0_30 : _GEN_2279; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2475 = 4'h4 == state ? plru0_31 : _GEN_2280; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2476 = 4'h4 == state ? plru0_32 : _GEN_2281; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2477 = 4'h4 == state ? plru0_33 : _GEN_2282; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2478 = 4'h4 == state ? plru0_34 : _GEN_2283; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2479 = 4'h4 == state ? plru0_35 : _GEN_2284; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2480 = 4'h4 == state ? plru0_36 : _GEN_2285; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2481 = 4'h4 == state ? plru0_37 : _GEN_2286; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2482 = 4'h4 == state ? plru0_38 : _GEN_2287; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2483 = 4'h4 == state ? plru0_39 : _GEN_2288; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2484 = 4'h4 == state ? plru0_40 : _GEN_2289; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2485 = 4'h4 == state ? plru0_41 : _GEN_2290; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2486 = 4'h4 == state ? plru0_42 : _GEN_2291; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2487 = 4'h4 == state ? plru0_43 : _GEN_2292; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2488 = 4'h4 == state ? plru0_44 : _GEN_2293; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2489 = 4'h4 == state ? plru0_45 : _GEN_2294; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2490 = 4'h4 == state ? plru0_46 : _GEN_2295; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2491 = 4'h4 == state ? plru0_47 : _GEN_2296; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2492 = 4'h4 == state ? plru0_48 : _GEN_2297; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2493 = 4'h4 == state ? plru0_49 : _GEN_2298; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2494 = 4'h4 == state ? plru0_50 : _GEN_2299; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2495 = 4'h4 == state ? plru0_51 : _GEN_2300; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2496 = 4'h4 == state ? plru0_52 : _GEN_2301; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2497 = 4'h4 == state ? plru0_53 : _GEN_2302; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2498 = 4'h4 == state ? plru0_54 : _GEN_2303; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2499 = 4'h4 == state ? plru0_55 : _GEN_2304; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2500 = 4'h4 == state ? plru0_56 : _GEN_2305; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2501 = 4'h4 == state ? plru0_57 : _GEN_2306; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2502 = 4'h4 == state ? plru0_58 : _GEN_2307; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2503 = 4'h4 == state ? plru0_59 : _GEN_2308; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2504 = 4'h4 == state ? plru0_60 : _GEN_2309; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2505 = 4'h4 == state ? plru0_61 : _GEN_2310; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2506 = 4'h4 == state ? plru0_62 : _GEN_2311; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2507 = 4'h4 == state ? plru0_63 : _GEN_2312; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2508 = 4'h4 == state ? plru1_0 : _GEN_2313; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2509 = 4'h4 == state ? plru1_1 : _GEN_2314; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2510 = 4'h4 == state ? plru1_2 : _GEN_2315; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2511 = 4'h4 == state ? plru1_3 : _GEN_2316; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2512 = 4'h4 == state ? plru1_4 : _GEN_2317; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2513 = 4'h4 == state ? plru1_5 : _GEN_2318; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2514 = 4'h4 == state ? plru1_6 : _GEN_2319; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2515 = 4'h4 == state ? plru1_7 : _GEN_2320; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2516 = 4'h4 == state ? plru1_8 : _GEN_2321; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2517 = 4'h4 == state ? plru1_9 : _GEN_2322; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2518 = 4'h4 == state ? plru1_10 : _GEN_2323; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2519 = 4'h4 == state ? plru1_11 : _GEN_2324; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2520 = 4'h4 == state ? plru1_12 : _GEN_2325; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2521 = 4'h4 == state ? plru1_13 : _GEN_2326; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2522 = 4'h4 == state ? plru1_14 : _GEN_2327; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2523 = 4'h4 == state ? plru1_15 : _GEN_2328; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2524 = 4'h4 == state ? plru1_16 : _GEN_2329; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2525 = 4'h4 == state ? plru1_17 : _GEN_2330; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2526 = 4'h4 == state ? plru1_18 : _GEN_2331; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2527 = 4'h4 == state ? plru1_19 : _GEN_2332; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2528 = 4'h4 == state ? plru1_20 : _GEN_2333; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2529 = 4'h4 == state ? plru1_21 : _GEN_2334; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2530 = 4'h4 == state ? plru1_22 : _GEN_2335; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2531 = 4'h4 == state ? plru1_23 : _GEN_2336; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2532 = 4'h4 == state ? plru1_24 : _GEN_2337; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2533 = 4'h4 == state ? plru1_25 : _GEN_2338; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2534 = 4'h4 == state ? plru1_26 : _GEN_2339; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2535 = 4'h4 == state ? plru1_27 : _GEN_2340; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2536 = 4'h4 == state ? plru1_28 : _GEN_2341; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2537 = 4'h4 == state ? plru1_29 : _GEN_2342; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2538 = 4'h4 == state ? plru1_30 : _GEN_2343; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2539 = 4'h4 == state ? plru1_31 : _GEN_2344; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2540 = 4'h4 == state ? plru1_32 : _GEN_2345; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2541 = 4'h4 == state ? plru1_33 : _GEN_2346; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2542 = 4'h4 == state ? plru1_34 : _GEN_2347; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2543 = 4'h4 == state ? plru1_35 : _GEN_2348; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2544 = 4'h4 == state ? plru1_36 : _GEN_2349; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2545 = 4'h4 == state ? plru1_37 : _GEN_2350; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2546 = 4'h4 == state ? plru1_38 : _GEN_2351; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2547 = 4'h4 == state ? plru1_39 : _GEN_2352; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2548 = 4'h4 == state ? plru1_40 : _GEN_2353; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2549 = 4'h4 == state ? plru1_41 : _GEN_2354; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2550 = 4'h4 == state ? plru1_42 : _GEN_2355; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2551 = 4'h4 == state ? plru1_43 : _GEN_2356; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2552 = 4'h4 == state ? plru1_44 : _GEN_2357; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2553 = 4'h4 == state ? plru1_45 : _GEN_2358; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2554 = 4'h4 == state ? plru1_46 : _GEN_2359; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2555 = 4'h4 == state ? plru1_47 : _GEN_2360; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2556 = 4'h4 == state ? plru1_48 : _GEN_2361; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2557 = 4'h4 == state ? plru1_49 : _GEN_2362; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2558 = 4'h4 == state ? plru1_50 : _GEN_2363; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2559 = 4'h4 == state ? plru1_51 : _GEN_2364; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2560 = 4'h4 == state ? plru1_52 : _GEN_2365; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2561 = 4'h4 == state ? plru1_53 : _GEN_2366; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2562 = 4'h4 == state ? plru1_54 : _GEN_2367; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2563 = 4'h4 == state ? plru1_55 : _GEN_2368; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2564 = 4'h4 == state ? plru1_56 : _GEN_2369; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2565 = 4'h4 == state ? plru1_57 : _GEN_2370; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2566 = 4'h4 == state ? plru1_58 : _GEN_2371; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2567 = 4'h4 == state ? plru1_59 : _GEN_2372; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2568 = 4'h4 == state ? plru1_60 : _GEN_2373; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2569 = 4'h4 == state ? plru1_61 : _GEN_2374; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2570 = 4'h4 == state ? plru1_62 : _GEN_2375; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2571 = 4'h4 == state ? plru1_63 : _GEN_2376; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2572 = 4'h4 == state ? plru2_0 : _GEN_2377; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2573 = 4'h4 == state ? plru2_1 : _GEN_2378; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2574 = 4'h4 == state ? plru2_2 : _GEN_2379; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2575 = 4'h4 == state ? plru2_3 : _GEN_2380; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2576 = 4'h4 == state ? plru2_4 : _GEN_2381; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2577 = 4'h4 == state ? plru2_5 : _GEN_2382; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2578 = 4'h4 == state ? plru2_6 : _GEN_2383; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2579 = 4'h4 == state ? plru2_7 : _GEN_2384; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2580 = 4'h4 == state ? plru2_8 : _GEN_2385; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2581 = 4'h4 == state ? plru2_9 : _GEN_2386; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2582 = 4'h4 == state ? plru2_10 : _GEN_2387; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2583 = 4'h4 == state ? plru2_11 : _GEN_2388; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2584 = 4'h4 == state ? plru2_12 : _GEN_2389; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2585 = 4'h4 == state ? plru2_13 : _GEN_2390; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2586 = 4'h4 == state ? plru2_14 : _GEN_2391; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2587 = 4'h4 == state ? plru2_15 : _GEN_2392; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2588 = 4'h4 == state ? plru2_16 : _GEN_2393; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2589 = 4'h4 == state ? plru2_17 : _GEN_2394; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2590 = 4'h4 == state ? plru2_18 : _GEN_2395; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2591 = 4'h4 == state ? plru2_19 : _GEN_2396; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2592 = 4'h4 == state ? plru2_20 : _GEN_2397; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2593 = 4'h4 == state ? plru2_21 : _GEN_2398; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2594 = 4'h4 == state ? plru2_22 : _GEN_2399; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2595 = 4'h4 == state ? plru2_23 : _GEN_2400; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2596 = 4'h4 == state ? plru2_24 : _GEN_2401; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2597 = 4'h4 == state ? plru2_25 : _GEN_2402; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2598 = 4'h4 == state ? plru2_26 : _GEN_2403; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2599 = 4'h4 == state ? plru2_27 : _GEN_2404; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2600 = 4'h4 == state ? plru2_28 : _GEN_2405; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2601 = 4'h4 == state ? plru2_29 : _GEN_2406; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2602 = 4'h4 == state ? plru2_30 : _GEN_2407; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2603 = 4'h4 == state ? plru2_31 : _GEN_2408; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2604 = 4'h4 == state ? plru2_32 : _GEN_2409; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2605 = 4'h4 == state ? plru2_33 : _GEN_2410; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2606 = 4'h4 == state ? plru2_34 : _GEN_2411; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2607 = 4'h4 == state ? plru2_35 : _GEN_2412; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2608 = 4'h4 == state ? plru2_36 : _GEN_2413; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2609 = 4'h4 == state ? plru2_37 : _GEN_2414; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2610 = 4'h4 == state ? plru2_38 : _GEN_2415; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2611 = 4'h4 == state ? plru2_39 : _GEN_2416; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2612 = 4'h4 == state ? plru2_40 : _GEN_2417; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2613 = 4'h4 == state ? plru2_41 : _GEN_2418; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2614 = 4'h4 == state ? plru2_42 : _GEN_2419; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2615 = 4'h4 == state ? plru2_43 : _GEN_2420; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2616 = 4'h4 == state ? plru2_44 : _GEN_2421; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2617 = 4'h4 == state ? plru2_45 : _GEN_2422; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2618 = 4'h4 == state ? plru2_46 : _GEN_2423; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2619 = 4'h4 == state ? plru2_47 : _GEN_2424; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2620 = 4'h4 == state ? plru2_48 : _GEN_2425; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2621 = 4'h4 == state ? plru2_49 : _GEN_2426; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2622 = 4'h4 == state ? plru2_50 : _GEN_2427; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2623 = 4'h4 == state ? plru2_51 : _GEN_2428; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2624 = 4'h4 == state ? plru2_52 : _GEN_2429; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2625 = 4'h4 == state ? plru2_53 : _GEN_2430; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2626 = 4'h4 == state ? plru2_54 : _GEN_2431; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2627 = 4'h4 == state ? plru2_55 : _GEN_2432; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2628 = 4'h4 == state ? plru2_56 : _GEN_2433; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2629 = 4'h4 == state ? plru2_57 : _GEN_2434; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2630 = 4'h4 == state ? plru2_58 : _GEN_2435; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2631 = 4'h4 == state ? plru2_59 : _GEN_2436; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2632 = 4'h4 == state ? plru2_60 : _GEN_2437; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2633 = 4'h4 == state ? plru2_61 : _GEN_2438; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2634 = 4'h4 == state ? plru2_62 : _GEN_2439; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2635 = 4'h4 == state ? plru2_63 : _GEN_2440; // @[Cache.scala 318:18 133:22]
  wire [63:0] _GEN_2636 = 4'h4 == state ? 64'h0 : _GEN_2441; // @[Cache.scala 318:18 289:22]
  wire  _GEN_2637 = 4'h3 == state ? _GEN_994 : pipeline_ready; // @[Cache.scala 318:18]
  wire [5:0] _GEN_2639 = 4'h3 == state ? _GEN_996 : _GEN_3; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2640 = 4'h3 == state ? _GEN_997 : 128'h0; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2641 = 4'h3 == state ? _GEN_998 : 21'h0; // @[Cache.scala 114:16 318:18]
  wire  _GEN_2643 = 4'h3 == state ? _GEN_1001 : pipeline_ready; // @[Cache.scala 318:18]
  wire [5:0] _GEN_2645 = 4'h3 == state ? _GEN_1003 : _GEN_3; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2646 = 4'h3 == state ? _GEN_1004 : 128'h0; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2647 = 4'h3 == state ? _GEN_1005 : 21'h0; // @[Cache.scala 114:16 318:18]
  wire  _GEN_2649 = 4'h3 == state ? _GEN_1008 : pipeline_ready; // @[Cache.scala 318:18]
  wire [5:0] _GEN_2651 = 4'h3 == state ? _GEN_1010 : _GEN_3; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2652 = 4'h3 == state ? _GEN_1011 : 128'h0; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2653 = 4'h3 == state ? _GEN_1012 : 21'h0; // @[Cache.scala 114:16 318:18]
  wire  _GEN_2655 = 4'h3 == state ? _GEN_1015 : pipeline_ready; // @[Cache.scala 318:18]
  wire [5:0] _GEN_2657 = 4'h3 == state ? _GEN_1017 : _GEN_3; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2658 = 4'h3 == state ? _GEN_1018 : 128'h0; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2659 = 4'h3 == state ? _GEN_1019 : 21'h0; // @[Cache.scala 114:16 318:18]
  wire [3:0] _GEN_2661 = 4'h3 == state ? _GEN_1341 : _GEN_2442; // @[Cache.scala 318:18]
  wire  _GEN_2662 = 4'h3 == state ? _GEN_1342 : _GEN_2444; // @[Cache.scala 318:18]
  wire  _GEN_2663 = 4'h3 == state ? _GEN_1343 : _GEN_2445; // @[Cache.scala 318:18]
  wire  _GEN_2664 = 4'h3 == state ? _GEN_1344 : _GEN_2446; // @[Cache.scala 318:18]
  wire  _GEN_2665 = 4'h3 == state ? _GEN_1345 : _GEN_2447; // @[Cache.scala 318:18]
  wire  _GEN_2666 = 4'h3 == state ? _GEN_1346 : _GEN_2448; // @[Cache.scala 318:18]
  wire  _GEN_2667 = 4'h3 == state ? _GEN_1347 : _GEN_2449; // @[Cache.scala 318:18]
  wire  _GEN_2668 = 4'h3 == state ? _GEN_1348 : _GEN_2450; // @[Cache.scala 318:18]
  wire  _GEN_2669 = 4'h3 == state ? _GEN_1349 : _GEN_2451; // @[Cache.scala 318:18]
  wire  _GEN_2670 = 4'h3 == state ? _GEN_1350 : _GEN_2452; // @[Cache.scala 318:18]
  wire  _GEN_2671 = 4'h3 == state ? _GEN_1351 : _GEN_2453; // @[Cache.scala 318:18]
  wire  _GEN_2672 = 4'h3 == state ? _GEN_1352 : _GEN_2454; // @[Cache.scala 318:18]
  wire  _GEN_2673 = 4'h3 == state ? _GEN_1353 : _GEN_2455; // @[Cache.scala 318:18]
  wire  _GEN_2674 = 4'h3 == state ? _GEN_1354 : _GEN_2456; // @[Cache.scala 318:18]
  wire  _GEN_2675 = 4'h3 == state ? _GEN_1355 : _GEN_2457; // @[Cache.scala 318:18]
  wire  _GEN_2676 = 4'h3 == state ? _GEN_1356 : _GEN_2458; // @[Cache.scala 318:18]
  wire  _GEN_2677 = 4'h3 == state ? _GEN_1357 : _GEN_2459; // @[Cache.scala 318:18]
  wire  _GEN_2678 = 4'h3 == state ? _GEN_1358 : _GEN_2460; // @[Cache.scala 318:18]
  wire  _GEN_2679 = 4'h3 == state ? _GEN_1359 : _GEN_2461; // @[Cache.scala 318:18]
  wire  _GEN_2680 = 4'h3 == state ? _GEN_1360 : _GEN_2462; // @[Cache.scala 318:18]
  wire  _GEN_2681 = 4'h3 == state ? _GEN_1361 : _GEN_2463; // @[Cache.scala 318:18]
  wire  _GEN_2682 = 4'h3 == state ? _GEN_1362 : _GEN_2464; // @[Cache.scala 318:18]
  wire  _GEN_2683 = 4'h3 == state ? _GEN_1363 : _GEN_2465; // @[Cache.scala 318:18]
  wire  _GEN_2684 = 4'h3 == state ? _GEN_1364 : _GEN_2466; // @[Cache.scala 318:18]
  wire  _GEN_2685 = 4'h3 == state ? _GEN_1365 : _GEN_2467; // @[Cache.scala 318:18]
  wire  _GEN_2686 = 4'h3 == state ? _GEN_1366 : _GEN_2468; // @[Cache.scala 318:18]
  wire  _GEN_2687 = 4'h3 == state ? _GEN_1367 : _GEN_2469; // @[Cache.scala 318:18]
  wire  _GEN_2688 = 4'h3 == state ? _GEN_1368 : _GEN_2470; // @[Cache.scala 318:18]
  wire  _GEN_2689 = 4'h3 == state ? _GEN_1369 : _GEN_2471; // @[Cache.scala 318:18]
  wire  _GEN_2690 = 4'h3 == state ? _GEN_1370 : _GEN_2472; // @[Cache.scala 318:18]
  wire  _GEN_2691 = 4'h3 == state ? _GEN_1371 : _GEN_2473; // @[Cache.scala 318:18]
  wire  _GEN_2692 = 4'h3 == state ? _GEN_1372 : _GEN_2474; // @[Cache.scala 318:18]
  wire  _GEN_2693 = 4'h3 == state ? _GEN_1373 : _GEN_2475; // @[Cache.scala 318:18]
  wire  _GEN_2694 = 4'h3 == state ? _GEN_1374 : _GEN_2476; // @[Cache.scala 318:18]
  wire  _GEN_2695 = 4'h3 == state ? _GEN_1375 : _GEN_2477; // @[Cache.scala 318:18]
  wire  _GEN_2696 = 4'h3 == state ? _GEN_1376 : _GEN_2478; // @[Cache.scala 318:18]
  wire  _GEN_2697 = 4'h3 == state ? _GEN_1377 : _GEN_2479; // @[Cache.scala 318:18]
  wire  _GEN_2698 = 4'h3 == state ? _GEN_1378 : _GEN_2480; // @[Cache.scala 318:18]
  wire  _GEN_2699 = 4'h3 == state ? _GEN_1379 : _GEN_2481; // @[Cache.scala 318:18]
  wire  _GEN_2700 = 4'h3 == state ? _GEN_1380 : _GEN_2482; // @[Cache.scala 318:18]
  wire  _GEN_2701 = 4'h3 == state ? _GEN_1381 : _GEN_2483; // @[Cache.scala 318:18]
  wire  _GEN_2702 = 4'h3 == state ? _GEN_1382 : _GEN_2484; // @[Cache.scala 318:18]
  wire  _GEN_2703 = 4'h3 == state ? _GEN_1383 : _GEN_2485; // @[Cache.scala 318:18]
  wire  _GEN_2704 = 4'h3 == state ? _GEN_1384 : _GEN_2486; // @[Cache.scala 318:18]
  wire  _GEN_2705 = 4'h3 == state ? _GEN_1385 : _GEN_2487; // @[Cache.scala 318:18]
  wire  _GEN_2706 = 4'h3 == state ? _GEN_1386 : _GEN_2488; // @[Cache.scala 318:18]
  wire  _GEN_2707 = 4'h3 == state ? _GEN_1387 : _GEN_2489; // @[Cache.scala 318:18]
  wire  _GEN_2708 = 4'h3 == state ? _GEN_1388 : _GEN_2490; // @[Cache.scala 318:18]
  wire  _GEN_2709 = 4'h3 == state ? _GEN_1389 : _GEN_2491; // @[Cache.scala 318:18]
  wire  _GEN_2710 = 4'h3 == state ? _GEN_1390 : _GEN_2492; // @[Cache.scala 318:18]
  wire  _GEN_2711 = 4'h3 == state ? _GEN_1391 : _GEN_2493; // @[Cache.scala 318:18]
  wire  _GEN_2712 = 4'h3 == state ? _GEN_1392 : _GEN_2494; // @[Cache.scala 318:18]
  wire  _GEN_2713 = 4'h3 == state ? _GEN_1393 : _GEN_2495; // @[Cache.scala 318:18]
  wire  _GEN_2714 = 4'h3 == state ? _GEN_1394 : _GEN_2496; // @[Cache.scala 318:18]
  wire  _GEN_2715 = 4'h3 == state ? _GEN_1395 : _GEN_2497; // @[Cache.scala 318:18]
  wire  _GEN_2716 = 4'h3 == state ? _GEN_1396 : _GEN_2498; // @[Cache.scala 318:18]
  wire  _GEN_2717 = 4'h3 == state ? _GEN_1397 : _GEN_2499; // @[Cache.scala 318:18]
  wire  _GEN_2718 = 4'h3 == state ? _GEN_1398 : _GEN_2500; // @[Cache.scala 318:18]
  wire  _GEN_2719 = 4'h3 == state ? _GEN_1399 : _GEN_2501; // @[Cache.scala 318:18]
  wire  _GEN_2720 = 4'h3 == state ? _GEN_1400 : _GEN_2502; // @[Cache.scala 318:18]
  wire  _GEN_2721 = 4'h3 == state ? _GEN_1401 : _GEN_2503; // @[Cache.scala 318:18]
  wire  _GEN_2722 = 4'h3 == state ? _GEN_1402 : _GEN_2504; // @[Cache.scala 318:18]
  wire  _GEN_2723 = 4'h3 == state ? _GEN_1403 : _GEN_2505; // @[Cache.scala 318:18]
  wire  _GEN_2724 = 4'h3 == state ? _GEN_1404 : _GEN_2506; // @[Cache.scala 318:18]
  wire  _GEN_2725 = 4'h3 == state ? _GEN_1405 : _GEN_2507; // @[Cache.scala 318:18]
  wire  _GEN_2726 = 4'h3 == state ? _GEN_1406 : _GEN_2508; // @[Cache.scala 318:18]
  wire  _GEN_2727 = 4'h3 == state ? _GEN_1407 : _GEN_2509; // @[Cache.scala 318:18]
  wire  _GEN_2728 = 4'h3 == state ? _GEN_1408 : _GEN_2510; // @[Cache.scala 318:18]
  wire  _GEN_2729 = 4'h3 == state ? _GEN_1409 : _GEN_2511; // @[Cache.scala 318:18]
  wire  _GEN_2730 = 4'h3 == state ? _GEN_1410 : _GEN_2512; // @[Cache.scala 318:18]
  wire  _GEN_2731 = 4'h3 == state ? _GEN_1411 : _GEN_2513; // @[Cache.scala 318:18]
  wire  _GEN_2732 = 4'h3 == state ? _GEN_1412 : _GEN_2514; // @[Cache.scala 318:18]
  wire  _GEN_2733 = 4'h3 == state ? _GEN_1413 : _GEN_2515; // @[Cache.scala 318:18]
  wire  _GEN_2734 = 4'h3 == state ? _GEN_1414 : _GEN_2516; // @[Cache.scala 318:18]
  wire  _GEN_2735 = 4'h3 == state ? _GEN_1415 : _GEN_2517; // @[Cache.scala 318:18]
  wire  _GEN_2736 = 4'h3 == state ? _GEN_1416 : _GEN_2518; // @[Cache.scala 318:18]
  wire  _GEN_2737 = 4'h3 == state ? _GEN_1417 : _GEN_2519; // @[Cache.scala 318:18]
  wire  _GEN_2738 = 4'h3 == state ? _GEN_1418 : _GEN_2520; // @[Cache.scala 318:18]
  wire  _GEN_2739 = 4'h3 == state ? _GEN_1419 : _GEN_2521; // @[Cache.scala 318:18]
  wire  _GEN_2740 = 4'h3 == state ? _GEN_1420 : _GEN_2522; // @[Cache.scala 318:18]
  wire  _GEN_2741 = 4'h3 == state ? _GEN_1421 : _GEN_2523; // @[Cache.scala 318:18]
  wire  _GEN_2742 = 4'h3 == state ? _GEN_1422 : _GEN_2524; // @[Cache.scala 318:18]
  wire  _GEN_2743 = 4'h3 == state ? _GEN_1423 : _GEN_2525; // @[Cache.scala 318:18]
  wire  _GEN_2744 = 4'h3 == state ? _GEN_1424 : _GEN_2526; // @[Cache.scala 318:18]
  wire  _GEN_2745 = 4'h3 == state ? _GEN_1425 : _GEN_2527; // @[Cache.scala 318:18]
  wire  _GEN_2746 = 4'h3 == state ? _GEN_1426 : _GEN_2528; // @[Cache.scala 318:18]
  wire  _GEN_2747 = 4'h3 == state ? _GEN_1427 : _GEN_2529; // @[Cache.scala 318:18]
  wire  _GEN_2748 = 4'h3 == state ? _GEN_1428 : _GEN_2530; // @[Cache.scala 318:18]
  wire  _GEN_2749 = 4'h3 == state ? _GEN_1429 : _GEN_2531; // @[Cache.scala 318:18]
  wire  _GEN_2750 = 4'h3 == state ? _GEN_1430 : _GEN_2532; // @[Cache.scala 318:18]
  wire  _GEN_2751 = 4'h3 == state ? _GEN_1431 : _GEN_2533; // @[Cache.scala 318:18]
  wire  _GEN_2752 = 4'h3 == state ? _GEN_1432 : _GEN_2534; // @[Cache.scala 318:18]
  wire  _GEN_2753 = 4'h3 == state ? _GEN_1433 : _GEN_2535; // @[Cache.scala 318:18]
  wire  _GEN_2754 = 4'h3 == state ? _GEN_1434 : _GEN_2536; // @[Cache.scala 318:18]
  wire  _GEN_2755 = 4'h3 == state ? _GEN_1435 : _GEN_2537; // @[Cache.scala 318:18]
  wire  _GEN_2756 = 4'h3 == state ? _GEN_1436 : _GEN_2538; // @[Cache.scala 318:18]
  wire  _GEN_2757 = 4'h3 == state ? _GEN_1437 : _GEN_2539; // @[Cache.scala 318:18]
  wire  _GEN_2758 = 4'h3 == state ? _GEN_1438 : _GEN_2540; // @[Cache.scala 318:18]
  wire  _GEN_2759 = 4'h3 == state ? _GEN_1439 : _GEN_2541; // @[Cache.scala 318:18]
  wire  _GEN_2760 = 4'h3 == state ? _GEN_1440 : _GEN_2542; // @[Cache.scala 318:18]
  wire  _GEN_2761 = 4'h3 == state ? _GEN_1441 : _GEN_2543; // @[Cache.scala 318:18]
  wire  _GEN_2762 = 4'h3 == state ? _GEN_1442 : _GEN_2544; // @[Cache.scala 318:18]
  wire  _GEN_2763 = 4'h3 == state ? _GEN_1443 : _GEN_2545; // @[Cache.scala 318:18]
  wire  _GEN_2764 = 4'h3 == state ? _GEN_1444 : _GEN_2546; // @[Cache.scala 318:18]
  wire  _GEN_2765 = 4'h3 == state ? _GEN_1445 : _GEN_2547; // @[Cache.scala 318:18]
  wire  _GEN_2766 = 4'h3 == state ? _GEN_1446 : _GEN_2548; // @[Cache.scala 318:18]
  wire  _GEN_2767 = 4'h3 == state ? _GEN_1447 : _GEN_2549; // @[Cache.scala 318:18]
  wire  _GEN_2768 = 4'h3 == state ? _GEN_1448 : _GEN_2550; // @[Cache.scala 318:18]
  wire  _GEN_2769 = 4'h3 == state ? _GEN_1449 : _GEN_2551; // @[Cache.scala 318:18]
  wire  _GEN_2770 = 4'h3 == state ? _GEN_1450 : _GEN_2552; // @[Cache.scala 318:18]
  wire  _GEN_2771 = 4'h3 == state ? _GEN_1451 : _GEN_2553; // @[Cache.scala 318:18]
  wire  _GEN_2772 = 4'h3 == state ? _GEN_1452 : _GEN_2554; // @[Cache.scala 318:18]
  wire  _GEN_2773 = 4'h3 == state ? _GEN_1453 : _GEN_2555; // @[Cache.scala 318:18]
  wire  _GEN_2774 = 4'h3 == state ? _GEN_1454 : _GEN_2556; // @[Cache.scala 318:18]
  wire  _GEN_2775 = 4'h3 == state ? _GEN_1455 : _GEN_2557; // @[Cache.scala 318:18]
  wire  _GEN_2776 = 4'h3 == state ? _GEN_1456 : _GEN_2558; // @[Cache.scala 318:18]
  wire  _GEN_2777 = 4'h3 == state ? _GEN_1457 : _GEN_2559; // @[Cache.scala 318:18]
  wire  _GEN_2778 = 4'h3 == state ? _GEN_1458 : _GEN_2560; // @[Cache.scala 318:18]
  wire  _GEN_2779 = 4'h3 == state ? _GEN_1459 : _GEN_2561; // @[Cache.scala 318:18]
  wire  _GEN_2780 = 4'h3 == state ? _GEN_1460 : _GEN_2562; // @[Cache.scala 318:18]
  wire  _GEN_2781 = 4'h3 == state ? _GEN_1461 : _GEN_2563; // @[Cache.scala 318:18]
  wire  _GEN_2782 = 4'h3 == state ? _GEN_1462 : _GEN_2564; // @[Cache.scala 318:18]
  wire  _GEN_2783 = 4'h3 == state ? _GEN_1463 : _GEN_2565; // @[Cache.scala 318:18]
  wire  _GEN_2784 = 4'h3 == state ? _GEN_1464 : _GEN_2566; // @[Cache.scala 318:18]
  wire  _GEN_2785 = 4'h3 == state ? _GEN_1465 : _GEN_2567; // @[Cache.scala 318:18]
  wire  _GEN_2786 = 4'h3 == state ? _GEN_1466 : _GEN_2568; // @[Cache.scala 318:18]
  wire  _GEN_2787 = 4'h3 == state ? _GEN_1467 : _GEN_2569; // @[Cache.scala 318:18]
  wire  _GEN_2788 = 4'h3 == state ? _GEN_1468 : _GEN_2570; // @[Cache.scala 318:18]
  wire  _GEN_2789 = 4'h3 == state ? _GEN_1469 : _GEN_2571; // @[Cache.scala 318:18]
  wire  _GEN_2790 = 4'h3 == state ? _GEN_1470 : _GEN_2572; // @[Cache.scala 318:18]
  wire  _GEN_2791 = 4'h3 == state ? _GEN_1471 : _GEN_2573; // @[Cache.scala 318:18]
  wire  _GEN_2792 = 4'h3 == state ? _GEN_1472 : _GEN_2574; // @[Cache.scala 318:18]
  wire  _GEN_2793 = 4'h3 == state ? _GEN_1473 : _GEN_2575; // @[Cache.scala 318:18]
  wire  _GEN_2794 = 4'h3 == state ? _GEN_1474 : _GEN_2576; // @[Cache.scala 318:18]
  wire  _GEN_2795 = 4'h3 == state ? _GEN_1475 : _GEN_2577; // @[Cache.scala 318:18]
  wire  _GEN_2796 = 4'h3 == state ? _GEN_1476 : _GEN_2578; // @[Cache.scala 318:18]
  wire  _GEN_2797 = 4'h3 == state ? _GEN_1477 : _GEN_2579; // @[Cache.scala 318:18]
  wire  _GEN_2798 = 4'h3 == state ? _GEN_1478 : _GEN_2580; // @[Cache.scala 318:18]
  wire  _GEN_2799 = 4'h3 == state ? _GEN_1479 : _GEN_2581; // @[Cache.scala 318:18]
  wire  _GEN_2800 = 4'h3 == state ? _GEN_1480 : _GEN_2582; // @[Cache.scala 318:18]
  wire  _GEN_2801 = 4'h3 == state ? _GEN_1481 : _GEN_2583; // @[Cache.scala 318:18]
  wire  _GEN_2802 = 4'h3 == state ? _GEN_1482 : _GEN_2584; // @[Cache.scala 318:18]
  wire  _GEN_2803 = 4'h3 == state ? _GEN_1483 : _GEN_2585; // @[Cache.scala 318:18]
  wire  _GEN_2804 = 4'h3 == state ? _GEN_1484 : _GEN_2586; // @[Cache.scala 318:18]
  wire  _GEN_2805 = 4'h3 == state ? _GEN_1485 : _GEN_2587; // @[Cache.scala 318:18]
  wire  _GEN_2806 = 4'h3 == state ? _GEN_1486 : _GEN_2588; // @[Cache.scala 318:18]
  wire  _GEN_2807 = 4'h3 == state ? _GEN_1487 : _GEN_2589; // @[Cache.scala 318:18]
  wire  _GEN_2808 = 4'h3 == state ? _GEN_1488 : _GEN_2590; // @[Cache.scala 318:18]
  wire  _GEN_2809 = 4'h3 == state ? _GEN_1489 : _GEN_2591; // @[Cache.scala 318:18]
  wire  _GEN_2810 = 4'h3 == state ? _GEN_1490 : _GEN_2592; // @[Cache.scala 318:18]
  wire  _GEN_2811 = 4'h3 == state ? _GEN_1491 : _GEN_2593; // @[Cache.scala 318:18]
  wire  _GEN_2812 = 4'h3 == state ? _GEN_1492 : _GEN_2594; // @[Cache.scala 318:18]
  wire  _GEN_2813 = 4'h3 == state ? _GEN_1493 : _GEN_2595; // @[Cache.scala 318:18]
  wire  _GEN_2814 = 4'h3 == state ? _GEN_1494 : _GEN_2596; // @[Cache.scala 318:18]
  wire  _GEN_2815 = 4'h3 == state ? _GEN_1495 : _GEN_2597; // @[Cache.scala 318:18]
  wire  _GEN_2816 = 4'h3 == state ? _GEN_1496 : _GEN_2598; // @[Cache.scala 318:18]
  wire  _GEN_2817 = 4'h3 == state ? _GEN_1497 : _GEN_2599; // @[Cache.scala 318:18]
  wire  _GEN_2818 = 4'h3 == state ? _GEN_1498 : _GEN_2600; // @[Cache.scala 318:18]
  wire  _GEN_2819 = 4'h3 == state ? _GEN_1499 : _GEN_2601; // @[Cache.scala 318:18]
  wire  _GEN_2820 = 4'h3 == state ? _GEN_1500 : _GEN_2602; // @[Cache.scala 318:18]
  wire  _GEN_2821 = 4'h3 == state ? _GEN_1501 : _GEN_2603; // @[Cache.scala 318:18]
  wire  _GEN_2822 = 4'h3 == state ? _GEN_1502 : _GEN_2604; // @[Cache.scala 318:18]
  wire  _GEN_2823 = 4'h3 == state ? _GEN_1503 : _GEN_2605; // @[Cache.scala 318:18]
  wire  _GEN_2824 = 4'h3 == state ? _GEN_1504 : _GEN_2606; // @[Cache.scala 318:18]
  wire  _GEN_2825 = 4'h3 == state ? _GEN_1505 : _GEN_2607; // @[Cache.scala 318:18]
  wire  _GEN_2826 = 4'h3 == state ? _GEN_1506 : _GEN_2608; // @[Cache.scala 318:18]
  wire  _GEN_2827 = 4'h3 == state ? _GEN_1507 : _GEN_2609; // @[Cache.scala 318:18]
  wire  _GEN_2828 = 4'h3 == state ? _GEN_1508 : _GEN_2610; // @[Cache.scala 318:18]
  wire  _GEN_2829 = 4'h3 == state ? _GEN_1509 : _GEN_2611; // @[Cache.scala 318:18]
  wire  _GEN_2830 = 4'h3 == state ? _GEN_1510 : _GEN_2612; // @[Cache.scala 318:18]
  wire  _GEN_2831 = 4'h3 == state ? _GEN_1511 : _GEN_2613; // @[Cache.scala 318:18]
  wire  _GEN_2832 = 4'h3 == state ? _GEN_1512 : _GEN_2614; // @[Cache.scala 318:18]
  wire  _GEN_2833 = 4'h3 == state ? _GEN_1513 : _GEN_2615; // @[Cache.scala 318:18]
  wire  _GEN_2834 = 4'h3 == state ? _GEN_1514 : _GEN_2616; // @[Cache.scala 318:18]
  wire  _GEN_2835 = 4'h3 == state ? _GEN_1515 : _GEN_2617; // @[Cache.scala 318:18]
  wire  _GEN_2836 = 4'h3 == state ? _GEN_1516 : _GEN_2618; // @[Cache.scala 318:18]
  wire  _GEN_2837 = 4'h3 == state ? _GEN_1517 : _GEN_2619; // @[Cache.scala 318:18]
  wire  _GEN_2838 = 4'h3 == state ? _GEN_1518 : _GEN_2620; // @[Cache.scala 318:18]
  wire  _GEN_2839 = 4'h3 == state ? _GEN_1519 : _GEN_2621; // @[Cache.scala 318:18]
  wire  _GEN_2840 = 4'h3 == state ? _GEN_1520 : _GEN_2622; // @[Cache.scala 318:18]
  wire  _GEN_2841 = 4'h3 == state ? _GEN_1521 : _GEN_2623; // @[Cache.scala 318:18]
  wire  _GEN_2842 = 4'h3 == state ? _GEN_1522 : _GEN_2624; // @[Cache.scala 318:18]
  wire  _GEN_2843 = 4'h3 == state ? _GEN_1523 : _GEN_2625; // @[Cache.scala 318:18]
  wire  _GEN_2844 = 4'h3 == state ? _GEN_1524 : _GEN_2626; // @[Cache.scala 318:18]
  wire  _GEN_2845 = 4'h3 == state ? _GEN_1525 : _GEN_2627; // @[Cache.scala 318:18]
  wire  _GEN_2846 = 4'h3 == state ? _GEN_1526 : _GEN_2628; // @[Cache.scala 318:18]
  wire  _GEN_2847 = 4'h3 == state ? _GEN_1527 : _GEN_2629; // @[Cache.scala 318:18]
  wire  _GEN_2848 = 4'h3 == state ? _GEN_1528 : _GEN_2630; // @[Cache.scala 318:18]
  wire  _GEN_2849 = 4'h3 == state ? _GEN_1529 : _GEN_2631; // @[Cache.scala 318:18]
  wire  _GEN_2850 = 4'h3 == state ? _GEN_1530 : _GEN_2632; // @[Cache.scala 318:18]
  wire  _GEN_2851 = 4'h3 == state ? _GEN_1531 : _GEN_2633; // @[Cache.scala 318:18]
  wire  _GEN_2852 = 4'h3 == state ? _GEN_1532 : _GEN_2634; // @[Cache.scala 318:18]
  wire  _GEN_2853 = 4'h3 == state ? _GEN_1533 : _GEN_2635; // @[Cache.scala 318:18]
  wire [63:0] _GEN_2855 = 4'h3 == state ? 64'h0 : _GEN_2636; // @[Cache.scala 318:18 289:22]
  wire [3:0] _GEN_2858 = 4'h2 == state ? _GEN_992 : _GEN_2661; // @[Cache.scala 318:18]
  wire  _GEN_2859 = 4'h2 == state ? pipeline_ready : _GEN_2637; // @[Cache.scala 318:18]
  wire  _GEN_2860 = 4'h2 == state ? 1'h0 : 4'h3 == state & _T_325; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_2861 = 4'h2 == state ? _GEN_3 : _GEN_2639; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2862 = 4'h2 == state ? 128'h0 : _GEN_2640; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2863 = 4'h2 == state ? 21'h0 : _GEN_2641; // @[Cache.scala 114:16 318:18]
  wire  _GEN_2865 = 4'h2 == state ? pipeline_ready : _GEN_2643; // @[Cache.scala 318:18]
  wire  _GEN_2866 = 4'h2 == state ? 1'h0 : 4'h3 == state & _T_389; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_2867 = 4'h2 == state ? _GEN_3 : _GEN_2645; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2868 = 4'h2 == state ? 128'h0 : _GEN_2646; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2869 = 4'h2 == state ? 21'h0 : _GEN_2647; // @[Cache.scala 114:16 318:18]
  wire  _GEN_2871 = 4'h2 == state ? pipeline_ready : _GEN_2649; // @[Cache.scala 318:18]
  wire  _GEN_2872 = 4'h2 == state ? 1'h0 : 4'h3 == state & _T_453; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_2873 = 4'h2 == state ? _GEN_3 : _GEN_2651; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2874 = 4'h2 == state ? 128'h0 : _GEN_2652; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2875 = 4'h2 == state ? 21'h0 : _GEN_2653; // @[Cache.scala 114:16 318:18]
  wire  _GEN_2877 = 4'h2 == state ? pipeline_ready : _GEN_2655; // @[Cache.scala 318:18]
  wire  _GEN_2878 = 4'h2 == state ? 1'h0 : 4'h3 == state & _T_517; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_2879 = 4'h2 == state ? _GEN_3 : _GEN_2657; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2880 = 4'h2 == state ? 128'h0 : _GEN_2658; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2881 = 4'h2 == state ? 21'h0 : _GEN_2659; // @[Cache.scala 114:16 318:18]
  wire [63:0] _GEN_3076 = 4'h2 == state ? 64'h0 : _GEN_2855; // @[Cache.scala 318:18 289:22]
  wire [3:0] _GEN_3077 = 4'h1 == state ? _GEN_986 : _GEN_2858; // @[Cache.scala 318:18]
  wire  _GEN_3080 = 4'h1 == state ? pipeline_ready : _GEN_2859; // @[Cache.scala 318:18]
  wire  _GEN_3081 = 4'h1 == state ? 1'h0 : _GEN_2860; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_3082 = 4'h1 == state ? _GEN_3 : _GEN_2861; // @[Cache.scala 318:18]
  wire [127:0] _GEN_3083 = 4'h1 == state ? 128'h0 : _GEN_2862; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_3084 = 4'h1 == state ? 21'h0 : _GEN_2863; // @[Cache.scala 114:16 318:18]
  wire  _GEN_3086 = 4'h1 == state ? pipeline_ready : _GEN_2865; // @[Cache.scala 318:18]
  wire  _GEN_3087 = 4'h1 == state ? 1'h0 : _GEN_2866; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_3088 = 4'h1 == state ? _GEN_3 : _GEN_2867; // @[Cache.scala 318:18]
  wire [127:0] _GEN_3089 = 4'h1 == state ? 128'h0 : _GEN_2868; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_3090 = 4'h1 == state ? 21'h0 : _GEN_2869; // @[Cache.scala 114:16 318:18]
  wire  _GEN_3092 = 4'h1 == state ? pipeline_ready : _GEN_2871; // @[Cache.scala 318:18]
  wire  _GEN_3093 = 4'h1 == state ? 1'h0 : _GEN_2872; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_3094 = 4'h1 == state ? _GEN_3 : _GEN_2873; // @[Cache.scala 318:18]
  wire [127:0] _GEN_3095 = 4'h1 == state ? 128'h0 : _GEN_2874; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_3096 = 4'h1 == state ? 21'h0 : _GEN_2875; // @[Cache.scala 114:16 318:18]
  wire  _GEN_3098 = 4'h1 == state ? pipeline_ready : _GEN_2877; // @[Cache.scala 318:18]
  wire  _GEN_3099 = 4'h1 == state ? 1'h0 : _GEN_2878; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_3100 = 4'h1 == state ? _GEN_3 : _GEN_2879; // @[Cache.scala 318:18]
  wire [127:0] _GEN_3101 = 4'h1 == state ? 128'h0 : _GEN_2880; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_3102 = 4'h1 == state ? 21'h0 : _GEN_2881; // @[Cache.scala 114:16 318:18]
  wire [63:0] _GEN_3297 = 4'h1 == state ? 64'h0 : _GEN_3076; // @[Cache.scala 318:18 289:22]
  wire  _T_610 = state == 4'h1; // @[Cache.scala 540:27]
  wire  _T_611 = state == 4'h4; // @[Cache.scala 541:27]
  wire  _T_612 = state == 4'h1 | _T_611; // @[Cache.scala 540:45]
  wire  _T_613 = state == 4'h5; // @[Cache.scala 542:27]
  wire [31:0] _T_622 = {s2_addr[31:4],4'h0}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3536 = _T_610 ? _T_622 : 32'h0; // @[Cache.scala 546:21 547:33 548:23]
  wire [31:0] _T_625 = {1'h1,s2_reg_tag_r,s2_idx,4'h0}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_3539 = _T_611 ? s2_reg_dat_w[63:0] : 64'h0; // @[Cache.scala 561:22 562:34 563:24]
  wire  _T_653 = state == 4'h6; // @[Cache.scala 584:28]
  ysyx_210128_Sram sram_0 ( // @[Cache.scala 89:22]
    .clock(sram_0_clock),
    .io_en(sram_0_io_en),
    .io_wen(sram_0_io_wen),
    .io_addr(sram_0_io_addr),
    .io_wdata(sram_0_io_wdata),
    .io_rdata(sram_0_io_rdata)
  );
  ysyx_210128_Sram sram_1 ( // @[Cache.scala 89:22]
    .clock(sram_1_clock),
    .io_en(sram_1_io_en),
    .io_wen(sram_1_io_wen),
    .io_addr(sram_1_io_addr),
    .io_wdata(sram_1_io_wdata),
    .io_rdata(sram_1_io_rdata)
  );
  ysyx_210128_Sram sram_2 ( // @[Cache.scala 89:22]
    .clock(sram_2_clock),
    .io_en(sram_2_io_en),
    .io_wen(sram_2_io_wen),
    .io_addr(sram_2_io_addr),
    .io_wdata(sram_2_io_wdata),
    .io_rdata(sram_2_io_rdata)
  );
  ysyx_210128_Sram sram_3 ( // @[Cache.scala 89:22]
    .clock(sram_3_clock),
    .io_en(sram_3_io_en),
    .io_wen(sram_3_io_wen),
    .io_addr(sram_3_io_addr),
    .io_wdata(sram_3_io_wdata),
    .io_rdata(sram_3_io_rdata)
  );
  ysyx_210128_Meta meta_0 ( // @[Cache.scala 97:22]
    .clock(meta_0_clock),
    .reset(meta_0_reset),
    .io_idx(meta_0_io_idx),
    .io_tag_r(meta_0_io_tag_r),
    .io_tag_w(meta_0_io_tag_w),
    .io_tag_wen(meta_0_io_tag_wen),
    .io_dirty_r_async(meta_0_io_dirty_r_async),
    .io_dirty_w(meta_0_io_dirty_w),
    .io_dirty_wen(meta_0_io_dirty_wen),
    .io_valid_r_async(meta_0_io_valid_r_async),
    .io_invalidate(meta_0_io_invalidate)
  );
  ysyx_210128_Meta meta_1 ( // @[Cache.scala 97:22]
    .clock(meta_1_clock),
    .reset(meta_1_reset),
    .io_idx(meta_1_io_idx),
    .io_tag_r(meta_1_io_tag_r),
    .io_tag_w(meta_1_io_tag_w),
    .io_tag_wen(meta_1_io_tag_wen),
    .io_dirty_r_async(meta_1_io_dirty_r_async),
    .io_dirty_w(meta_1_io_dirty_w),
    .io_dirty_wen(meta_1_io_dirty_wen),
    .io_valid_r_async(meta_1_io_valid_r_async),
    .io_invalidate(meta_1_io_invalidate)
  );
  ysyx_210128_Meta meta_2 ( // @[Cache.scala 97:22]
    .clock(meta_2_clock),
    .reset(meta_2_reset),
    .io_idx(meta_2_io_idx),
    .io_tag_r(meta_2_io_tag_r),
    .io_tag_w(meta_2_io_tag_w),
    .io_tag_wen(meta_2_io_tag_wen),
    .io_dirty_r_async(meta_2_io_dirty_r_async),
    .io_dirty_w(meta_2_io_dirty_w),
    .io_dirty_wen(meta_2_io_dirty_wen),
    .io_valid_r_async(meta_2_io_valid_r_async),
    .io_invalidate(meta_2_io_invalidate)
  );
  ysyx_210128_Meta meta_3 ( // @[Cache.scala 97:22]
    .clock(meta_3_clock),
    .reset(meta_3_reset),
    .io_idx(meta_3_io_idx),
    .io_tag_r(meta_3_io_tag_r),
    .io_tag_w(meta_3_io_tag_w),
    .io_tag_wen(meta_3_io_tag_wen),
    .io_dirty_r_async(meta_3_io_dirty_r_async),
    .io_dirty_w(meta_3_io_dirty_w),
    .io_dirty_wen(meta_3_io_dirty_wen),
    .io_valid_r_async(meta_3_io_valid_r_async),
    .io_invalidate(meta_3_io_invalidate)
  );
  assign io_in_req_ready = pipeline_ready & ~fi_valid; // @[Cache.scala 287:34]
  assign io_in_resp_valid = s2_hit_real & state != 4'h8 | _T_18; // @[Cache.scala 288:71]
  assign io_in_resp_bits_rdata = 4'h0 == state ? _GEN_230 : _GEN_3297; // @[Cache.scala 318:18]
  assign io_in_resp_bits_user = s2_user; // @[Cache.scala 292:33]
  assign io_out_req_valid = _T_612 | _T_613; // @[Cache.scala 541:46]
  assign io_out_req_bits_addr = _T_611 ? _T_625 : _GEN_3536; // @[Cache.scala 550:34 553:23]
  assign io_out_req_bits_aen = _T_610 | _T_611; // @[Cache.scala 558:48]
  assign io_out_req_bits_wdata = _T_613 ? s2_reg_dat_w[127:64] : _GEN_3539; // @[Cache.scala 565:34 566:24]
  assign io_out_req_bits_wlast = state == 4'h5; // @[Cache.scala 575:32]
  assign io_out_req_bits_wen = _T_611 | _T_613; // @[Cache.scala 577:49]
  assign io_out_resp_ready = state == 4'h2 | _T_653; // @[Cache.scala 583:47]
  assign sram_0_clock = clock;
  assign sram_0_io_en = 4'h0 == state ? pipeline_ready : _GEN_3080; // @[Cache.scala 318:18]
  assign sram_0_io_wen = 4'h0 == state ? 1'h0 : _GEN_3081; // @[Cache.scala 318:18]
  assign sram_0_io_addr = 4'h0 == state ? _GEN_3 : _GEN_3082; // @[Cache.scala 318:18]
  assign sram_0_io_wdata = 4'h0 == state ? 128'h0 : _GEN_3083; // @[Cache.scala 318:18]
  assign sram_1_clock = clock;
  assign sram_1_io_en = 4'h0 == state ? pipeline_ready : _GEN_3086; // @[Cache.scala 318:18]
  assign sram_1_io_wen = 4'h0 == state ? 1'h0 : _GEN_3087; // @[Cache.scala 318:18]
  assign sram_1_io_addr = 4'h0 == state ? _GEN_3 : _GEN_3088; // @[Cache.scala 318:18]
  assign sram_1_io_wdata = 4'h0 == state ? 128'h0 : _GEN_3089; // @[Cache.scala 318:18]
  assign sram_2_clock = clock;
  assign sram_2_io_en = 4'h0 == state ? pipeline_ready : _GEN_3092; // @[Cache.scala 318:18]
  assign sram_2_io_wen = 4'h0 == state ? 1'h0 : _GEN_3093; // @[Cache.scala 318:18]
  assign sram_2_io_addr = 4'h0 == state ? _GEN_3 : _GEN_3094; // @[Cache.scala 318:18]
  assign sram_2_io_wdata = 4'h0 == state ? 128'h0 : _GEN_3095; // @[Cache.scala 318:18]
  assign sram_3_clock = clock;
  assign sram_3_io_en = 4'h0 == state ? pipeline_ready : _GEN_3098; // @[Cache.scala 318:18]
  assign sram_3_io_wen = 4'h0 == state ? 1'h0 : _GEN_3099; // @[Cache.scala 318:18]
  assign sram_3_io_addr = 4'h0 == state ? _GEN_3 : _GEN_3100; // @[Cache.scala 318:18]
  assign sram_3_io_wdata = 4'h0 == state ? 128'h0 : _GEN_3101; // @[Cache.scala 318:18]
  assign meta_0_clock = clock;
  assign meta_0_reset = reset;
  assign meta_0_io_idx = 4'h0 == state ? _GEN_3 : _GEN_3082; // @[Cache.scala 318:18]
  assign meta_0_io_tag_w = 4'h0 == state ? 21'h0 : _GEN_3084; // @[Cache.scala 114:16 318:18]
  assign meta_0_io_tag_wen = 4'h0 == state ? 1'h0 : _GEN_3081; // @[Cache.scala 115:18 318:18]
  assign meta_0_io_dirty_w = 1'h0; // @[Cache.scala 318:18]
  assign meta_0_io_dirty_wen = 4'h0 == state ? 1'h0 : _GEN_3081; // @[Cache.scala 318:18]
  assign meta_0_io_invalidate = fi_valid & fi_ready; // @[Cache.scala 164:26]
  assign meta_1_clock = clock;
  assign meta_1_reset = reset;
  assign meta_1_io_idx = 4'h0 == state ? _GEN_3 : _GEN_3088; // @[Cache.scala 318:18]
  assign meta_1_io_tag_w = 4'h0 == state ? 21'h0 : _GEN_3090; // @[Cache.scala 114:16 318:18]
  assign meta_1_io_tag_wen = 4'h0 == state ? 1'h0 : _GEN_3087; // @[Cache.scala 115:18 318:18]
  assign meta_1_io_dirty_w = 1'h0; // @[Cache.scala 318:18]
  assign meta_1_io_dirty_wen = 4'h0 == state ? 1'h0 : _GEN_3087; // @[Cache.scala 318:18]
  assign meta_1_io_invalidate = fi_valid & fi_ready; // @[Cache.scala 164:26]
  assign meta_2_clock = clock;
  assign meta_2_reset = reset;
  assign meta_2_io_idx = 4'h0 == state ? _GEN_3 : _GEN_3094; // @[Cache.scala 318:18]
  assign meta_2_io_tag_w = 4'h0 == state ? 21'h0 : _GEN_3096; // @[Cache.scala 114:16 318:18]
  assign meta_2_io_tag_wen = 4'h0 == state ? 1'h0 : _GEN_3093; // @[Cache.scala 115:18 318:18]
  assign meta_2_io_dirty_w = 1'h0; // @[Cache.scala 318:18]
  assign meta_2_io_dirty_wen = 4'h0 == state ? 1'h0 : _GEN_3093; // @[Cache.scala 318:18]
  assign meta_2_io_invalidate = fi_valid & fi_ready; // @[Cache.scala 164:26]
  assign meta_3_clock = clock;
  assign meta_3_reset = reset;
  assign meta_3_io_idx = 4'h0 == state ? _GEN_3 : _GEN_3100; // @[Cache.scala 318:18]
  assign meta_3_io_tag_w = 4'h0 == state ? 21'h0 : _GEN_3102; // @[Cache.scala 114:16 318:18]
  assign meta_3_io_tag_wen = 4'h0 == state ? 1'h0 : _GEN_3099; // @[Cache.scala 115:18 318:18]
  assign meta_3_io_dirty_w = 1'h0; // @[Cache.scala 318:18]
  assign meta_3_io_dirty_wen = 4'h0 == state ? 1'h0 : _GEN_3099; // @[Cache.scala 318:18]
  assign meta_3_io_invalidate = fi_valid & fi_ready; // @[Cache.scala 164:26]
  always @(posedge clock) begin
    REG <= meta_0_io_valid_r_async; // @[Cache.scala 123:59]
    REG_1 <= meta_1_io_valid_r_async; // @[Cache.scala 123:59]
    REG_2 <= meta_2_io_valid_r_async; // @[Cache.scala 123:59]
    REG_3 <= meta_3_io_valid_r_async; // @[Cache.scala 123:59]
    REG_4 <= meta_0_io_dirty_r_async; // @[Cache.scala 124:59]
    REG_5 <= meta_1_io_dirty_r_async; // @[Cache.scala 124:59]
    REG_6 <= meta_2_io_dirty_r_async; // @[Cache.scala 124:59]
    REG_7 <= meta_3_io_dirty_r_async; // @[Cache.scala 124:59]
    if (reset) begin // @[Cache.scala 129:22]
      plru0_0 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_0 <= _GEN_231;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_0 <= _GEN_2662;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_1 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_1 <= _GEN_232;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_1 <= _GEN_2663;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_2 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_2 <= _GEN_233;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_2 <= _GEN_2664;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_3 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_3 <= _GEN_234;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_3 <= _GEN_2665;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_4 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_4 <= _GEN_235;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_4 <= _GEN_2666;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_5 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_5 <= _GEN_236;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_5 <= _GEN_2667;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_6 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_6 <= _GEN_237;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_6 <= _GEN_2668;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_7 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_7 <= _GEN_238;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_7 <= _GEN_2669;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_8 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_8 <= _GEN_239;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_8 <= _GEN_2670;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_9 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_9 <= _GEN_240;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_9 <= _GEN_2671;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_10 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_10 <= _GEN_241;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_10 <= _GEN_2672;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_11 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_11 <= _GEN_242;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_11 <= _GEN_2673;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_12 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_12 <= _GEN_243;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_12 <= _GEN_2674;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_13 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_13 <= _GEN_244;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_13 <= _GEN_2675;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_14 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_14 <= _GEN_245;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_14 <= _GEN_2676;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_15 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_15 <= _GEN_246;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_15 <= _GEN_2677;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_16 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_16 <= _GEN_247;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_16 <= _GEN_2678;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_17 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_17 <= _GEN_248;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_17 <= _GEN_2679;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_18 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_18 <= _GEN_249;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_18 <= _GEN_2680;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_19 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_19 <= _GEN_250;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_19 <= _GEN_2681;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_20 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_20 <= _GEN_251;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_20 <= _GEN_2682;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_21 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_21 <= _GEN_252;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_21 <= _GEN_2683;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_22 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_22 <= _GEN_253;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_22 <= _GEN_2684;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_23 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_23 <= _GEN_254;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_23 <= _GEN_2685;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_24 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_24 <= _GEN_255;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_24 <= _GEN_2686;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_25 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_25 <= _GEN_256;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_25 <= _GEN_2687;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_26 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_26 <= _GEN_257;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_26 <= _GEN_2688;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_27 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_27 <= _GEN_258;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_27 <= _GEN_2689;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_28 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_28 <= _GEN_259;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_28 <= _GEN_2690;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_29 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_29 <= _GEN_260;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_29 <= _GEN_2691;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_30 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_30 <= _GEN_261;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_30 <= _GEN_2692;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_31 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_31 <= _GEN_262;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_31 <= _GEN_2693;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_32 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_32 <= _GEN_263;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_32 <= _GEN_2694;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_33 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_33 <= _GEN_264;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_33 <= _GEN_2695;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_34 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_34 <= _GEN_265;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_34 <= _GEN_2696;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_35 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_35 <= _GEN_266;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_35 <= _GEN_2697;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_36 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_36 <= _GEN_267;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_36 <= _GEN_2698;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_37 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_37 <= _GEN_268;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_37 <= _GEN_2699;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_38 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_38 <= _GEN_269;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_38 <= _GEN_2700;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_39 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_39 <= _GEN_270;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_39 <= _GEN_2701;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_40 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_40 <= _GEN_271;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_40 <= _GEN_2702;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_41 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_41 <= _GEN_272;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_41 <= _GEN_2703;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_42 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_42 <= _GEN_273;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_42 <= _GEN_2704;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_43 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_43 <= _GEN_274;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_43 <= _GEN_2705;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_44 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_44 <= _GEN_275;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_44 <= _GEN_2706;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_45 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_45 <= _GEN_276;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_45 <= _GEN_2707;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_46 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_46 <= _GEN_277;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_46 <= _GEN_2708;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_47 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_47 <= _GEN_278;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_47 <= _GEN_2709;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_48 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_48 <= _GEN_279;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_48 <= _GEN_2710;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_49 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_49 <= _GEN_280;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_49 <= _GEN_2711;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_50 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_50 <= _GEN_281;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_50 <= _GEN_2712;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_51 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_51 <= _GEN_282;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_51 <= _GEN_2713;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_52 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_52 <= _GEN_283;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_52 <= _GEN_2714;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_53 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_53 <= _GEN_284;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_53 <= _GEN_2715;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_54 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_54 <= _GEN_285;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_54 <= _GEN_2716;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_55 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_55 <= _GEN_286;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_55 <= _GEN_2717;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_56 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_56 <= _GEN_287;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_56 <= _GEN_2718;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_57 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_57 <= _GEN_288;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_57 <= _GEN_2719;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_58 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_58 <= _GEN_289;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_58 <= _GEN_2720;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_59 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_59 <= _GEN_290;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_59 <= _GEN_2721;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_60 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_60 <= _GEN_291;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_60 <= _GEN_2722;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_61 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_61 <= _GEN_292;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_61 <= _GEN_2723;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_62 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_62 <= _GEN_293;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_62 <= _GEN_2724;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_63 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_63 <= _GEN_294;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_63 <= _GEN_2725;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_0 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_0 <= _GEN_423;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_0 <= _GEN_2726;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_1 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_1 <= _GEN_424;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_1 <= _GEN_2727;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_2 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_2 <= _GEN_425;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_2 <= _GEN_2728;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_3 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_3 <= _GEN_426;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_3 <= _GEN_2729;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_4 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_4 <= _GEN_427;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_4 <= _GEN_2730;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_5 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_5 <= _GEN_428;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_5 <= _GEN_2731;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_6 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_6 <= _GEN_429;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_6 <= _GEN_2732;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_7 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_7 <= _GEN_430;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_7 <= _GEN_2733;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_8 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_8 <= _GEN_431;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_8 <= _GEN_2734;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_9 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_9 <= _GEN_432;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_9 <= _GEN_2735;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_10 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_10 <= _GEN_433;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_10 <= _GEN_2736;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_11 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_11 <= _GEN_434;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_11 <= _GEN_2737;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_12 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_12 <= _GEN_435;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_12 <= _GEN_2738;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_13 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_13 <= _GEN_436;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_13 <= _GEN_2739;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_14 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_14 <= _GEN_437;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_14 <= _GEN_2740;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_15 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_15 <= _GEN_438;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_15 <= _GEN_2741;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_16 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_16 <= _GEN_439;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_16 <= _GEN_2742;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_17 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_17 <= _GEN_440;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_17 <= _GEN_2743;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_18 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_18 <= _GEN_441;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_18 <= _GEN_2744;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_19 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_19 <= _GEN_442;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_19 <= _GEN_2745;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_20 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_20 <= _GEN_443;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_20 <= _GEN_2746;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_21 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_21 <= _GEN_444;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_21 <= _GEN_2747;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_22 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_22 <= _GEN_445;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_22 <= _GEN_2748;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_23 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_23 <= _GEN_446;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_23 <= _GEN_2749;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_24 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_24 <= _GEN_447;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_24 <= _GEN_2750;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_25 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_25 <= _GEN_448;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_25 <= _GEN_2751;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_26 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_26 <= _GEN_449;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_26 <= _GEN_2752;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_27 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_27 <= _GEN_450;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_27 <= _GEN_2753;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_28 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_28 <= _GEN_451;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_28 <= _GEN_2754;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_29 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_29 <= _GEN_452;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_29 <= _GEN_2755;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_30 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_30 <= _GEN_453;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_30 <= _GEN_2756;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_31 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_31 <= _GEN_454;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_31 <= _GEN_2757;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_32 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_32 <= _GEN_455;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_32 <= _GEN_2758;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_33 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_33 <= _GEN_456;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_33 <= _GEN_2759;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_34 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_34 <= _GEN_457;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_34 <= _GEN_2760;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_35 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_35 <= _GEN_458;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_35 <= _GEN_2761;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_36 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_36 <= _GEN_459;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_36 <= _GEN_2762;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_37 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_37 <= _GEN_460;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_37 <= _GEN_2763;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_38 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_38 <= _GEN_461;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_38 <= _GEN_2764;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_39 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_39 <= _GEN_462;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_39 <= _GEN_2765;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_40 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_40 <= _GEN_463;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_40 <= _GEN_2766;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_41 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_41 <= _GEN_464;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_41 <= _GEN_2767;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_42 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_42 <= _GEN_465;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_42 <= _GEN_2768;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_43 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_43 <= _GEN_466;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_43 <= _GEN_2769;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_44 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_44 <= _GEN_467;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_44 <= _GEN_2770;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_45 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_45 <= _GEN_468;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_45 <= _GEN_2771;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_46 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_46 <= _GEN_469;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_46 <= _GEN_2772;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_47 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_47 <= _GEN_470;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_47 <= _GEN_2773;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_48 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_48 <= _GEN_471;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_48 <= _GEN_2774;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_49 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_49 <= _GEN_472;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_49 <= _GEN_2775;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_50 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_50 <= _GEN_473;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_50 <= _GEN_2776;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_51 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_51 <= _GEN_474;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_51 <= _GEN_2777;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_52 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_52 <= _GEN_475;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_52 <= _GEN_2778;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_53 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_53 <= _GEN_476;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_53 <= _GEN_2779;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_54 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_54 <= _GEN_477;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_54 <= _GEN_2780;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_55 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_55 <= _GEN_478;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_55 <= _GEN_2781;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_56 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_56 <= _GEN_479;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_56 <= _GEN_2782;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_57 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_57 <= _GEN_480;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_57 <= _GEN_2783;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_58 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_58 <= _GEN_481;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_58 <= _GEN_2784;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_59 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_59 <= _GEN_482;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_59 <= _GEN_2785;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_60 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_60 <= _GEN_483;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_60 <= _GEN_2786;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_61 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_61 <= _GEN_484;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_61 <= _GEN_2787;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_62 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_62 <= _GEN_485;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_62 <= _GEN_2788;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_63 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_63 <= _GEN_486;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_63 <= _GEN_2789;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_0 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_0 <= _GEN_487;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_0 <= _GEN_2790;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_1 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_1 <= _GEN_488;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_1 <= _GEN_2791;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_2 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_2 <= _GEN_489;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_2 <= _GEN_2792;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_3 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_3 <= _GEN_490;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_3 <= _GEN_2793;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_4 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_4 <= _GEN_491;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_4 <= _GEN_2794;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_5 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_5 <= _GEN_492;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_5 <= _GEN_2795;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_6 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_6 <= _GEN_493;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_6 <= _GEN_2796;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_7 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_7 <= _GEN_494;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_7 <= _GEN_2797;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_8 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_8 <= _GEN_495;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_8 <= _GEN_2798;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_9 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_9 <= _GEN_496;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_9 <= _GEN_2799;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_10 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_10 <= _GEN_497;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_10 <= _GEN_2800;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_11 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_11 <= _GEN_498;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_11 <= _GEN_2801;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_12 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_12 <= _GEN_499;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_12 <= _GEN_2802;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_13 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_13 <= _GEN_500;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_13 <= _GEN_2803;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_14 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_14 <= _GEN_501;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_14 <= _GEN_2804;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_15 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_15 <= _GEN_502;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_15 <= _GEN_2805;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_16 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_16 <= _GEN_503;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_16 <= _GEN_2806;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_17 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_17 <= _GEN_504;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_17 <= _GEN_2807;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_18 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_18 <= _GEN_505;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_18 <= _GEN_2808;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_19 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_19 <= _GEN_506;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_19 <= _GEN_2809;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_20 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_20 <= _GEN_507;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_20 <= _GEN_2810;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_21 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_21 <= _GEN_508;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_21 <= _GEN_2811;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_22 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_22 <= _GEN_509;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_22 <= _GEN_2812;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_23 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_23 <= _GEN_510;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_23 <= _GEN_2813;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_24 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_24 <= _GEN_511;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_24 <= _GEN_2814;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_25 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_25 <= _GEN_512;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_25 <= _GEN_2815;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_26 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_26 <= _GEN_513;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_26 <= _GEN_2816;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_27 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_27 <= _GEN_514;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_27 <= _GEN_2817;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_28 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_28 <= _GEN_515;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_28 <= _GEN_2818;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_29 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_29 <= _GEN_516;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_29 <= _GEN_2819;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_30 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_30 <= _GEN_517;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_30 <= _GEN_2820;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_31 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_31 <= _GEN_518;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_31 <= _GEN_2821;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_32 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_32 <= _GEN_519;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_32 <= _GEN_2822;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_33 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_33 <= _GEN_520;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_33 <= _GEN_2823;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_34 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_34 <= _GEN_521;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_34 <= _GEN_2824;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_35 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_35 <= _GEN_522;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_35 <= _GEN_2825;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_36 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_36 <= _GEN_523;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_36 <= _GEN_2826;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_37 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_37 <= _GEN_524;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_37 <= _GEN_2827;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_38 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_38 <= _GEN_525;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_38 <= _GEN_2828;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_39 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_39 <= _GEN_526;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_39 <= _GEN_2829;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_40 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_40 <= _GEN_527;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_40 <= _GEN_2830;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_41 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_41 <= _GEN_528;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_41 <= _GEN_2831;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_42 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_42 <= _GEN_529;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_42 <= _GEN_2832;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_43 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_43 <= _GEN_530;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_43 <= _GEN_2833;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_44 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_44 <= _GEN_531;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_44 <= _GEN_2834;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_45 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_45 <= _GEN_532;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_45 <= _GEN_2835;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_46 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_46 <= _GEN_533;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_46 <= _GEN_2836;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_47 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_47 <= _GEN_534;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_47 <= _GEN_2837;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_48 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_48 <= _GEN_535;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_48 <= _GEN_2838;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_49 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_49 <= _GEN_536;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_49 <= _GEN_2839;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_50 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_50 <= _GEN_537;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_50 <= _GEN_2840;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_51 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_51 <= _GEN_538;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_51 <= _GEN_2841;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_52 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_52 <= _GEN_539;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_52 <= _GEN_2842;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_53 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_53 <= _GEN_540;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_53 <= _GEN_2843;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_54 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_54 <= _GEN_541;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_54 <= _GEN_2844;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_55 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_55 <= _GEN_542;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_55 <= _GEN_2845;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_56 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_56 <= _GEN_543;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_56 <= _GEN_2846;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_57 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_57 <= _GEN_544;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_57 <= _GEN_2847;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_58 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_58 <= _GEN_545;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_58 <= _GEN_2848;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_59 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_59 <= _GEN_546;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_59 <= _GEN_2849;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_60 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_60 <= _GEN_547;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_60 <= _GEN_2850;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_61 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_61 <= _GEN_548;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_61 <= _GEN_2851;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_62 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_62 <= _GEN_549;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_62 <= _GEN_2852;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_63 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_63 <= _GEN_550;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_63 <= _GEN_2853;
      end
    end
    REG_9 <= (hit_ready | _T_18) & io_in_resp_ready | invalid_ready; // @[Cache.scala 282:66]
    if (reset) begin // @[Cache.scala 215:25]
      s2_addr <= 32'h0; // @[Cache.scala 215:25]
    end else if (pipeline_ready) begin // @[Cache.scala 246:24]
      s2_addr <= io_in_req_bits_addr; // @[Cache.scala 248:14]
    end
    if (reset) begin // @[Cache.scala 239:27]
      s2_reg_hit <= 1'h0; // @[Cache.scala 239:27]
    end else if (!(pipeline_ready)) begin // @[Cache.scala 246:24]
      if (~pipeline_ready & REG_8) begin // @[Cache.scala 256:58]
        s2_reg_hit <= s2_hit; // @[Cache.scala 259:18]
      end
    end
    if (reset) begin // @[Cache.scala 213:22]
      state <= 4'h8; // @[Cache.scala 213:22]
    end else if (fi_fire) begin // @[Cache.scala 447:18]
      state <= 4'h8; // @[Cache.scala 448:11]
    end else if (pipeline_ready) begin // @[Cache.scala 417:24]
      if (io_in_req_valid) begin // @[Cache.scala 418:17]
        state <= 4'h0;
      end else begin
        state <= 4'h8;
      end
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      state <= _GEN_985;
    end else begin
      state <= _GEN_3077;
    end
    if (reset) begin // @[Utils.scala 34:20]
      fi_valid <= 1'h0; // @[Utils.scala 34:20]
    end else if (dcache_fi_complete) begin // @[Utils.scala 41:19]
      fi_valid <= 1'h0; // @[Utils.scala 41:23]
    end else begin
      fi_valid <= _GEN_0;
    end
    if (reset) begin // @[Cache.scala 222:25]
      s2_user <= 68'h0; // @[Cache.scala 222:25]
    end else if (pipeline_ready) begin // @[Cache.scala 246:24]
      s2_user <= io_in_req_bits_user; // @[Cache.scala 253:15]
    end
    if (reset) begin // @[Cache.scala 241:29]
      s2_reg_rdata <= 128'h0; // @[Cache.scala 241:29]
    end else if (!(pipeline_ready)) begin // @[Cache.scala 246:24]
      if (~pipeline_ready & REG_8) begin // @[Cache.scala 256:58]
        if (2'h3 == s2_way) begin // @[Cache.scala 261:18]
          s2_reg_rdata <= sram_out_3; // @[Cache.scala 261:18]
        end else begin
          s2_reg_rdata <= _GEN_6;
        end
      end
    end
    if (reset) begin // @[Cache.scala 242:29]
      s2_reg_dirty <= 1'h0; // @[Cache.scala 242:29]
    end else if (!(pipeline_ready)) begin // @[Cache.scala 246:24]
      if (~pipeline_ready & REG_8) begin // @[Cache.scala 256:58]
        if (2'h3 == replace_way) begin // @[Cache.scala 262:18]
          s2_reg_dirty <= REG_7; // @[Cache.scala 262:18]
        end else begin
          s2_reg_dirty <= _GEN_10;
        end
      end
    end
    if (reset) begin // @[Cache.scala 243:29]
      s2_reg_tag_r <= 21'h0; // @[Cache.scala 243:29]
    end else if (!(pipeline_ready)) begin // @[Cache.scala 246:24]
      if (~pipeline_ready & REG_8) begin // @[Cache.scala 256:58]
        if (2'h3 == replace_way) begin // @[Cache.scala 263:18]
          s2_reg_tag_r <= tag_out_3; // @[Cache.scala 263:18]
        end else begin
          s2_reg_tag_r <= _GEN_14;
        end
      end
    end
    if (reset) begin // @[Cache.scala 244:29]
      s2_reg_dat_w <= 128'h0; // @[Cache.scala 244:29]
    end else if (!(pipeline_ready)) begin // @[Cache.scala 246:24]
      if (~pipeline_ready & REG_8) begin // @[Cache.scala 256:58]
        if (2'h3 == replace_way) begin // @[Cache.scala 264:18]
          s2_reg_dat_w <= sram_out_3; // @[Cache.scala 264:18]
        end else begin
          s2_reg_dat_w <= _GEN_18;
        end
      end
    end
    REG_8 <= (hit_ready | _T_18) & io_in_resp_ready | invalid_ready; // @[Cache.scala 282:66]
    if (reset) begin // @[Cache.scala 270:23]
      wdata1 <= 64'h0; // @[Cache.scala 270:23]
    end else if (!(4'h0 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
        if (4'h2 == state) begin // @[Cache.scala 318:18]
          wdata1 <= _GEN_990;
        end
      end
    end
    if (reset) begin // @[Cache.scala 271:23]
      wdata2 <= 64'h0; // @[Cache.scala 271:23]
    end else if (!(4'h0 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
        if (4'h2 == state) begin // @[Cache.scala 318:18]
          wdata2 <= _GEN_991;
        end
      end
    end
    REG_10 <= (hit_ready | _T_18) & io_in_resp_ready | invalid_ready; // @[Cache.scala 282:66]
    REG_11 <= (hit_ready | _T_18) & io_in_resp_ready | invalid_ready; // @[Cache.scala 282:66]
    if (s2_offs) begin // @[Cache.scala 410:40]
      REG_12 <= wdata2;
    end else begin
      REG_12 <= wdata1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  REG_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  REG_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  REG_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  plru0_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  plru0_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  plru0_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  plru0_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  plru0_4 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  plru0_5 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  plru0_6 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  plru0_7 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  plru0_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  plru0_9 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  plru0_10 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  plru0_11 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  plru0_12 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  plru0_13 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  plru0_14 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  plru0_15 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  plru0_16 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  plru0_17 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  plru0_18 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  plru0_19 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  plru0_20 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  plru0_21 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  plru0_22 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  plru0_23 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  plru0_24 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  plru0_25 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  plru0_26 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  plru0_27 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  plru0_28 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  plru0_29 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  plru0_30 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  plru0_31 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  plru0_32 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  plru0_33 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  plru0_34 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  plru0_35 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  plru0_36 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  plru0_37 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  plru0_38 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  plru0_39 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  plru0_40 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  plru0_41 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  plru0_42 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  plru0_43 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  plru0_44 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  plru0_45 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  plru0_46 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  plru0_47 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  plru0_48 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  plru0_49 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  plru0_50 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  plru0_51 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  plru0_52 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  plru0_53 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  plru0_54 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  plru0_55 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  plru0_56 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  plru0_57 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  plru0_58 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  plru0_59 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  plru0_60 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  plru0_61 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  plru0_62 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  plru0_63 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  plru1_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  plru1_1 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  plru1_2 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  plru1_3 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  plru1_4 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  plru1_5 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  plru1_6 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  plru1_7 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  plru1_8 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  plru1_9 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  plru1_10 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  plru1_11 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  plru1_12 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  plru1_13 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  plru1_14 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  plru1_15 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  plru1_16 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  plru1_17 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  plru1_18 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  plru1_19 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  plru1_20 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  plru1_21 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  plru1_22 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  plru1_23 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  plru1_24 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  plru1_25 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  plru1_26 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  plru1_27 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  plru1_28 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  plru1_29 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  plru1_30 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  plru1_31 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  plru1_32 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  plru1_33 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  plru1_34 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  plru1_35 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  plru1_36 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  plru1_37 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  plru1_38 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  plru1_39 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  plru1_40 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  plru1_41 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  plru1_42 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  plru1_43 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  plru1_44 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  plru1_45 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  plru1_46 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  plru1_47 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  plru1_48 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  plru1_49 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  plru1_50 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  plru1_51 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  plru1_52 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  plru1_53 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  plru1_54 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  plru1_55 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  plru1_56 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  plru1_57 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  plru1_58 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  plru1_59 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  plru1_60 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  plru1_61 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  plru1_62 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  plru1_63 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  plru2_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  plru2_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  plru2_2 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  plru2_3 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  plru2_4 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  plru2_5 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  plru2_6 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  plru2_7 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  plru2_8 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  plru2_9 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  plru2_10 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  plru2_11 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  plru2_12 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  plru2_13 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  plru2_14 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  plru2_15 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  plru2_16 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  plru2_17 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  plru2_18 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  plru2_19 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  plru2_20 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  plru2_21 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  plru2_22 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  plru2_23 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  plru2_24 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  plru2_25 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  plru2_26 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  plru2_27 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  plru2_28 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  plru2_29 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  plru2_30 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  plru2_31 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  plru2_32 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  plru2_33 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  plru2_34 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  plru2_35 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  plru2_36 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  plru2_37 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  plru2_38 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  plru2_39 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  plru2_40 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  plru2_41 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  plru2_42 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  plru2_43 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  plru2_44 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  plru2_45 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  plru2_46 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  plru2_47 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  plru2_48 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  plru2_49 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  plru2_50 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  plru2_51 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  plru2_52 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  plru2_53 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  plru2_54 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  plru2_55 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  plru2_56 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  plru2_57 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  plru2_58 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  plru2_59 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  plru2_60 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  plru2_61 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  plru2_62 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  plru2_63 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  REG_9 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  s2_addr = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  s2_reg_hit = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  state = _RAND_203[3:0];
  _RAND_204 = {1{`RANDOM}};
  fi_valid = _RAND_204[0:0];
  _RAND_205 = {3{`RANDOM}};
  s2_user = _RAND_205[67:0];
  _RAND_206 = {4{`RANDOM}};
  s2_reg_rdata = _RAND_206[127:0];
  _RAND_207 = {1{`RANDOM}};
  s2_reg_dirty = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  s2_reg_tag_r = _RAND_208[20:0];
  _RAND_209 = {4{`RANDOM}};
  s2_reg_dat_w = _RAND_209[127:0];
  _RAND_210 = {1{`RANDOM}};
  REG_8 = _RAND_210[0:0];
  _RAND_211 = {2{`RANDOM}};
  wdata1 = _RAND_211[63:0];
  _RAND_212 = {2{`RANDOM}};
  wdata2 = _RAND_212[63:0];
  _RAND_213 = {1{`RANDOM}};
  REG_10 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  REG_11 = _RAND_214[0:0];
  _RAND_215 = {2{`RANDOM}};
  REG_12 = _RAND_215[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_Uncache(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [67:0] io_in_req_bits_user,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output [67:0] io_in_resp_bits_user,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [1:0]  io_out_req_bits_size,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [95:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Uncache.scala 17:22]
  reg [31:0] addr; // @[Uncache.scala 20:22]
  reg [1:0] size; // @[Uncache.scala 24:22]
  reg [67:0] in_user; // @[Uncache.scala 26:24]
  reg [31:0] rdata_1; // @[Uncache.scala 29:24]
  reg [31:0] rdata_2; // @[Uncache.scala 30:24]
  wire  req_split = size == 2'h3 & addr[2:0] == 3'h0; // @[Uncache.scala 34:35]
  wire  _T_5 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_10 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _T_14 = req_split ? 3'h3 : 3'h5; // @[Uncache.scala 68:21]
  wire [31:0] _GEN_11 = _T_12 ? io_out_resp_bits_rdata[31:0] : rdata_1; // @[Uncache.scala 66:30 67:17 29:24]
  wire [2:0] _GEN_12 = _T_12 ? _T_14 : state; // @[Uncache.scala 66:30 68:15 17:22]
  wire [2:0] _GEN_13 = _T_10 ? 3'h4 : state; // @[Uncache.scala 72:29 73:15 17:22]
  wire [31:0] _GEN_14 = _T_12 ? io_out_resp_bits_rdata[31:0] : rdata_2; // @[Uncache.scala 77:30 79:19 30:24]
  wire [2:0] _GEN_15 = _T_12 ? 3'h5 : state; // @[Uncache.scala 77:30 83:15 17:22]
  wire  _T_21 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_16 = _T_21 ? 3'h0 : state; // @[Uncache.scala 87:29 88:15 17:22]
  wire [2:0] _GEN_17 = 3'h5 == state ? _GEN_16 : state; // @[Uncache.scala 36:18 17:22]
  wire [31:0] _GEN_18 = 3'h4 == state ? _GEN_14 : rdata_2; // @[Uncache.scala 36:18 30:24]
  wire [2:0] _GEN_19 = 3'h4 == state ? _GEN_15 : _GEN_17; // @[Uncache.scala 36:18]
  wire [2:0] _GEN_20 = 3'h3 == state ? _GEN_13 : _GEN_19; // @[Uncache.scala 36:18]
  wire [31:0] _GEN_21 = 3'h3 == state ? rdata_2 : _GEN_18; // @[Uncache.scala 36:18 30:24]
  wire  _T_24 = state == 3'h3; // @[Uncache.scala 98:55]
  wire [31:0] _T_34 = addr + 32'h4; // @[Uncache.scala 115:70]
  assign io_in_req_ready = state == 3'h0; // @[Uncache.scala 97:34]
  assign io_in_resp_valid = state == 3'h5; // @[Uncache.scala 106:34]
  assign io_in_resp_bits_rdata = {rdata_2,rdata_1}; // @[Cat.scala 30:58]
  assign io_in_resp_bits_user = in_user; // @[Uncache.scala 111:33]
  assign io_out_req_valid = state == 3'h1 | state == 3'h3; // @[Uncache.scala 98:46]
  assign io_out_req_bits_addr = req_split & _T_24 ? _T_34 : addr; // @[Uncache.scala 115:30]
  assign io_out_req_bits_size = req_split ? 2'h2 : size; // @[Uncache.scala 118:30]
  assign io_out_resp_ready = state == 3'h2 | state == 3'h4; // @[Uncache.scala 105:47]
  always @(posedge clock) begin
    if (reset) begin // @[Uncache.scala 17:22]
      state <= 3'h0; // @[Uncache.scala 17:22]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        if (~io_in_req_bits_addr[2]) begin // @[Uncache.scala 52:21]
          state <= 3'h1;
        end else begin
          state <= 3'h3;
        end
      end
    end else if (3'h1 == state) begin // @[Uncache.scala 36:18]
      if (_T_10) begin // @[Uncache.scala 61:29]
        state <= 3'h2; // @[Uncache.scala 62:15]
      end
    end else if (3'h2 == state) begin // @[Uncache.scala 36:18]
      state <= _GEN_12;
    end else begin
      state <= _GEN_20;
    end
    if (reset) begin // @[Uncache.scala 20:22]
      addr <= 32'h0; // @[Uncache.scala 20:22]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        addr <= io_in_req_bits_addr; // @[Uncache.scala 39:15]
      end
    end
    if (reset) begin // @[Uncache.scala 24:22]
      size <= 2'h0; // @[Uncache.scala 24:22]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        size <= 2'h3; // @[Uncache.scala 43:15]
      end
    end
    if (reset) begin // @[Uncache.scala 26:24]
      in_user <= 68'h0; // @[Uncache.scala 26:24]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        in_user <= io_in_req_bits_user; // @[Uncache.scala 47:19]
      end
    end
    if (reset) begin // @[Uncache.scala 29:24]
      rdata_1 <= 32'h0; // @[Uncache.scala 29:24]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        rdata_1 <= 32'h0; // @[Uncache.scala 50:17]
      end
    end else if (!(3'h1 == state)) begin // @[Uncache.scala 36:18]
      if (3'h2 == state) begin // @[Uncache.scala 36:18]
        rdata_1 <= _GEN_11;
      end
    end
    if (reset) begin // @[Uncache.scala 30:24]
      rdata_2 <= 32'h0; // @[Uncache.scala 30:24]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        rdata_2 <= 32'h0; // @[Uncache.scala 51:17]
      end
    end else if (!(3'h1 == state)) begin // @[Uncache.scala 36:18]
      if (!(3'h2 == state)) begin // @[Uncache.scala 36:18]
        rdata_2 <= _GEN_21;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  size = _RAND_2[1:0];
  _RAND_3 = {3{`RANDOM}};
  in_user = _RAND_3[67:0];
  _RAND_4 = {1{`RANDOM}};
  rdata_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  rdata_2 = _RAND_5[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_CacheBusCrossbar1to2(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [67:0] io_in_req_bits_user,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output [67:0] io_in_resp_bits_user,
  input         io_out_0_req_ready,
  output        io_out_0_req_valid,
  output [31:0] io_out_0_req_bits_addr,
  output [67:0] io_out_0_req_bits_user,
  output        io_out_0_resp_ready,
  input         io_out_0_resp_valid,
  input  [63:0] io_out_0_resp_bits_rdata,
  input  [67:0] io_out_0_resp_bits_user,
  input         io_out_1_req_ready,
  output        io_out_1_req_valid,
  output [31:0] io_out_1_req_bits_addr,
  output [67:0] io_out_1_req_bits_user,
  output        io_out_1_resp_ready,
  input         io_out_1_resp_valid,
  input  [63:0] io_out_1_resp_bits_rdata,
  input  [67:0] io_out_1_resp_bits_user,
  input         io_to_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] in_flight_req_0; // @[Crossbar.scala 87:30]
  reg [7:0] in_flight_req_1; // @[Crossbar.scala 87:30]
  wire  _T = io_out_0_req_ready & io_out_0_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_1 = io_out_0_resp_ready & io_out_0_resp_valid; // @[Decoupled.scala 40:37]
  wire [7:0] _T_5 = in_flight_req_0 + 8'h1; // @[Crossbar.scala 90:44]
  wire [7:0] _T_11 = in_flight_req_0 - 8'h1; // @[Crossbar.scala 95:44]
  wire  _T_12 = io_out_1_req_ready & io_out_1_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_13 = io_out_1_resp_ready & io_out_1_resp_valid; // @[Decoupled.scala 40:37]
  wire [7:0] _T_17 = in_flight_req_1 + 8'h1; // @[Crossbar.scala 90:44]
  wire [7:0] _T_23 = in_flight_req_1 - 8'h1; // @[Crossbar.scala 95:44]
  wire  req_0_ready = in_flight_req_1 == 8'h0; // @[Crossbar.scala 102:39]
  wire  req_1_ready = in_flight_req_0 == 8'h0; // @[Crossbar.scala 103:39]
  reg  channel; // @[Crossbar.scala 105:24]
  wire  _GEN_4 = _T ? 1'h0 : channel; // @[Crossbar.scala 107:33 108:15 105:24]
  wire  _GEN_5 = _T_12 | _GEN_4; // @[Crossbar.scala 107:33 108:15]
  wire  _T_34 = ~channel; // @[Crossbar.scala 120:57]
  wire [67:0] _GEN_6 = _T_34 ? io_out_0_resp_bits_user : 68'h0; // @[Crossbar.scala 130:28 131:23 125:25]
  wire [63:0] _GEN_7 = _T_34 ? io_out_0_resp_bits_rdata : 64'h0; // @[Crossbar.scala 130:28 131:23 127:25]
  wire  _GEN_9 = _T_34 & io_out_0_resp_valid; // @[Crossbar.scala 130:28 132:24 128:25]
  assign io_in_req_ready = io_to_1 ? io_out_1_req_ready & req_1_ready : io_out_0_req_ready & req_0_ready; // @[Crossbar.scala 117:29]
  assign io_in_resp_valid = channel ? io_out_1_resp_valid : _GEN_9; // @[Crossbar.scala 130:28 132:24]
  assign io_in_resp_bits_rdata = channel ? io_out_1_resp_bits_rdata : _GEN_7; // @[Crossbar.scala 130:28 131:23]
  assign io_in_resp_bits_user = channel ? io_out_1_resp_bits_user : _GEN_6; // @[Crossbar.scala 130:28 131:23]
  assign io_out_0_req_valid = io_in_req_valid & ~io_to_1 & req_0_ready; // @[Crossbar.scala 115:54]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 113:23]
  assign io_out_0_req_bits_user = io_in_req_bits_user; // @[Crossbar.scala 113:23]
  assign io_out_0_resp_ready = io_in_resp_ready & ~channel; // @[Crossbar.scala 120:45]
  assign io_out_1_req_valid = io_in_req_valid & io_to_1 & req_1_ready; // @[Crossbar.scala 116:53]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 114:23]
  assign io_out_1_req_bits_user = io_in_req_bits_user; // @[Crossbar.scala 114:23]
  assign io_out_1_resp_ready = io_in_resp_ready & channel; // @[Crossbar.scala 121:45]
  always @(posedge clock) begin
    if (reset) begin // @[Crossbar.scala 87:30]
      in_flight_req_0 <= 8'h0; // @[Crossbar.scala 87:30]
    end else if (_T & ~_T_1) begin // @[Crossbar.scala 89:59]
      in_flight_req_0 <= _T_5; // @[Crossbar.scala 90:24]
    end else if (_T_1 & ~_T) begin // @[Crossbar.scala 94:66]
      in_flight_req_0 <= _T_11; // @[Crossbar.scala 95:24]
    end
    if (reset) begin // @[Crossbar.scala 87:30]
      in_flight_req_1 <= 8'h0; // @[Crossbar.scala 87:30]
    end else if (_T_12 & ~_T_13) begin // @[Crossbar.scala 89:59]
      in_flight_req_1 <= _T_17; // @[Crossbar.scala 90:24]
    end else if (_T_13 & ~_T_12) begin // @[Crossbar.scala 94:66]
      in_flight_req_1 <= _T_23; // @[Crossbar.scala 95:24]
    end
    if (reset) begin // @[Crossbar.scala 105:24]
      channel <= 1'h0; // @[Crossbar.scala 105:24]
    end else begin
      channel <= _GEN_5;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_req_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_req_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  channel = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_CacheController(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [67:0] io_in_req_bits_user,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output [67:0] io_in_resp_bits_user,
  input         io_out_cache_req_ready,
  output        io_out_cache_req_valid,
  output [31:0] io_out_cache_req_bits_addr,
  output        io_out_cache_req_bits_aen,
  output [63:0] io_out_cache_req_bits_wdata,
  output        io_out_cache_req_bits_wlast,
  output        io_out_cache_req_bits_wen,
  output        io_out_cache_resp_ready,
  input         io_out_cache_resp_valid,
  input  [63:0] io_out_cache_resp_bits_rdata,
  input         io_out_cache_resp_bits_rlast,
  input         io_out_uncache_req_ready,
  output        io_out_uncache_req_valid,
  output [31:0] io_out_uncache_req_bits_addr,
  output [1:0]  io_out_uncache_req_bits_size,
  output        io_out_uncache_resp_ready,
  input         io_out_uncache_resp_valid,
  input  [63:0] io_out_uncache_resp_bits_rdata,
  input         fence_i,
  input         _WIRE_10,
  input         empty
);
  wire  cache_clock; // @[CacheController.scala 14:21]
  wire  cache_reset; // @[CacheController.scala 14:21]
  wire  cache_io_in_req_ready; // @[CacheController.scala 14:21]
  wire  cache_io_in_req_valid; // @[CacheController.scala 14:21]
  wire [31:0] cache_io_in_req_bits_addr; // @[CacheController.scala 14:21]
  wire [67:0] cache_io_in_req_bits_user; // @[CacheController.scala 14:21]
  wire  cache_io_in_resp_ready; // @[CacheController.scala 14:21]
  wire  cache_io_in_resp_valid; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_in_resp_bits_rdata; // @[CacheController.scala 14:21]
  wire [67:0] cache_io_in_resp_bits_user; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_ready; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_valid; // @[CacheController.scala 14:21]
  wire [31:0] cache_io_out_req_bits_addr; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_bits_aen; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_out_req_bits_wdata; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_bits_wlast; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_bits_wen; // @[CacheController.scala 14:21]
  wire  cache_io_out_resp_ready; // @[CacheController.scala 14:21]
  wire  cache_io_out_resp_valid; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_out_resp_bits_rdata; // @[CacheController.scala 14:21]
  wire  cache_io_out_resp_bits_rlast; // @[CacheController.scala 14:21]
  wire  cache_fence_i_0; // @[CacheController.scala 14:21]
  wire  cache_dcache_fi_complete; // @[CacheController.scala 14:21]
  wire  cache_sq_empty_0; // @[CacheController.scala 14:21]
  wire  uncache_clock; // @[CacheController.scala 15:23]
  wire  uncache_reset; // @[CacheController.scala 15:23]
  wire  uncache_io_in_req_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_in_req_valid; // @[CacheController.scala 15:23]
  wire [31:0] uncache_io_in_req_bits_addr; // @[CacheController.scala 15:23]
  wire [67:0] uncache_io_in_req_bits_user; // @[CacheController.scala 15:23]
  wire  uncache_io_in_resp_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_in_resp_valid; // @[CacheController.scala 15:23]
  wire [63:0] uncache_io_in_resp_bits_rdata; // @[CacheController.scala 15:23]
  wire [67:0] uncache_io_in_resp_bits_user; // @[CacheController.scala 15:23]
  wire  uncache_io_out_req_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_out_req_valid; // @[CacheController.scala 15:23]
  wire [31:0] uncache_io_out_req_bits_addr; // @[CacheController.scala 15:23]
  wire [1:0] uncache_io_out_req_bits_size; // @[CacheController.scala 15:23]
  wire  uncache_io_out_resp_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_out_resp_valid; // @[CacheController.scala 15:23]
  wire [63:0] uncache_io_out_resp_bits_rdata; // @[CacheController.scala 15:23]
  wire  crossbar1to2_clock; // @[CacheController.scala 17:28]
  wire  crossbar1to2_reset; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_req_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_req_valid; // @[CacheController.scala 17:28]
  wire [31:0] crossbar1to2_io_in_req_bits_addr; // @[CacheController.scala 17:28]
  wire [67:0] crossbar1to2_io_in_req_bits_user; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_resp_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_resp_valid; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_in_resp_bits_rdata; // @[CacheController.scala 17:28]
  wire [67:0] crossbar1to2_io_in_resp_bits_user; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_req_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_req_valid; // @[CacheController.scala 17:28]
  wire [31:0] crossbar1to2_io_out_0_req_bits_addr; // @[CacheController.scala 17:28]
  wire [67:0] crossbar1to2_io_out_0_req_bits_user; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_resp_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_resp_valid; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_out_0_resp_bits_rdata; // @[CacheController.scala 17:28]
  wire [67:0] crossbar1to2_io_out_0_resp_bits_user; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_req_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_req_valid; // @[CacheController.scala 17:28]
  wire [31:0] crossbar1to2_io_out_1_req_bits_addr; // @[CacheController.scala 17:28]
  wire [67:0] crossbar1to2_io_out_1_req_bits_user; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_resp_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_resp_valid; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_out_1_resp_bits_rdata; // @[CacheController.scala 17:28]
  wire [67:0] crossbar1to2_io_out_1_resp_bits_user; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_to_1; // @[CacheController.scala 17:28]
  ysyx_210128_Cache cache ( // @[CacheController.scala 14:21]
    .clock(cache_clock),
    .reset(cache_reset),
    .io_in_req_ready(cache_io_in_req_ready),
    .io_in_req_valid(cache_io_in_req_valid),
    .io_in_req_bits_addr(cache_io_in_req_bits_addr),
    .io_in_req_bits_user(cache_io_in_req_bits_user),
    .io_in_resp_ready(cache_io_in_resp_ready),
    .io_in_resp_valid(cache_io_in_resp_valid),
    .io_in_resp_bits_rdata(cache_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(cache_io_in_resp_bits_user),
    .io_out_req_ready(cache_io_out_req_ready),
    .io_out_req_valid(cache_io_out_req_valid),
    .io_out_req_bits_addr(cache_io_out_req_bits_addr),
    .io_out_req_bits_aen(cache_io_out_req_bits_aen),
    .io_out_req_bits_wdata(cache_io_out_req_bits_wdata),
    .io_out_req_bits_wlast(cache_io_out_req_bits_wlast),
    .io_out_req_bits_wen(cache_io_out_req_bits_wen),
    .io_out_resp_ready(cache_io_out_resp_ready),
    .io_out_resp_valid(cache_io_out_resp_valid),
    .io_out_resp_bits_rdata(cache_io_out_resp_bits_rdata),
    .io_out_resp_bits_rlast(cache_io_out_resp_bits_rlast),
    .fence_i_0(cache_fence_i_0),
    .dcache_fi_complete(cache_dcache_fi_complete),
    .sq_empty_0(cache_sq_empty_0)
  );
  ysyx_210128_Uncache uncache ( // @[CacheController.scala 15:23]
    .clock(uncache_clock),
    .reset(uncache_reset),
    .io_in_req_ready(uncache_io_in_req_ready),
    .io_in_req_valid(uncache_io_in_req_valid),
    .io_in_req_bits_addr(uncache_io_in_req_bits_addr),
    .io_in_req_bits_user(uncache_io_in_req_bits_user),
    .io_in_resp_ready(uncache_io_in_resp_ready),
    .io_in_resp_valid(uncache_io_in_resp_valid),
    .io_in_resp_bits_rdata(uncache_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(uncache_io_in_resp_bits_user),
    .io_out_req_ready(uncache_io_out_req_ready),
    .io_out_req_valid(uncache_io_out_req_valid),
    .io_out_req_bits_addr(uncache_io_out_req_bits_addr),
    .io_out_req_bits_size(uncache_io_out_req_bits_size),
    .io_out_resp_ready(uncache_io_out_resp_ready),
    .io_out_resp_valid(uncache_io_out_resp_valid),
    .io_out_resp_bits_rdata(uncache_io_out_resp_bits_rdata)
  );
  ysyx_210128_CacheBusCrossbar1to2 crossbar1to2 ( // @[CacheController.scala 17:28]
    .clock(crossbar1to2_clock),
    .reset(crossbar1to2_reset),
    .io_in_req_ready(crossbar1to2_io_in_req_ready),
    .io_in_req_valid(crossbar1to2_io_in_req_valid),
    .io_in_req_bits_addr(crossbar1to2_io_in_req_bits_addr),
    .io_in_req_bits_user(crossbar1to2_io_in_req_bits_user),
    .io_in_resp_ready(crossbar1to2_io_in_resp_ready),
    .io_in_resp_valid(crossbar1to2_io_in_resp_valid),
    .io_in_resp_bits_rdata(crossbar1to2_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(crossbar1to2_io_in_resp_bits_user),
    .io_out_0_req_ready(crossbar1to2_io_out_0_req_ready),
    .io_out_0_req_valid(crossbar1to2_io_out_0_req_valid),
    .io_out_0_req_bits_addr(crossbar1to2_io_out_0_req_bits_addr),
    .io_out_0_req_bits_user(crossbar1to2_io_out_0_req_bits_user),
    .io_out_0_resp_ready(crossbar1to2_io_out_0_resp_ready),
    .io_out_0_resp_valid(crossbar1to2_io_out_0_resp_valid),
    .io_out_0_resp_bits_rdata(crossbar1to2_io_out_0_resp_bits_rdata),
    .io_out_0_resp_bits_user(crossbar1to2_io_out_0_resp_bits_user),
    .io_out_1_req_ready(crossbar1to2_io_out_1_req_ready),
    .io_out_1_req_valid(crossbar1to2_io_out_1_req_valid),
    .io_out_1_req_bits_addr(crossbar1to2_io_out_1_req_bits_addr),
    .io_out_1_req_bits_user(crossbar1to2_io_out_1_req_bits_user),
    .io_out_1_resp_ready(crossbar1to2_io_out_1_resp_ready),
    .io_out_1_resp_valid(crossbar1to2_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(crossbar1to2_io_out_1_resp_bits_rdata),
    .io_out_1_resp_bits_user(crossbar1to2_io_out_1_resp_bits_user),
    .io_to_1(crossbar1to2_io_to_1)
  );
  assign io_in_req_ready = crossbar1to2_io_in_req_ready; // @[CacheController.scala 19:22]
  assign io_in_resp_valid = crossbar1to2_io_in_resp_valid; // @[CacheController.scala 19:22]
  assign io_in_resp_bits_rdata = crossbar1to2_io_in_resp_bits_rdata; // @[CacheController.scala 19:22]
  assign io_in_resp_bits_user = crossbar1to2_io_in_resp_bits_user; // @[CacheController.scala 19:22]
  assign io_out_cache_req_valid = cache_io_out_req_valid; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_addr = cache_io_out_req_bits_addr; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_aen = cache_io_out_req_bits_aen; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_wdata = cache_io_out_req_bits_wdata; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_wlast = cache_io_out_req_bits_wlast; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_wen = cache_io_out_req_bits_wen; // @[CacheController.scala 23:16]
  assign io_out_cache_resp_ready = cache_io_out_resp_ready; // @[CacheController.scala 23:16]
  assign io_out_uncache_req_valid = uncache_io_out_req_valid; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_addr = uncache_io_out_req_bits_addr; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_size = uncache_io_out_req_bits_size; // @[CacheController.scala 24:18]
  assign io_out_uncache_resp_ready = uncache_io_out_resp_ready; // @[CacheController.scala 24:18]
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_io_in_req_valid = crossbar1to2_io_out_0_req_valid; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_addr = crossbar1to2_io_out_0_req_bits_addr; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_user = crossbar1to2_io_out_0_req_bits_user; // @[CacheController.scala 20:26]
  assign cache_io_in_resp_ready = crossbar1to2_io_out_0_resp_ready; // @[CacheController.scala 20:26]
  assign cache_io_out_req_ready = io_out_cache_req_ready; // @[CacheController.scala 23:16]
  assign cache_io_out_resp_valid = io_out_cache_resp_valid; // @[CacheController.scala 23:16]
  assign cache_io_out_resp_bits_rdata = io_out_cache_resp_bits_rdata; // @[CacheController.scala 23:16]
  assign cache_io_out_resp_bits_rlast = io_out_cache_resp_bits_rlast; // @[CacheController.scala 23:16]
  assign cache_fence_i_0 = fence_i;
  assign cache_dcache_fi_complete = _WIRE_10;
  assign cache_sq_empty_0 = empty;
  assign uncache_clock = clock;
  assign uncache_reset = reset;
  assign uncache_io_in_req_valid = crossbar1to2_io_out_1_req_valid; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_addr = crossbar1to2_io_out_1_req_bits_addr; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_user = crossbar1to2_io_out_1_req_bits_user; // @[CacheController.scala 21:26]
  assign uncache_io_in_resp_ready = crossbar1to2_io_out_1_resp_ready; // @[CacheController.scala 21:26]
  assign uncache_io_out_req_ready = io_out_uncache_req_ready; // @[CacheController.scala 24:18]
  assign uncache_io_out_resp_valid = io_out_uncache_resp_valid; // @[CacheController.scala 24:18]
  assign uncache_io_out_resp_bits_rdata = io_out_uncache_resp_bits_rdata; // @[CacheController.scala 24:18]
  assign crossbar1to2_clock = clock;
  assign crossbar1to2_reset = reset;
  assign crossbar1to2_io_in_req_valid = io_in_req_valid; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_addr = io_in_req_bits_addr; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_user = io_in_req_bits_user; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_resp_ready = io_in_resp_ready; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_out_0_req_ready = cache_io_in_req_ready; // @[CacheController.scala 20:26]
  assign crossbar1to2_io_out_0_resp_valid = cache_io_in_resp_valid; // @[CacheController.scala 20:26]
  assign crossbar1to2_io_out_0_resp_bits_rdata = cache_io_in_resp_bits_rdata; // @[CacheController.scala 20:26]
  assign crossbar1to2_io_out_0_resp_bits_user = cache_io_in_resp_bits_user; // @[CacheController.scala 20:26]
  assign crossbar1to2_io_out_1_req_ready = uncache_io_in_req_ready; // @[CacheController.scala 21:26]
  assign crossbar1to2_io_out_1_resp_valid = uncache_io_in_resp_valid; // @[CacheController.scala 21:26]
  assign crossbar1to2_io_out_1_resp_bits_rdata = uncache_io_in_resp_bits_rdata; // @[CacheController.scala 21:26]
  assign crossbar1to2_io_out_1_resp_bits_user = uncache_io_in_resp_bits_user; // @[CacheController.scala 21:26]
  assign crossbar1to2_io_to_1 = ~io_in_req_bits_addr[31]; // @[CacheController.scala 13:45]
endmodule
module ysyx_210128_InstBuffer(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_vec_0_pc,
  input  [31:0] io_in_bits_vec_0_inst,
  input         io_in_bits_vec_0_pred_br,
  input  [31:0] io_in_bits_vec_0_pred_bpc,
  input         io_in_bits_vec_0_valid,
  input  [31:0] io_in_bits_vec_1_pc,
  input  [31:0] io_in_bits_vec_1_inst,
  input         io_in_bits_vec_1_pred_br,
  input  [31:0] io_in_bits_vec_1_pred_bpc,
  input         io_in_bits_vec_1_valid,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_vec_0_pc,
  output [31:0] io_out_bits_vec_0_inst,
  output        io_out_bits_vec_0_pred_br,
  output [31:0] io_out_bits_vec_0_pred_bpc,
  output        io_out_bits_vec_0_valid,
  output [31:0] io_out_bits_vec_1_pc,
  output [31:0] io_out_bits_vec_1_inst,
  output        io_out_bits_vec_1_pred_br,
  output [31:0] io_out_bits_vec_1_pred_bpc,
  output        io_out_bits_vec_1_valid,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] buf_pc [0:7]; // @[InstBuffer.scala 48:24]
//   wire  buf_pc_MPORT_2_en; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pc_MPORT_2_addr; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pc_MPORT_2_data; // @[InstBuffer.scala 48:24]
//   wire  buf_pc_MPORT_3_en; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pc_MPORT_3_addr; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pc_MPORT_3_data; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pc_MPORT_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pc_MPORT_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pc_MPORT_1_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pc_MPORT_1_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_1_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_1_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pc_MPORT_4_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pc_MPORT_4_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_4_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_4_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pc_MPORT_5_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pc_MPORT_5_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_5_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_5_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pc_MPORT_6_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pc_MPORT_6_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_6_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_6_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pc_MPORT_7_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pc_MPORT_7_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_7_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_7_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pc_MPORT_8_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pc_MPORT_8_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_8_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_8_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pc_MPORT_9_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pc_MPORT_9_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_9_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_9_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pc_MPORT_10_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pc_MPORT_10_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_10_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_10_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pc_MPORT_11_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pc_MPORT_11_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_11_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pc_MPORT_11_en; // @[InstBuffer.scala 48:24]
//   reg  buf_pc_MPORT_2_en_pipe_0;
  reg [2:0] buf_pc_MPORT_2_addr_pipe_0;
//   reg  buf_pc_MPORT_3_en_pipe_0;
  reg [2:0] buf_pc_MPORT_3_addr_pipe_0;
  reg [31:0] buf_inst [0:7]; // @[InstBuffer.scala 48:24]
//   wire  buf_inst_MPORT_2_en; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_inst_MPORT_2_addr; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_inst_MPORT_2_data; // @[InstBuffer.scala 48:24]
//   wire  buf_inst_MPORT_3_en; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_inst_MPORT_3_addr; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_inst_MPORT_3_data; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_inst_MPORT_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_inst_MPORT_addr; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_mask; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_inst_MPORT_1_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_inst_MPORT_1_addr; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_1_mask; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_1_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_inst_MPORT_4_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_inst_MPORT_4_addr; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_4_mask; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_4_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_inst_MPORT_5_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_inst_MPORT_5_addr; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_5_mask; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_5_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_inst_MPORT_6_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_inst_MPORT_6_addr; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_6_mask; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_6_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_inst_MPORT_7_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_inst_MPORT_7_addr; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_7_mask; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_7_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_inst_MPORT_8_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_inst_MPORT_8_addr; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_8_mask; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_8_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_inst_MPORT_9_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_inst_MPORT_9_addr; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_9_mask; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_9_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_inst_MPORT_10_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_inst_MPORT_10_addr; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_10_mask; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_10_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_inst_MPORT_11_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_inst_MPORT_11_addr; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_11_mask; // @[InstBuffer.scala 48:24]
  wire  buf_inst_MPORT_11_en; // @[InstBuffer.scala 48:24]
//   reg  buf_inst_MPORT_2_en_pipe_0;
  reg [2:0] buf_inst_MPORT_2_addr_pipe_0;
//   reg  buf_inst_MPORT_3_en_pipe_0;
  reg [2:0] buf_inst_MPORT_3_addr_pipe_0;
  reg  buf_pred_br [0:7]; // @[InstBuffer.scala 48:24]
//   wire  buf_pred_br_MPORT_2_en; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_br_MPORT_2_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_2_data; // @[InstBuffer.scala 48:24]
//   wire  buf_pred_br_MPORT_3_en; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_br_MPORT_3_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_3_data; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_br_MPORT_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_en; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_1_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_br_MPORT_1_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_1_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_1_en; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_4_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_br_MPORT_4_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_4_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_4_en; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_5_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_br_MPORT_5_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_5_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_5_en; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_6_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_br_MPORT_6_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_6_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_6_en; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_7_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_br_MPORT_7_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_7_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_7_en; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_8_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_br_MPORT_8_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_8_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_8_en; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_9_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_br_MPORT_9_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_9_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_9_en; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_10_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_br_MPORT_10_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_10_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_10_en; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_11_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_br_MPORT_11_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_11_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_br_MPORT_11_en; // @[InstBuffer.scala 48:24]
//   reg  buf_pred_br_MPORT_2_en_pipe_0;
  reg [2:0] buf_pred_br_MPORT_2_addr_pipe_0;
//   reg  buf_pred_br_MPORT_3_en_pipe_0;
  reg [2:0] buf_pred_br_MPORT_3_addr_pipe_0;
  reg [31:0] buf_pred_bpc [0:7]; // @[InstBuffer.scala 48:24]
//   wire  buf_pred_bpc_MPORT_2_en; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_bpc_MPORT_2_addr; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pred_bpc_MPORT_2_data; // @[InstBuffer.scala 48:24]
//   wire  buf_pred_bpc_MPORT_3_en; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_bpc_MPORT_3_addr; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pred_bpc_MPORT_3_data; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pred_bpc_MPORT_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_bpc_MPORT_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pred_bpc_MPORT_1_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_bpc_MPORT_1_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_1_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_1_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pred_bpc_MPORT_4_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_bpc_MPORT_4_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_4_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_4_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pred_bpc_MPORT_5_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_bpc_MPORT_5_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_5_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_5_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pred_bpc_MPORT_6_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_bpc_MPORT_6_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_6_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_6_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pred_bpc_MPORT_7_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_bpc_MPORT_7_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_7_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_7_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pred_bpc_MPORT_8_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_bpc_MPORT_8_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_8_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_8_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pred_bpc_MPORT_9_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_bpc_MPORT_9_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_9_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_9_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pred_bpc_MPORT_10_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_bpc_MPORT_10_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_10_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_10_en; // @[InstBuffer.scala 48:24]
  wire [31:0] buf_pred_bpc_MPORT_11_data; // @[InstBuffer.scala 48:24]
  wire [2:0] buf_pred_bpc_MPORT_11_addr; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_11_mask; // @[InstBuffer.scala 48:24]
  wire  buf_pred_bpc_MPORT_11_en; // @[InstBuffer.scala 48:24]
//   reg  buf_pred_bpc_MPORT_2_en_pipe_0;
  reg [2:0] buf_pred_bpc_MPORT_2_addr_pipe_0;
//   reg  buf_pred_bpc_MPORT_3_en_pipe_0;
  reg [2:0] buf_pred_bpc_MPORT_3_addr_pipe_0;
  reg [3:0] enq_vec_0; // @[InstBuffer.scala 50:24]
  reg [3:0] enq_vec_1; // @[InstBuffer.scala 50:24]
  reg [3:0] deq_vec_0; // @[InstBuffer.scala 51:24]
  reg [3:0] deq_vec_1; // @[InstBuffer.scala 51:24]
  wire [2:0] enq_ptr = enq_vec_0[2:0]; // @[InstBuffer.scala 45:32]
  wire [2:0] deq_ptr = deq_vec_0[2:0]; // @[InstBuffer.scala 45:32]
  wire  enq_flag = enq_vec_0[3]; // @[InstBuffer.scala 46:33]
  wire  deq_flag = deq_vec_0[3]; // @[InstBuffer.scala 46:33]
  wire [2:0] _T_4 = enq_ptr - deq_ptr; // @[InstBuffer.scala 57:50]
  wire [3:0] _GEN_85 = {{1'd0}, enq_ptr}; // @[InstBuffer.scala 57:71]
  wire [3:0] _T_6 = 4'h8 + _GEN_85; // @[InstBuffer.scala 57:71]
  wire [3:0] _GEN_86 = {{1'd0}, deq_ptr}; // @[InstBuffer.scala 57:81]
  wire [3:0] _T_8 = _T_6 - _GEN_86; // @[InstBuffer.scala 57:81]
  wire [3:0] count = enq_flag == deq_flag ? {{1'd0}, _T_4} : _T_8; // @[InstBuffer.scala 57:18]
  reg  enq_ready; // @[InstBuffer.scala 58:26]
  wire  _T_9 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_10 = io_in_bits_vec_0_valid + io_in_bits_vec_1_valid; // @[Bitwise.scala 47:55]
  wire [1:0] num_enq = _T_9 ? _T_10 : 2'h0; // @[InstBuffer.scala 60:20]
  wire  _T_12 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_13 = io_out_bits_vec_0_valid + io_out_bits_vec_1_valid; // @[Bitwise.scala 47:55]
  wire [1:0] num_deq = _T_12 ? _T_13 : 2'h0; // @[InstBuffer.scala 61:20]
  wire  _T_15 = count >= 4'h2; // @[InstBuffer.scala 63:31]
  wire [3:0] num_try_deq = count >= 4'h2 ? 4'h2 : count; // @[InstBuffer.scala 63:24]
  wire [3:0] _GEN_87 = {{2'd0}, num_enq}; // @[InstBuffer.scala 64:29]
  wire [4:0] num_after_enq = count + _GEN_87; // @[InstBuffer.scala 64:29]
  wire [4:0] _GEN_88 = {{1'd0}, num_try_deq}; // @[InstBuffer.scala 65:58]
  wire [4:0] _T_17 = num_after_enq - _GEN_88; // @[InstBuffer.scala 65:58]
  wire [4:0] next_valid_entry = io_out_ready ? _T_17 : num_after_enq; // @[InstBuffer.scala 65:29]
  wire  _T_21 = io_in_bits_vec_0_valid & _T_9; // @[InstBuffer.scala 85:35]
  wire  _T_22 = ~io_flush; // @[InstBuffer.scala 85:54]
  wire  _T_26 = io_in_bits_vec_1_valid & _T_9; // @[InstBuffer.scala 85:35]
  wire [3:0] _GEN_12 = io_in_bits_vec_0_valid ? enq_vec_1 : enq_vec_0; // @[InstBuffer.scala 45:{32,32}]
  wire [3:0] next_enq_vec_0 = enq_vec_0 + _GEN_87; // @[InstBuffer.scala 92:44]
  wire [3:0] next_enq_vec_1 = enq_vec_1 + _GEN_87; // @[InstBuffer.scala 92:44]
  wire  shiftAmount = count[0]; // @[OneHot.scala 64:49]
  wire [1:0] _T_38 = 2'h1 << shiftAmount; // @[OneHot.scala 65:12]
  wire [1:0] _T_41 = _T_38 - 2'h1; // @[InstBuffer.scala 102:98]
  wire [1:0] valid_vec = _T_15 ? 2'h3 : _T_41; // @[InstBuffer.scala 102:22]
  wire [3:0] _GEN_91 = {{2'd0}, num_deq}; // @[InstBuffer.scala 103:44]
  wire [3:0] next_deq_vec_0 = deq_vec_0 + _GEN_91; // @[InstBuffer.scala 103:44]
  wire [3:0] next_deq_vec_1 = deq_vec_1 + _GEN_91; // @[InstBuffer.scala 103:44]
  wire [1:0] _T_54 = {io_out_bits_vec_0_valid,io_out_bits_vec_1_valid}; // @[Cat.scala 30:58]
  wire  _GEN_30 = io_flush | 5'h6 >= next_valid_entry; // @[InstBuffer.scala 116:19 117:15 67:13]
//   assign buf_pc_MPORT_2_en = buf_pc_MPORT_2_en_pipe_0;
  assign buf_pc_MPORT_2_addr = buf_pc_MPORT_2_addr_pipe_0;
  assign buf_pc_MPORT_2_data = buf_pc[buf_pc_MPORT_2_addr]; // @[InstBuffer.scala 48:24]
//   assign buf_pc_MPORT_3_en = buf_pc_MPORT_3_en_pipe_0;
  assign buf_pc_MPORT_3_addr = buf_pc_MPORT_3_addr_pipe_0;
  assign buf_pc_MPORT_3_data = buf_pc[buf_pc_MPORT_3_addr]; // @[InstBuffer.scala 48:24]
  assign buf_pc_MPORT_data = io_in_bits_vec_0_pc;
  assign buf_pc_MPORT_addr = enq_vec_0[2:0];
  assign buf_pc_MPORT_mask = 1'h1;
  assign buf_pc_MPORT_en = _T_21 & _T_22;
  assign buf_pc_MPORT_1_data = io_in_bits_vec_1_pc;
  assign buf_pc_MPORT_1_addr = _GEN_12[2:0];
  assign buf_pc_MPORT_1_mask = 1'h1;
  assign buf_pc_MPORT_1_en = _T_26 & _T_22;
  assign buf_pc_MPORT_4_data = 32'h0;
  assign buf_pc_MPORT_4_addr = 3'h0;
  assign buf_pc_MPORT_4_mask = 1'h1;
  assign buf_pc_MPORT_4_en = reset;
  assign buf_pc_MPORT_5_data = 32'h0;
  assign buf_pc_MPORT_5_addr = 3'h1;
  assign buf_pc_MPORT_5_mask = 1'h1;
  assign buf_pc_MPORT_5_en = reset;
  assign buf_pc_MPORT_6_data = 32'h0;
  assign buf_pc_MPORT_6_addr = 3'h2;
  assign buf_pc_MPORT_6_mask = 1'h1;
  assign buf_pc_MPORT_6_en = reset;
  assign buf_pc_MPORT_7_data = 32'h0;
  assign buf_pc_MPORT_7_addr = 3'h3;
  assign buf_pc_MPORT_7_mask = 1'h1;
  assign buf_pc_MPORT_7_en = reset;
  assign buf_pc_MPORT_8_data = 32'h0;
  assign buf_pc_MPORT_8_addr = 3'h4;
  assign buf_pc_MPORT_8_mask = 1'h1;
  assign buf_pc_MPORT_8_en = reset;
  assign buf_pc_MPORT_9_data = 32'h0;
  assign buf_pc_MPORT_9_addr = 3'h5;
  assign buf_pc_MPORT_9_mask = 1'h1;
  assign buf_pc_MPORT_9_en = reset;
  assign buf_pc_MPORT_10_data = 32'h0;
  assign buf_pc_MPORT_10_addr = 3'h6;
  assign buf_pc_MPORT_10_mask = 1'h1;
  assign buf_pc_MPORT_10_en = reset;
  assign buf_pc_MPORT_11_data = 32'h0;
  assign buf_pc_MPORT_11_addr = 3'h7;
  assign buf_pc_MPORT_11_mask = 1'h1;
  assign buf_pc_MPORT_11_en = reset;
//   assign buf_inst_MPORT_2_en = buf_inst_MPORT_2_en_pipe_0;
  assign buf_inst_MPORT_2_addr = buf_inst_MPORT_2_addr_pipe_0;
  assign buf_inst_MPORT_2_data = buf_inst[buf_inst_MPORT_2_addr]; // @[InstBuffer.scala 48:24]
//   assign buf_inst_MPORT_3_en = buf_inst_MPORT_3_en_pipe_0;
  assign buf_inst_MPORT_3_addr = buf_inst_MPORT_3_addr_pipe_0;
  assign buf_inst_MPORT_3_data = buf_inst[buf_inst_MPORT_3_addr]; // @[InstBuffer.scala 48:24]
  assign buf_inst_MPORT_data = io_in_bits_vec_0_inst;
  assign buf_inst_MPORT_addr = enq_vec_0[2:0];
  assign buf_inst_MPORT_mask = 1'h1;
  assign buf_inst_MPORT_en = _T_21 & _T_22;
  assign buf_inst_MPORT_1_data = io_in_bits_vec_1_inst;
  assign buf_inst_MPORT_1_addr = _GEN_12[2:0];
  assign buf_inst_MPORT_1_mask = 1'h1;
  assign buf_inst_MPORT_1_en = _T_26 & _T_22;
  assign buf_inst_MPORT_4_data = 32'h0;
  assign buf_inst_MPORT_4_addr = 3'h0;
  assign buf_inst_MPORT_4_mask = 1'h1;
  assign buf_inst_MPORT_4_en = reset;
  assign buf_inst_MPORT_5_data = 32'h0;
  assign buf_inst_MPORT_5_addr = 3'h1;
  assign buf_inst_MPORT_5_mask = 1'h1;
  assign buf_inst_MPORT_5_en = reset;
  assign buf_inst_MPORT_6_data = 32'h0;
  assign buf_inst_MPORT_6_addr = 3'h2;
  assign buf_inst_MPORT_6_mask = 1'h1;
  assign buf_inst_MPORT_6_en = reset;
  assign buf_inst_MPORT_7_data = 32'h0;
  assign buf_inst_MPORT_7_addr = 3'h3;
  assign buf_inst_MPORT_7_mask = 1'h1;
  assign buf_inst_MPORT_7_en = reset;
  assign buf_inst_MPORT_8_data = 32'h0;
  assign buf_inst_MPORT_8_addr = 3'h4;
  assign buf_inst_MPORT_8_mask = 1'h1;
  assign buf_inst_MPORT_8_en = reset;
  assign buf_inst_MPORT_9_data = 32'h0;
  assign buf_inst_MPORT_9_addr = 3'h5;
  assign buf_inst_MPORT_9_mask = 1'h1;
  assign buf_inst_MPORT_9_en = reset;
  assign buf_inst_MPORT_10_data = 32'h0;
  assign buf_inst_MPORT_10_addr = 3'h6;
  assign buf_inst_MPORT_10_mask = 1'h1;
  assign buf_inst_MPORT_10_en = reset;
  assign buf_inst_MPORT_11_data = 32'h0;
  assign buf_inst_MPORT_11_addr = 3'h7;
  assign buf_inst_MPORT_11_mask = 1'h1;
  assign buf_inst_MPORT_11_en = reset;
//   assign buf_pred_br_MPORT_2_en = buf_pred_br_MPORT_2_en_pipe_0;
  assign buf_pred_br_MPORT_2_addr = buf_pred_br_MPORT_2_addr_pipe_0;
  assign buf_pred_br_MPORT_2_data = buf_pred_br[buf_pred_br_MPORT_2_addr]; // @[InstBuffer.scala 48:24]
//   assign buf_pred_br_MPORT_3_en = buf_pred_br_MPORT_3_en_pipe_0;
  assign buf_pred_br_MPORT_3_addr = buf_pred_br_MPORT_3_addr_pipe_0;
  assign buf_pred_br_MPORT_3_data = buf_pred_br[buf_pred_br_MPORT_3_addr]; // @[InstBuffer.scala 48:24]
  assign buf_pred_br_MPORT_data = io_in_bits_vec_0_pred_br;
  assign buf_pred_br_MPORT_addr = enq_vec_0[2:0];
  assign buf_pred_br_MPORT_mask = 1'h1;
  assign buf_pred_br_MPORT_en = _T_21 & _T_22;
  assign buf_pred_br_MPORT_1_data = io_in_bits_vec_1_pred_br;
  assign buf_pred_br_MPORT_1_addr = _GEN_12[2:0];
  assign buf_pred_br_MPORT_1_mask = 1'h1;
  assign buf_pred_br_MPORT_1_en = _T_26 & _T_22;
  assign buf_pred_br_MPORT_4_data = 1'h0;
  assign buf_pred_br_MPORT_4_addr = 3'h0;
  assign buf_pred_br_MPORT_4_mask = 1'h1;
  assign buf_pred_br_MPORT_4_en = reset;
  assign buf_pred_br_MPORT_5_data = 1'h0;
  assign buf_pred_br_MPORT_5_addr = 3'h1;
  assign buf_pred_br_MPORT_5_mask = 1'h1;
  assign buf_pred_br_MPORT_5_en = reset;
  assign buf_pred_br_MPORT_6_data = 1'h0;
  assign buf_pred_br_MPORT_6_addr = 3'h2;
  assign buf_pred_br_MPORT_6_mask = 1'h1;
  assign buf_pred_br_MPORT_6_en = reset;
  assign buf_pred_br_MPORT_7_data = 1'h0;
  assign buf_pred_br_MPORT_7_addr = 3'h3;
  assign buf_pred_br_MPORT_7_mask = 1'h1;
  assign buf_pred_br_MPORT_7_en = reset;
  assign buf_pred_br_MPORT_8_data = 1'h0;
  assign buf_pred_br_MPORT_8_addr = 3'h4;
  assign buf_pred_br_MPORT_8_mask = 1'h1;
  assign buf_pred_br_MPORT_8_en = reset;
  assign buf_pred_br_MPORT_9_data = 1'h0;
  assign buf_pred_br_MPORT_9_addr = 3'h5;
  assign buf_pred_br_MPORT_9_mask = 1'h1;
  assign buf_pred_br_MPORT_9_en = reset;
  assign buf_pred_br_MPORT_10_data = 1'h0;
  assign buf_pred_br_MPORT_10_addr = 3'h6;
  assign buf_pred_br_MPORT_10_mask = 1'h1;
  assign buf_pred_br_MPORT_10_en = reset;
  assign buf_pred_br_MPORT_11_data = 1'h0;
  assign buf_pred_br_MPORT_11_addr = 3'h7;
  assign buf_pred_br_MPORT_11_mask = 1'h1;
  assign buf_pred_br_MPORT_11_en = reset;
//   assign buf_pred_bpc_MPORT_2_en = buf_pred_bpc_MPORT_2_en_pipe_0;
  assign buf_pred_bpc_MPORT_2_addr = buf_pred_bpc_MPORT_2_addr_pipe_0;
  assign buf_pred_bpc_MPORT_2_data = buf_pred_bpc[buf_pred_bpc_MPORT_2_addr]; // @[InstBuffer.scala 48:24]
//   assign buf_pred_bpc_MPORT_3_en = buf_pred_bpc_MPORT_3_en_pipe_0;
  assign buf_pred_bpc_MPORT_3_addr = buf_pred_bpc_MPORT_3_addr_pipe_0;
  assign buf_pred_bpc_MPORT_3_data = buf_pred_bpc[buf_pred_bpc_MPORT_3_addr]; // @[InstBuffer.scala 48:24]
  assign buf_pred_bpc_MPORT_data = io_in_bits_vec_0_pred_bpc;
  assign buf_pred_bpc_MPORT_addr = enq_vec_0[2:0];
  assign buf_pred_bpc_MPORT_mask = 1'h1;
  assign buf_pred_bpc_MPORT_en = _T_21 & _T_22;
  assign buf_pred_bpc_MPORT_1_data = io_in_bits_vec_1_pred_bpc;
  assign buf_pred_bpc_MPORT_1_addr = _GEN_12[2:0];
  assign buf_pred_bpc_MPORT_1_mask = 1'h1;
  assign buf_pred_bpc_MPORT_1_en = _T_26 & _T_22;
  assign buf_pred_bpc_MPORT_4_data = 32'h0;
  assign buf_pred_bpc_MPORT_4_addr = 3'h0;
  assign buf_pred_bpc_MPORT_4_mask = 1'h1;
  assign buf_pred_bpc_MPORT_4_en = reset;
  assign buf_pred_bpc_MPORT_5_data = 32'h0;
  assign buf_pred_bpc_MPORT_5_addr = 3'h1;
  assign buf_pred_bpc_MPORT_5_mask = 1'h1;
  assign buf_pred_bpc_MPORT_5_en = reset;
  assign buf_pred_bpc_MPORT_6_data = 32'h0;
  assign buf_pred_bpc_MPORT_6_addr = 3'h2;
  assign buf_pred_bpc_MPORT_6_mask = 1'h1;
  assign buf_pred_bpc_MPORT_6_en = reset;
  assign buf_pred_bpc_MPORT_7_data = 32'h0;
  assign buf_pred_bpc_MPORT_7_addr = 3'h3;
  assign buf_pred_bpc_MPORT_7_mask = 1'h1;
  assign buf_pred_bpc_MPORT_7_en = reset;
  assign buf_pred_bpc_MPORT_8_data = 32'h0;
  assign buf_pred_bpc_MPORT_8_addr = 3'h4;
  assign buf_pred_bpc_MPORT_8_mask = 1'h1;
  assign buf_pred_bpc_MPORT_8_en = reset;
  assign buf_pred_bpc_MPORT_9_data = 32'h0;
  assign buf_pred_bpc_MPORT_9_addr = 3'h5;
  assign buf_pred_bpc_MPORT_9_mask = 1'h1;
  assign buf_pred_bpc_MPORT_9_en = reset;
  assign buf_pred_bpc_MPORT_10_data = 32'h0;
  assign buf_pred_bpc_MPORT_10_addr = 3'h6;
  assign buf_pred_bpc_MPORT_10_mask = 1'h1;
  assign buf_pred_bpc_MPORT_10_en = reset;
  assign buf_pred_bpc_MPORT_11_data = 32'h0;
  assign buf_pred_bpc_MPORT_11_addr = 3'h7;
  assign buf_pred_bpc_MPORT_11_mask = 1'h1;
  assign buf_pred_bpc_MPORT_11_en = reset;
  assign io_in_ready = enq_ready; // @[InstBuffer.scala 98:15]
  assign io_out_valid = |_T_54; // @[InstBuffer.scala 112:53]
  assign io_out_bits_vec_0_pc = buf_pc_MPORT_2_data; // @[InstBuffer.scala 108:24]
  assign io_out_bits_vec_0_inst = buf_inst_MPORT_2_data; // @[InstBuffer.scala 108:24]
  assign io_out_bits_vec_0_pred_br = buf_pred_br_MPORT_2_data; // @[InstBuffer.scala 108:24]
  assign io_out_bits_vec_0_pred_bpc = buf_pred_bpc_MPORT_2_data; // @[InstBuffer.scala 108:24]
  assign io_out_bits_vec_0_valid = valid_vec[0]; // @[InstBuffer.scala 109:42]
  assign io_out_bits_vec_1_pc = buf_pc_MPORT_3_data; // @[InstBuffer.scala 108:24]
  assign io_out_bits_vec_1_inst = buf_inst_MPORT_3_data; // @[InstBuffer.scala 108:24]
  assign io_out_bits_vec_1_pred_br = buf_pred_br_MPORT_3_data; // @[InstBuffer.scala 108:24]
  assign io_out_bits_vec_1_pred_bpc = buf_pred_bpc_MPORT_3_data; // @[InstBuffer.scala 108:24]
  assign io_out_bits_vec_1_valid = valid_vec[1]; // @[InstBuffer.scala 109:42]
  always @(posedge clock) begin
    if (buf_pc_MPORT_en & buf_pc_MPORT_mask) begin
      buf_pc[buf_pc_MPORT_addr] <= buf_pc_MPORT_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pc_MPORT_1_en & buf_pc_MPORT_1_mask) begin
      buf_pc[buf_pc_MPORT_1_addr] <= buf_pc_MPORT_1_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pc_MPORT_4_en & buf_pc_MPORT_4_mask) begin
      buf_pc[buf_pc_MPORT_4_addr] <= buf_pc_MPORT_4_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pc_MPORT_5_en & buf_pc_MPORT_5_mask) begin
      buf_pc[buf_pc_MPORT_5_addr] <= buf_pc_MPORT_5_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pc_MPORT_6_en & buf_pc_MPORT_6_mask) begin
      buf_pc[buf_pc_MPORT_6_addr] <= buf_pc_MPORT_6_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pc_MPORT_7_en & buf_pc_MPORT_7_mask) begin
      buf_pc[buf_pc_MPORT_7_addr] <= buf_pc_MPORT_7_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pc_MPORT_8_en & buf_pc_MPORT_8_mask) begin
      buf_pc[buf_pc_MPORT_8_addr] <= buf_pc_MPORT_8_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pc_MPORT_9_en & buf_pc_MPORT_9_mask) begin
      buf_pc[buf_pc_MPORT_9_addr] <= buf_pc_MPORT_9_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pc_MPORT_10_en & buf_pc_MPORT_10_mask) begin
      buf_pc[buf_pc_MPORT_10_addr] <= buf_pc_MPORT_10_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pc_MPORT_11_en & buf_pc_MPORT_11_mask) begin
      buf_pc[buf_pc_MPORT_11_addr] <= buf_pc_MPORT_11_data; // @[InstBuffer.scala 48:24]
    end
//     buf_pc_MPORT_2_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      buf_pc_MPORT_2_addr_pipe_0 <= next_deq_vec_0[2:0];
    end
//     buf_pc_MPORT_3_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      buf_pc_MPORT_3_addr_pipe_0 <= next_deq_vec_1[2:0];
    end
    if (buf_inst_MPORT_en & buf_inst_MPORT_mask) begin
      buf_inst[buf_inst_MPORT_addr] <= buf_inst_MPORT_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_inst_MPORT_1_en & buf_inst_MPORT_1_mask) begin
      buf_inst[buf_inst_MPORT_1_addr] <= buf_inst_MPORT_1_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_inst_MPORT_4_en & buf_inst_MPORT_4_mask) begin
      buf_inst[buf_inst_MPORT_4_addr] <= buf_inst_MPORT_4_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_inst_MPORT_5_en & buf_inst_MPORT_5_mask) begin
      buf_inst[buf_inst_MPORT_5_addr] <= buf_inst_MPORT_5_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_inst_MPORT_6_en & buf_inst_MPORT_6_mask) begin
      buf_inst[buf_inst_MPORT_6_addr] <= buf_inst_MPORT_6_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_inst_MPORT_7_en & buf_inst_MPORT_7_mask) begin
      buf_inst[buf_inst_MPORT_7_addr] <= buf_inst_MPORT_7_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_inst_MPORT_8_en & buf_inst_MPORT_8_mask) begin
      buf_inst[buf_inst_MPORT_8_addr] <= buf_inst_MPORT_8_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_inst_MPORT_9_en & buf_inst_MPORT_9_mask) begin
      buf_inst[buf_inst_MPORT_9_addr] <= buf_inst_MPORT_9_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_inst_MPORT_10_en & buf_inst_MPORT_10_mask) begin
      buf_inst[buf_inst_MPORT_10_addr] <= buf_inst_MPORT_10_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_inst_MPORT_11_en & buf_inst_MPORT_11_mask) begin
      buf_inst[buf_inst_MPORT_11_addr] <= buf_inst_MPORT_11_data; // @[InstBuffer.scala 48:24]
    end
//     buf_inst_MPORT_2_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      buf_inst_MPORT_2_addr_pipe_0 <= next_deq_vec_0[2:0];
    end
//     buf_inst_MPORT_3_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      buf_inst_MPORT_3_addr_pipe_0 <= next_deq_vec_1[2:0];
    end
    if (buf_pred_br_MPORT_en & buf_pred_br_MPORT_mask) begin
      buf_pred_br[buf_pred_br_MPORT_addr] <= buf_pred_br_MPORT_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_br_MPORT_1_en & buf_pred_br_MPORT_1_mask) begin
      buf_pred_br[buf_pred_br_MPORT_1_addr] <= buf_pred_br_MPORT_1_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_br_MPORT_4_en & buf_pred_br_MPORT_4_mask) begin
      buf_pred_br[buf_pred_br_MPORT_4_addr] <= buf_pred_br_MPORT_4_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_br_MPORT_5_en & buf_pred_br_MPORT_5_mask) begin
      buf_pred_br[buf_pred_br_MPORT_5_addr] <= buf_pred_br_MPORT_5_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_br_MPORT_6_en & buf_pred_br_MPORT_6_mask) begin
      buf_pred_br[buf_pred_br_MPORT_6_addr] <= buf_pred_br_MPORT_6_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_br_MPORT_7_en & buf_pred_br_MPORT_7_mask) begin
      buf_pred_br[buf_pred_br_MPORT_7_addr] <= buf_pred_br_MPORT_7_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_br_MPORT_8_en & buf_pred_br_MPORT_8_mask) begin
      buf_pred_br[buf_pred_br_MPORT_8_addr] <= buf_pred_br_MPORT_8_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_br_MPORT_9_en & buf_pred_br_MPORT_9_mask) begin
      buf_pred_br[buf_pred_br_MPORT_9_addr] <= buf_pred_br_MPORT_9_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_br_MPORT_10_en & buf_pred_br_MPORT_10_mask) begin
      buf_pred_br[buf_pred_br_MPORT_10_addr] <= buf_pred_br_MPORT_10_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_br_MPORT_11_en & buf_pred_br_MPORT_11_mask) begin
      buf_pred_br[buf_pred_br_MPORT_11_addr] <= buf_pred_br_MPORT_11_data; // @[InstBuffer.scala 48:24]
    end
//     buf_pred_br_MPORT_2_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      buf_pred_br_MPORT_2_addr_pipe_0 <= next_deq_vec_0[2:0];
    end
//     buf_pred_br_MPORT_3_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      buf_pred_br_MPORT_3_addr_pipe_0 <= next_deq_vec_1[2:0];
    end
    if (buf_pred_bpc_MPORT_en & buf_pred_bpc_MPORT_mask) begin
      buf_pred_bpc[buf_pred_bpc_MPORT_addr] <= buf_pred_bpc_MPORT_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_bpc_MPORT_1_en & buf_pred_bpc_MPORT_1_mask) begin
      buf_pred_bpc[buf_pred_bpc_MPORT_1_addr] <= buf_pred_bpc_MPORT_1_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_bpc_MPORT_4_en & buf_pred_bpc_MPORT_4_mask) begin
      buf_pred_bpc[buf_pred_bpc_MPORT_4_addr] <= buf_pred_bpc_MPORT_4_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_bpc_MPORT_5_en & buf_pred_bpc_MPORT_5_mask) begin
      buf_pred_bpc[buf_pred_bpc_MPORT_5_addr] <= buf_pred_bpc_MPORT_5_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_bpc_MPORT_6_en & buf_pred_bpc_MPORT_6_mask) begin
      buf_pred_bpc[buf_pred_bpc_MPORT_6_addr] <= buf_pred_bpc_MPORT_6_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_bpc_MPORT_7_en & buf_pred_bpc_MPORT_7_mask) begin
      buf_pred_bpc[buf_pred_bpc_MPORT_7_addr] <= buf_pred_bpc_MPORT_7_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_bpc_MPORT_8_en & buf_pred_bpc_MPORT_8_mask) begin
      buf_pred_bpc[buf_pred_bpc_MPORT_8_addr] <= buf_pred_bpc_MPORT_8_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_bpc_MPORT_9_en & buf_pred_bpc_MPORT_9_mask) begin
      buf_pred_bpc[buf_pred_bpc_MPORT_9_addr] <= buf_pred_bpc_MPORT_9_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_bpc_MPORT_10_en & buf_pred_bpc_MPORT_10_mask) begin
      buf_pred_bpc[buf_pred_bpc_MPORT_10_addr] <= buf_pred_bpc_MPORT_10_data; // @[InstBuffer.scala 48:24]
    end
    if (buf_pred_bpc_MPORT_11_en & buf_pred_bpc_MPORT_11_mask) begin
      buf_pred_bpc[buf_pred_bpc_MPORT_11_addr] <= buf_pred_bpc_MPORT_11_data; // @[InstBuffer.scala 48:24]
    end
//     buf_pred_bpc_MPORT_2_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      buf_pred_bpc_MPORT_2_addr_pipe_0 <= next_deq_vec_0[2:0];
    end
//     buf_pred_bpc_MPORT_3_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      buf_pred_bpc_MPORT_3_addr_pipe_0 <= next_deq_vec_1[2:0];
    end
    if (reset) begin // @[InstBuffer.scala 50:24]
      enq_vec_0 <= 4'h0; // @[InstBuffer.scala 50:24]
    end else if (io_flush) begin // @[InstBuffer.scala 116:19]
      enq_vec_0 <= 4'h0; // @[InstBuffer.scala 118:13]
    end else if (_T_9 & _T_22) begin // @[InstBuffer.scala 94:36]
      enq_vec_0 <= next_enq_vec_0; // @[InstBuffer.scala 95:13]
    end
    if (reset) begin // @[InstBuffer.scala 50:24]
      enq_vec_1 <= 4'h1; // @[InstBuffer.scala 50:24]
    end else if (io_flush) begin // @[InstBuffer.scala 116:19]
      enq_vec_1 <= 4'h1; // @[InstBuffer.scala 118:13]
    end else if (_T_9 & _T_22) begin // @[InstBuffer.scala 94:36]
      enq_vec_1 <= next_enq_vec_1; // @[InstBuffer.scala 95:13]
    end
    if (reset) begin // @[InstBuffer.scala 51:24]
      deq_vec_0 <= 4'h0; // @[InstBuffer.scala 51:24]
    end else if (io_flush) begin // @[InstBuffer.scala 116:19]
      deq_vec_0 <= 4'h0; // @[InstBuffer.scala 119:13]
    end else begin
      deq_vec_0 <= next_deq_vec_0; // @[InstBuffer.scala 104:11]
    end
    if (reset) begin // @[InstBuffer.scala 51:24]
      deq_vec_1 <= 4'h1; // @[InstBuffer.scala 51:24]
    end else if (io_flush) begin // @[InstBuffer.scala 116:19]
      deq_vec_1 <= 4'h1; // @[InstBuffer.scala 119:13]
    end else begin
      deq_vec_1 <= next_deq_vec_1; // @[InstBuffer.scala 104:11]
    end
    enq_ready <= reset | _GEN_30; // @[InstBuffer.scala 58:{26,26}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    buf_pc[initvar] = _RAND_0[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    buf_inst[initvar] = _RAND_5[31:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    buf_pred_br[initvar] = _RAND_10[0:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    buf_pred_bpc[initvar] = _RAND_15[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
//   buf_pc_MPORT_2_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  buf_pc_MPORT_2_addr_pipe_0 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
//   buf_pc_MPORT_3_en_pipe_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  buf_pc_MPORT_3_addr_pipe_0 = _RAND_4[2:0];
  _RAND_6 = {1{`RANDOM}};
//   buf_inst_MPORT_2_en_pipe_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  buf_inst_MPORT_2_addr_pipe_0 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
//   buf_inst_MPORT_3_en_pipe_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  buf_inst_MPORT_3_addr_pipe_0 = _RAND_9[2:0];
  _RAND_11 = {1{`RANDOM}};
//   buf_pred_br_MPORT_2_en_pipe_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  buf_pred_br_MPORT_2_addr_pipe_0 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
//   buf_pred_br_MPORT_3_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  buf_pred_br_MPORT_3_addr_pipe_0 = _RAND_14[2:0];
  _RAND_16 = {1{`RANDOM}};
//   buf_pred_bpc_MPORT_2_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  buf_pred_bpc_MPORT_2_addr_pipe_0 = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
//   buf_pred_bpc_MPORT_3_en_pipe_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  buf_pred_bpc_MPORT_3_addr_pipe_0 = _RAND_19[2:0];
  _RAND_20 = {1{`RANDOM}};
  enq_vec_0 = _RAND_20[3:0];
  _RAND_21 = {1{`RANDOM}};
  enq_vec_1 = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  deq_vec_0 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  deq_vec_1 = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  enq_ready = _RAND_24[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_Decoder(
  input  [31:0] io_in__pc,
  input  [31:0] io_in__inst,
  input         io_in__pred_br,
  input  [31:0] io_in__pred_bpc,
  input         io_in__valid,
  input         io_in_valid,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_npc,
  output [31:0] io_out_inst,
  output [2:0]  io_out_fu_code,
  output [3:0]  io_out_alu_code,
  output [3:0]  io_out_jmp_code,
  output [1:0]  io_out_mem_code,
  output [1:0]  io_out_mem_size,
  output [2:0]  io_out_sys_code,
  output        io_out_w_type,
  output [1:0]  io_out_rs1_src,
  output [1:0]  io_out_rs2_src,
  output [4:0]  io_out_rs1_addr,
  output [4:0]  io_out_rs2_addr,
  output [4:0]  io_out_rd_addr,
  output        io_out_rd_en,
  output [31:0] io_out_imm,
  output        io_out_pred_br,
  output [31:0] io_out_pred_bpc
);
  wire [31:0] uop_npc = io_in__pc + 32'h4; // @[Decode.scala 63:23]
  wire [4:0] uop_rs1_addr = io_in__inst[19:15]; // @[Decode.scala 66:23]
  wire [4:0] uop_rs2_addr = io_in__inst[24:20]; // @[Decode.scala 67:23]
  wire [4:0] uop_rd_addr = io_in__inst[11:7]; // @[Decode.scala 68:22]
  wire [31:0] invInputs = ~io_in__inst; // @[pla.scala 77:21]
  wire  andMatrixInput_0 = io_in__inst[0]; // @[pla.scala 89:45]
  wire  andMatrixInput_1 = io_in__inst[1]; // @[pla.scala 89:45]
  wire  andMatrixInput_2 = invInputs[2]; // @[pla.scala 90:29]
  wire  andMatrixInput_3 = io_in__inst[3]; // @[pla.scala 89:45]
  wire  andMatrixInput_4 = io_in__inst[4]; // @[pla.scala 89:45]
  wire  andMatrixInput_5 = invInputs[5]; // @[pla.scala 90:29]
  wire  andMatrixInput_6 = invInputs[6]; // @[pla.scala 90:29]
  wire  andMatrixInput_7 = invInputs[12]; // @[pla.scala 90:29]
  wire  andMatrixInput_8 = invInputs[13]; // @[pla.scala 90:29]
  wire  andMatrixInput_9 = invInputs[14]; // @[pla.scala 90:29]
  wire [9:0] _T_5 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3,andMatrixInput_4,
    andMatrixInput_5,andMatrixInput_6,andMatrixInput_7,andMatrixInput_8,andMatrixInput_9}; // @[Cat.scala 30:58]
  wire  _T_6 = &_T_5; // @[pla.scala 97:74]
  wire  andMatrixInput_1_1 = io_in__inst[5]; // @[pla.scala 89:45]
  wire  andMatrixInput_3_1 = io_in__inst[13]; // @[pla.scala 89:45]
  wire [3:0] _T_7 = {andMatrixInput_2,andMatrixInput_1_1,andMatrixInput_7,andMatrixInput_3_1}; // @[Cat.scala 30:58]
  wire  _T_8 = &_T_7; // @[pla.scala 97:74]
  wire  andMatrixInput_1_2 = io_in__inst[12]; // @[pla.scala 89:45]
  wire  andMatrixInput_3_2 = io_in__inst[30]; // @[pla.scala 89:45]
  wire [3:0] _T_9 = {andMatrixInput_2,andMatrixInput_1_2,andMatrixInput_8,andMatrixInput_3_2}; // @[Cat.scala 30:58]
  wire  _T_10 = &_T_9; // @[pla.scala 97:74]
  wire  andMatrixInput_3_3 = invInputs[3]; // @[pla.scala 90:29]
  wire  andMatrixInput_6_1 = io_in__inst[6]; // @[pla.scala 89:45]
  wire [7:0] _T_11 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3_3,andMatrixInput_4,
    andMatrixInput_1_1,andMatrixInput_6_1,andMatrixInput_1_2}; // @[Cat.scala 30:58]
  wire  _T_12 = &_T_11; // @[pla.scala 97:74]
  wire  andMatrixInput_4_2 = invInputs[4]; // @[pla.scala 90:29]
  wire [7:0] _T_13 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3_3,andMatrixInput_4_2,
    andMatrixInput_5,andMatrixInput_6,andMatrixInput_9}; // @[Cat.scala 30:58]
  wire  _T_14 = &_T_13; // @[pla.scala 97:74]
  wire  andMatrixInput_8_1 = io_in__inst[14]; // @[pla.scala 89:45]
  wire  andMatrixInput_9_1 = invInputs[25]; // @[pla.scala 90:29]
  wire  andMatrixInput_10 = invInputs[26]; // @[pla.scala 90:29]
  wire  andMatrixInput_11 = invInputs[27]; // @[pla.scala 90:29]
  wire  andMatrixInput_12 = invInputs[28]; // @[pla.scala 90:29]
  wire  andMatrixInput_13 = invInputs[29]; // @[pla.scala 90:29]
  wire  andMatrixInput_14 = invInputs[31]; // @[pla.scala 90:29]
  wire [6:0] lo_5 = {andMatrixInput_8_1,andMatrixInput_9_1,andMatrixInput_10,andMatrixInput_11,andMatrixInput_12,
    andMatrixInput_13,andMatrixInput_14}; // @[Cat.scala 30:58]
  wire [1:0] hi_hi_lo = {andMatrixInput_2,andMatrixInput_3}; // @[Cat.scala 30:58]
  wire [14:0] _T_15 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3,andMatrixInput_4,
    andMatrixInput_6,andMatrixInput_1_2,andMatrixInput_8,lo_5}; // @[Cat.scala 30:58]
  wire  _T_16 = &_T_15; // @[pla.scala 97:74]
  wire  _T_17 = &andMatrixInput_5; // @[pla.scala 97:74]
  wire  andMatrixInput_10_1 = invInputs[30]; // @[pla.scala 90:29]
  wire [5:0] lo_6 = {andMatrixInput_10,andMatrixInput_11,andMatrixInput_12,andMatrixInput_13,andMatrixInput_10_1,
    andMatrixInput_14}; // @[Cat.scala 30:58]
  wire [11:0] _T_18 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_3_3,andMatrixInput_4,andMatrixInput_5,
    andMatrixInput_6,lo_6}; // @[Cat.scala 30:58]
  wire  _T_19 = &_T_18; // @[pla.scala 97:74]
  wire [7:0] _T_20 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3_3,andMatrixInput_4,
    andMatrixInput_1_1,andMatrixInput_6_1,andMatrixInput_3_1}; // @[Cat.scala 30:58]
  wire  _T_21 = &_T_20; // @[pla.scala 97:74]
  wire  andMatrixInput_7_6 = invInputs[7]; // @[pla.scala 90:29]
  wire  andMatrixInput_8_3 = invInputs[8]; // @[pla.scala 90:29]
  wire  andMatrixInput_9_3 = invInputs[9]; // @[pla.scala 90:29]
  wire  andMatrixInput_10_2 = invInputs[10]; // @[pla.scala 90:29]
  wire  andMatrixInput_11_2 = invInputs[11]; // @[pla.scala 90:29]
  wire  andMatrixInput_13_1 = invInputs[15]; // @[pla.scala 90:29]
  wire  andMatrixInput_14_1 = invInputs[16]; // @[pla.scala 90:29]
  wire  andMatrixInput_15 = invInputs[17]; // @[pla.scala 90:29]
  wire  andMatrixInput_16 = invInputs[18]; // @[pla.scala 90:29]
  wire  andMatrixInput_17 = invInputs[19]; // @[pla.scala 90:29]
  wire  andMatrixInput_18 = invInputs[20]; // @[pla.scala 90:29]
  wire  andMatrixInput_19 = io_in__inst[21]; // @[pla.scala 89:45]
  wire  andMatrixInput_20 = invInputs[22]; // @[pla.scala 90:29]
  wire  andMatrixInput_21 = invInputs[23]; // @[pla.scala 90:29]
  wire  andMatrixInput_22 = invInputs[24]; // @[pla.scala 90:29]
  wire  andMatrixInput_26 = io_in__inst[28]; // @[pla.scala 89:45]
  wire  andMatrixInput_27 = io_in__inst[29]; // @[pla.scala 89:45]
  wire [6:0] lo_lo_6 = {andMatrixInput_9_1,andMatrixInput_10,andMatrixInput_11,andMatrixInput_26,andMatrixInput_27,
    andMatrixInput_10_1,andMatrixInput_14}; // @[Cat.scala 30:58]
  wire [14:0] lo_8 = {andMatrixInput_15,andMatrixInput_16,andMatrixInput_17,andMatrixInput_18,andMatrixInput_19,
    andMatrixInput_20,andMatrixInput_21,andMatrixInput_22,lo_lo_6}; // @[Cat.scala 30:58]
  wire [6:0] hi_lo_6 = {andMatrixInput_8_3,andMatrixInput_9_3,andMatrixInput_10_2,andMatrixInput_11_2,andMatrixInput_9,
    andMatrixInput_13_1,andMatrixInput_14_1}; // @[Cat.scala 30:58]
  wire [29:0] _T_22 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3_3,andMatrixInput_4,
    andMatrixInput_1_1,andMatrixInput_6_1,andMatrixInput_7_6,hi_lo_6,lo_8}; // @[Cat.scala 30:58]
  wire  _T_23 = &_T_22; // @[pla.scala 97:74]
  wire [3:0] _T_24 = {andMatrixInput_2,andMatrixInput_7,andMatrixInput_8,andMatrixInput_8_1}; // @[Cat.scala 30:58]
  wire  _T_25 = &_T_24; // @[pla.scala 97:74]
  wire  andMatrixInput_0_11 = io_in__inst[2]; // @[pla.scala 89:45]
  wire [1:0] _T_26 = {andMatrixInput_0_11,andMatrixInput_5}; // @[Cat.scala 30:58]
  wire  _T_27 = &_T_26; // @[pla.scala 97:74]
  wire [2:0] _T_28 = {andMatrixInput_3_3,andMatrixInput_6_1,andMatrixInput_18}; // @[Cat.scala 30:58]
  wire  _T_29 = &_T_28; // @[pla.scala 97:74]
  wire [5:0] _T_30 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_0_11,andMatrixInput_3_3,andMatrixInput_4,
    andMatrixInput_6}; // @[Cat.scala 30:58]
  wire  _T_31 = &_T_30; // @[pla.scala 97:74]
  wire [2:0] _T_32 = {andMatrixInput_4,andMatrixInput_6_1,andMatrixInput_8_1}; // @[Cat.scala 30:58]
  wire  _T_33 = &_T_32; // @[pla.scala 97:74]
  wire [6:0] lo_11 = {andMatrixInput_9,andMatrixInput_9_1,andMatrixInput_10,andMatrixInput_11,andMatrixInput_12,
    andMatrixInput_13,andMatrixInput_14}; // @[Cat.scala 30:58]
  wire [13:0] _T_34 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_4,andMatrixInput_6,
    andMatrixInput_7,andMatrixInput_8,lo_11}; // @[Cat.scala 30:58]
  wire  _T_35 = &_T_34; // @[pla.scala 97:74]
  wire [5:0] lo_12 = {andMatrixInput_8_1,andMatrixInput_10,andMatrixInput_11,andMatrixInput_12,andMatrixInput_13,
    andMatrixInput_14}; // @[Cat.scala 30:58]
  wire [11:0] _T_36 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_3_3,andMatrixInput_4,andMatrixInput_5,
    andMatrixInput_6,lo_12}; // @[Cat.scala 30:58]
  wire  _T_37 = &_T_36; // @[pla.scala 97:74]
  wire [6:0] _T_38 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3_3,andMatrixInput_5,
    andMatrixInput_6,andMatrixInput_7}; // @[Cat.scala 30:58]
  wire  _T_39 = &_T_38; // @[pla.scala 97:74]
  wire [2:0] _T_40 = {andMatrixInput_2,andMatrixInput_4,andMatrixInput_6}; // @[Cat.scala 30:58]
  wire  _T_41 = &_T_40; // @[pla.scala 97:74]
  wire [2:0] _T_42 = {andMatrixInput_1_2,andMatrixInput_8_1,andMatrixInput_10_1}; // @[Cat.scala 30:58]
  wire  _T_43 = &_T_42; // @[pla.scala 97:74]
  wire [3:0] _T_44 = {andMatrixInput_2,andMatrixInput_1_1,andMatrixInput_1_2,andMatrixInput_3_1}; // @[Cat.scala 30:58]
  wire  _T_45 = &_T_44; // @[pla.scala 97:74]
  wire [8:0] _T_46 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_0_11,andMatrixInput_4_2,andMatrixInput_1_1,
    andMatrixInput_6_1,andMatrixInput_7,andMatrixInput_8,andMatrixInput_9}; // @[Cat.scala 30:58]
  wire  _T_47 = &_T_46; // @[pla.scala 97:74]
  wire  andMatrixInput_18_1 = io_in__inst[20]; // @[pla.scala 89:45]
  wire  andMatrixInput_19_1 = invInputs[21]; // @[pla.scala 90:29]
  wire  andMatrixInput_20_1 = io_in__inst[22]; // @[pla.scala 89:45]
  wire [6:0] lo_lo_10 = {andMatrixInput_9_1,andMatrixInput_10,andMatrixInput_11,andMatrixInput_26,andMatrixInput_13,
    andMatrixInput_10_1,andMatrixInput_14}; // @[Cat.scala 30:58]
  wire [14:0] lo_16 = {andMatrixInput_15,andMatrixInput_16,andMatrixInput_17,andMatrixInput_18_1,andMatrixInput_19_1,
    andMatrixInput_20_1,andMatrixInput_21,andMatrixInput_22,lo_lo_10}; // @[Cat.scala 30:58]
  wire [29:0] _T_48 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3_3,andMatrixInput_4,
    andMatrixInput_1_1,andMatrixInput_6_1,andMatrixInput_7_6,hi_lo_6,lo_16}; // @[Cat.scala 30:58]
  wire  _T_49 = &_T_48; // @[pla.scala 97:74]
  wire [3:0] _T_50 = {andMatrixInput_4_2,andMatrixInput_5,andMatrixInput_8,andMatrixInput_9}; // @[Cat.scala 30:58]
  wire  _T_51 = &_T_50; // @[pla.scala 97:74]
  wire [13:0] _T_52 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_4,andMatrixInput_6,
    andMatrixInput_1_2,andMatrixInput_8,lo_5}; // @[Cat.scala 30:58]
  wire  _T_53 = &_T_52; // @[pla.scala 97:74]
  wire [1:0] _T_54 = {andMatrixInput_0_11,andMatrixInput_3}; // @[Cat.scala 30:58]
  wire  _T_55 = &_T_54; // @[pla.scala 97:74]
  wire [6:0] _T_56 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3_3,andMatrixInput_4_2,
    andMatrixInput_6,andMatrixInput_9}; // @[Cat.scala 30:58]
  wire  _T_57 = &_T_56; // @[pla.scala 97:74]
  wire [7:0] _T_58 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3_3,andMatrixInput_4_2,
    andMatrixInput_1_1,andMatrixInput_6_1,andMatrixInput_8_1}; // @[Cat.scala 30:58]
  wire  _T_59 = &_T_58; // @[pla.scala 97:74]
  wire [7:0] _T_60 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3_3,andMatrixInput_4_2,
    andMatrixInput_5,andMatrixInput_6,andMatrixInput_8}; // @[Cat.scala 30:58]
  wire  _T_61 = &_T_60; // @[pla.scala 97:74]
  wire [6:0] lo_lo_14 = {andMatrixInput_9_1,andMatrixInput_10,andMatrixInput_11,andMatrixInput_12,andMatrixInput_13,
    andMatrixInput_10_1,andMatrixInput_14}; // @[Cat.scala 30:58]
  wire [14:0] lo_22 = {andMatrixInput_15,andMatrixInput_16,andMatrixInput_17,andMatrixInput_18,andMatrixInput_19_1,
    andMatrixInput_20,andMatrixInput_21,andMatrixInput_22,lo_lo_14}; // @[Cat.scala 30:58]
  wire [6:0] hi_lo_16 = {andMatrixInput_10_2,andMatrixInput_11_2,andMatrixInput_7,andMatrixInput_8,andMatrixInput_9,
    andMatrixInput_13_1,andMatrixInput_14_1}; // @[Cat.scala 30:58]
  wire [29:0] _T_62 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_1_1,andMatrixInput_6_1,
    andMatrixInput_7_6,andMatrixInput_8_3,andMatrixInput_9_3,hi_lo_16,lo_22}; // @[Cat.scala 30:58]
  wire  _T_63 = &_T_62; // @[pla.scala 97:74]
  wire [3:0] _T_64 = {andMatrixInput_3_3,andMatrixInput_6_1,andMatrixInput_7,andMatrixInput_9}; // @[Cat.scala 30:58]
  wire  _T_65 = &_T_64; // @[pla.scala 97:74]
  wire [4:0] _T_66 = {andMatrixInput_2,andMatrixInput_4_2,andMatrixInput_1_2,andMatrixInput_8,andMatrixInput_8_1}; // @[Cat.scala 30:58]
  wire  _T_67 = &_T_66; // @[pla.scala 97:74]
  wire [6:0] _T_68 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_0_11,andMatrixInput_3,andMatrixInput_4_2,
    andMatrixInput_1_1,andMatrixInput_6_1}; // @[Cat.scala 30:58]
  wire  _T_69 = &_T_68; // @[pla.scala 97:74]
  wire [7:0] _T_70 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3_3,andMatrixInput_4_2,
    andMatrixInput_1_1,andMatrixInput_6_1,andMatrixInput_8}; // @[Cat.scala 30:58]
  wire  _T_71 = &_T_70; // @[pla.scala 97:74]
  wire [1:0] _T_72 = {andMatrixInput_8,andMatrixInput_19}; // @[Cat.scala 30:58]
  wire  _T_73 = &_T_72; // @[pla.scala 97:74]
  wire [14:0] _T_74 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3,andMatrixInput_4,
    andMatrixInput_6,andMatrixInput_1_2,andMatrixInput_8,lo_lo_14}; // @[Cat.scala 30:58]
  wire  _T_75 = &_T_74; // @[pla.scala 97:74]
  wire [3:0] _T_76 = {andMatrixInput_4,andMatrixInput_6_1,andMatrixInput_1_2,andMatrixInput_9}; // @[Cat.scala 30:58]
  wire  _T_77 = &_T_76; // @[pla.scala 97:74]
  wire [2:0] _T_78 = {andMatrixInput_2,andMatrixInput_3_1,andMatrixInput_8_1}; // @[Cat.scala 30:58]
  wire  _T_79 = &_T_78; // @[pla.scala 97:74]
  wire [3:0] _T_80 = {andMatrixInput_2,andMatrixInput_5,andMatrixInput_1_2,andMatrixInput_3_1}; // @[Cat.scala 30:58]
  wire  _T_81 = &_T_80; // @[pla.scala 97:74]
  wire [2:0] _T_82 = {andMatrixInput_1_2,andMatrixInput_3_1,andMatrixInput_8_1}; // @[Cat.scala 30:58]
  wire  _T_83 = &_T_82; // @[pla.scala 97:74]
  wire [6:0] _T_84 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_3_3,andMatrixInput_4,andMatrixInput_5,
    andMatrixInput_6,andMatrixInput_3_1}; // @[Cat.scala 30:58]
  wire  _T_85 = &_T_84; // @[pla.scala 97:74]
  wire [9:0] _T_86 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_0_11,andMatrixInput_3,andMatrixInput_4_2,
    andMatrixInput_5,andMatrixInput_6,andMatrixInput_1_2,andMatrixInput_8,andMatrixInput_9}; // @[Cat.scala 30:58]
  wire  _T_87 = &_T_86; // @[pla.scala 97:74]
  wire [3:0] _T_88 = {andMatrixInput_2,andMatrixInput_5,andMatrixInput_7,andMatrixInput_9}; // @[Cat.scala 30:58]
  wire  _T_89 = &_T_88; // @[pla.scala 97:74]
  wire [3:0] _T_90 = {andMatrixInput_2,andMatrixInput_1_1,andMatrixInput_1_2,andMatrixInput_8}; // @[Cat.scala 30:58]
  wire  _T_91 = &_T_90; // @[pla.scala 97:74]
  wire [2:0] _T_92 = {andMatrixInput_2,andMatrixInput_7,andMatrixInput_3_1}; // @[Cat.scala 30:58]
  wire  _T_93 = &_T_92; // @[pla.scala 97:74]
  wire [3:0] _T_94 = {andMatrixInput_4,andMatrixInput_7,andMatrixInput_9,andMatrixInput_10_1}; // @[Cat.scala 30:58]
  wire  _T_95 = &_T_94; // @[pla.scala 97:74]
  wire [4:0] _T_96 = {andMatrixInput_2,andMatrixInput_3_3,andMatrixInput_4,andMatrixInput_1_2,andMatrixInput_8}; // @[Cat.scala 30:58]
  wire  _T_97 = &_T_96; // @[pla.scala 97:74]
  wire  _T_99 = &hi_hi_lo; // @[pla.scala 97:74]
  wire [2:0] _T_100 = {andMatrixInput_3_3,andMatrixInput_4_2,andMatrixInput_6_1}; // @[Cat.scala 30:58]
  wire  _T_101 = &_T_100; // @[pla.scala 97:74]
  wire [1:0] _T_102 = {andMatrixInput_0_11,andMatrixInput_4}; // @[Cat.scala 30:58]
  wire  _T_103 = &_T_102; // @[pla.scala 97:74]
  wire [3:0] _T_104 = {andMatrixInput_2,andMatrixInput_6_1,andMatrixInput_3_1,andMatrixInput_9}; // @[Cat.scala 30:58]
  wire  _T_105 = &_T_104; // @[pla.scala 97:74]
  wire [14:0] _T_106 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3,andMatrixInput_4,
    andMatrixInput_6,andMatrixInput_7,andMatrixInput_8,lo_11}; // @[Cat.scala 30:58]
  wire  _T_107 = &_T_106; // @[pla.scala 97:74]
  wire [2:0] _T_108 = {andMatrixInput_2,andMatrixInput_1_2,andMatrixInput_8}; // @[Cat.scala 30:58]
  wire  _T_109 = &_T_108; // @[pla.scala 97:74]
  wire [11:0] _T_110 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_3_3,andMatrixInput_4,andMatrixInput_6,
    andMatrixInput_9_1,lo_6}; // @[Cat.scala 30:58]
  wire  _T_111 = &_T_110; // @[pla.scala 97:74]
  wire [3:0] _T_112 = {andMatrixInput_2,andMatrixInput_1_1,andMatrixInput_7,andMatrixInput_8}; // @[Cat.scala 30:58]
  wire  _T_113 = &_T_112; // @[pla.scala 97:74]
  wire [2:0] _T_114 = {andMatrixInput_2,andMatrixInput_4_2,andMatrixInput_6}; // @[Cat.scala 30:58]
  wire  _T_115 = &_T_114; // @[pla.scala 97:74]
  wire [2:0] _T_116 = {andMatrixInput_2,andMatrixInput_1_1,andMatrixInput_3_2}; // @[Cat.scala 30:58]
  wire  _T_117 = &_T_116; // @[pla.scala 97:74]
  wire [9:0] _orMatrixOutputs_T = {_T_25,_T_33,_T_51,_T_55,_T_67,_T_79,_T_81,_T_89,_T_99,_T_101}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_1 = |_orMatrixOutputs_T; // @[pla.scala 113:41]
  wire [4:0] _orMatrixOutputs_T_2 = {_T_8,_T_45,_T_91,_T_97,_T_113}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_3 = |_orMatrixOutputs_T_2; // @[pla.scala 113:41]
  wire [3:0] _orMatrixOutputs_T_4 = {_T_33,_T_55,_T_97,_T_103}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_5 = |_orMatrixOutputs_T_4; // @[pla.scala 113:41]
  wire [7:0] orMatrixOutputs_lo_3 = {_T_39,_T_47,_T_53,_T_61,_T_69,_T_75,_T_85,_T_111}; // @[Cat.scala 30:58]
  wire [15:0] _orMatrixOutputs_T_6 = {_T_6,_T_12,_T_14,_T_19,_T_21,_T_31,_T_35,_T_37,orMatrixOutputs_lo_3}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_7 = |_orMatrixOutputs_T_6; // @[pla.scala 113:41]
  wire [4:0] _orMatrixOutputs_T_8 = {_T_8,_T_45,_T_65,_T_91,_T_113}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_9 = |_orMatrixOutputs_T_8; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_10 = {_T_17,_T_55,_T_103}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_11 = |_orMatrixOutputs_T_10; // @[pla.scala 113:41]
  wire [6:0] _orMatrixOutputs_T_12 = {_T_27,_T_41,_T_55,_T_77,_T_101,_T_105,_T_115}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_13 = |_orMatrixOutputs_T_12; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_14 = {_T_27,_T_33,_T_55}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_15 = |_orMatrixOutputs_T_14; // @[pla.scala 113:41]
  wire [3:0] _orMatrixOutputs_T_16 = {_T_6,_T_16,_T_75,_T_107}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_17 = |_orMatrixOutputs_T_16; // @[pla.scala 113:41]
  wire [3:0] _orMatrixOutputs_T_18 = {_T_27,_T_45,_T_73,_T_91}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_19 = |_orMatrixOutputs_T_18; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_20 = {_T_8,_T_27,_T_45}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_21 = |_orMatrixOutputs_T_20; // @[pla.scala 113:41]
  wire [1:0] _orMatrixOutputs_T_22 = {_T_27,_T_113}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_23 = |_orMatrixOutputs_T_22; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_24 = {_T_45,_T_81,_T_109}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_25 = |_orMatrixOutputs_T_24; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_26 = {_T_45,_T_81,_T_93}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_27 = |_orMatrixOutputs_T_26; // @[pla.scala 113:41]
  wire [5:0] _orMatrixOutputs_T_28 = {_T_8,_T_45,_T_51,_T_89,_T_91,_T_113}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_29 = |_orMatrixOutputs_T_28; // @[pla.scala 113:41]
  wire [7:0] _orMatrixOutputs_T_30 = {_T_8,_T_25,_T_45,_T_67,_T_79,_T_81,_T_91,_T_113}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_31 = |_orMatrixOutputs_T_30; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_32 = {_T_8,_T_55,_T_113}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_33 = |_orMatrixOutputs_T_32; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_34 = {_T_8,_T_65,_T_67}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_35 = |_orMatrixOutputs_T_34; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_36 = {_T_8,_T_25,_T_91}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_37 = |_orMatrixOutputs_T_36; // @[pla.scala 113:41]
  wire  _orMatrixOutputs_T_38 = |_T_45; // @[pla.scala 113:41]
  wire [5:0] _orMatrixOutputs_T_39 = {_T_25,_T_43,_T_83,_T_89,_T_95,_T_103}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_40 = |_orMatrixOutputs_T_39; // @[pla.scala 113:41]
  wire [3:0] _orMatrixOutputs_T_41 = {_T_10,_T_79,_T_93,_T_117}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_42 = |_orMatrixOutputs_T_41; // @[pla.scala 113:41]
  wire [3:0] _orMatrixOutputs_T_43 = {_T_25,_T_45,_T_79,_T_81}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_44 = |_orMatrixOutputs_T_43; // @[pla.scala 113:41]
  wire  _orMatrixOutputs_T_45 = |_T_109; // @[pla.scala 113:41]
  wire [7:0] _orMatrixOutputs_T_46 = {_T_27,_T_33,_T_41,_T_77,_T_95,_T_99,_T_103,_T_105}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_47 = |_orMatrixOutputs_T_46; // @[pla.scala 113:41]
  wire [5:0] _orMatrixOutputs_T_48 = {_T_29,_T_33,_T_55,_T_77,_T_101,_T_105}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_49 = |_orMatrixOutputs_T_48; // @[pla.scala 113:41]
  wire  _orMatrixOutputs_T_50 = |_T_115; // @[pla.scala 113:41]
  wire [4:0] orMatrixOutputs_lo_lo_4 = {_T_71,_T_75,_T_85,_T_87,_T_111}; // @[Cat.scala 30:58]
  wire [10:0] orMatrixOutputs_lo_15 = {_T_53,_T_57,_T_59,_T_61,_T_63,_T_69,orMatrixOutputs_lo_lo_4}; // @[Cat.scala 30:58]
  wire [4:0] orMatrixOutputs_hi_lo_5 = {_T_35,_T_37,_T_39,_T_47,_T_49}; // @[Cat.scala 30:58]
  wire [21:0] _orMatrixOutputs_T_51 = {_T_6,_T_12,_T_19,_T_21,_T_23,_T_31,orMatrixOutputs_hi_lo_5,orMatrixOutputs_lo_15}
    ; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_52 = |_orMatrixOutputs_T_51; // @[pla.scala 113:41]
  wire [6:0] orMatrixOutputs_lo_lo_5 = {_orMatrixOutputs_T_13,_orMatrixOutputs_T_11,_orMatrixOutputs_T_9,
    _orMatrixOutputs_T_7,_orMatrixOutputs_T_5,_orMatrixOutputs_T_3,_orMatrixOutputs_T_1}; // @[Cat.scala 30:58]
  wire [13:0] orMatrixOutputs_lo_16 = {_orMatrixOutputs_T_27,_orMatrixOutputs_T_25,_orMatrixOutputs_T_23,
    _orMatrixOutputs_T_21,_orMatrixOutputs_T_19,_orMatrixOutputs_T_17,_orMatrixOutputs_T_15,orMatrixOutputs_lo_lo_5}; // @[Cat.scala 30:58]
  wire [6:0] orMatrixOutputs_hi_lo_6 = {_orMatrixOutputs_T_40,_orMatrixOutputs_T_38,_orMatrixOutputs_T_37,
    _orMatrixOutputs_T_35,_orMatrixOutputs_T_33,_orMatrixOutputs_T_31,_orMatrixOutputs_T_29}; // @[Cat.scala 30:58]
  wire [27:0] orMatrixOutputs = {_orMatrixOutputs_T_52,_orMatrixOutputs_T_50,_orMatrixOutputs_T_49,_orMatrixOutputs_T_47
    ,_orMatrixOutputs_T_45,_orMatrixOutputs_T_44,_orMatrixOutputs_T_42,orMatrixOutputs_hi_lo_6,orMatrixOutputs_lo_16}; // @[Cat.scala 30:58]
  wire [6:0] invMatrixOutputs_lo_lo = {orMatrixOutputs[6],orMatrixOutputs[5],orMatrixOutputs[4],orMatrixOutputs[3],
    orMatrixOutputs[2],orMatrixOutputs[1],orMatrixOutputs[0]}; // @[Cat.scala 30:58]
  wire [13:0] invMatrixOutputs_lo = {orMatrixOutputs[13],orMatrixOutputs[12],orMatrixOutputs[11],orMatrixOutputs[10],
    orMatrixOutputs[9],orMatrixOutputs[8],orMatrixOutputs[7],invMatrixOutputs_lo_lo}; // @[Cat.scala 30:58]
  wire [6:0] invMatrixOutputs_hi_lo = {orMatrixOutputs[20],orMatrixOutputs[19],orMatrixOutputs[18],orMatrixOutputs[17],
    orMatrixOutputs[16],orMatrixOutputs[15],orMatrixOutputs[14]}; // @[Cat.scala 30:58]
  wire [27:0] invMatrixOutputs = {orMatrixOutputs[27],orMatrixOutputs[26],orMatrixOutputs[25],orMatrixOutputs[24],
    orMatrixOutputs[23],orMatrixOutputs[22],orMatrixOutputs[21],invMatrixOutputs_hi_lo,invMatrixOutputs_lo}; // @[Cat.scala 30:58]
  wire [1:0] uop_rs2_src = invMatrixOutputs[5:4]; // @[MicroOp.scala 56:20]
  wire [1:0] uop_rs1_src = invMatrixOutputs[7:6]; // @[MicroOp.scala 56:20]
  wire  uop_w_type = invMatrixOutputs[8]; // @[MicroOp.scala 54:20]
  wire [2:0] uop_sys_code = invMatrixOutputs[11:9]; // @[MicroOp.scala 56:20]
  wire [1:0] uop_mem_size = invMatrixOutputs[13:12]; // @[MicroOp.scala 56:20]
  wire [1:0] uop_mem_code = invMatrixOutputs[15:14]; // @[MicroOp.scala 56:20]
  wire [3:0] uop_jmp_code = invMatrixOutputs[19:16]; // @[MicroOp.scala 56:20]
  wire [3:0] uop_alu_code = invMatrixOutputs[23:20]; // @[MicroOp.scala 56:20]
  wire [2:0] uop_fu_code = invMatrixOutputs[26:24]; // @[MicroOp.scala 56:20]
  wire  uop_valid = invMatrixOutputs[27]; // @[MicroOp.scala 54:20]
  wire  uop_rd_en = invMatrixOutputs[3] & uop_rd_addr != 5'h0; // @[MicroOp.scala 61:24]
  wire [20:0] _T_135 = io_in__inst[31] ? 21'h1fffff : 21'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_137 = {_T_135,io_in__inst[30:20]}; // @[Cat.scala 30:58]
  wire [31:0] _T_143 = {_T_135,io_in__inst[30:25],uop_rd_addr}; // @[Cat.scala 30:58]
  wire [19:0] _T_146 = io_in__inst[31] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_150 = {_T_146,io_in__inst[7],io_in__inst[30:25],io_in__inst[11:8],1'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_153 = {io_in__inst[31:12],12'h0}; // @[Cat.scala 30:58]
  wire [11:0] _T_156 = io_in__inst[31] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_160 = {_T_156,io_in__inst[19:12],andMatrixInput_18_1,io_in__inst[30:21],1'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_163 = {27'h0,uop_rs2_addr}; // @[Cat.scala 30:58]
  wire [31:0] _T_166 = {26'h0,io_in__inst[25:20]}; // @[Cat.scala 30:58]
  wire [31:0] _T_167 = uop_w_type ? _T_163 : _T_166; // @[MicroOp.scala 68:24]
  wire [31:0] _T_170 = {27'h0,uop_rs1_addr}; // @[Cat.scala 30:58]
  wire [31:0] _T_172 = 3'h1 == invMatrixOutputs[2:0] ? _T_137 : 32'h0; // @[Mux.scala 80:57]
  wire [31:0] _T_174 = 3'h2 == invMatrixOutputs[2:0] ? _T_143 : _T_172; // @[Mux.scala 80:57]
  wire [31:0] _T_176 = 3'h3 == invMatrixOutputs[2:0] ? _T_150 : _T_174; // @[Mux.scala 80:57]
  wire [31:0] _T_178 = 3'h4 == invMatrixOutputs[2:0] ? _T_153 : _T_176; // @[Mux.scala 80:57]
  wire [31:0] _T_180 = 3'h5 == invMatrixOutputs[2:0] ? _T_160 : _T_178; // @[Mux.scala 80:57]
  wire [31:0] _T_182 = 3'h6 == invMatrixOutputs[2:0] ? _T_167 : _T_180; // @[Mux.scala 80:57]
  wire [31:0] uop_imm = 3'h7 == invMatrixOutputs[2:0] ? _T_170 : _T_182; // @[Mux.scala 80:57]
  assign io_out_valid = io_in_valid & io_in__valid & uop_valid; // @[Decode.scala 79:16]
  assign io_out_pc = io_in_valid & io_in__valid ? io_in__pc : 32'h0; // @[Decode.scala 79:16]
  assign io_out_npc = io_in_valid & io_in__valid ? uop_npc : 32'h0; // @[Decode.scala 79:16]
  assign io_out_inst = io_in_valid & io_in__valid ? io_in__inst : 32'h0; // @[Decode.scala 79:16]
  assign io_out_fu_code = io_in_valid & io_in__valid ? uop_fu_code : 3'h0; // @[Decode.scala 79:16]
  assign io_out_alu_code = io_in_valid & io_in__valid ? uop_alu_code : 4'h0; // @[Decode.scala 79:16]
  assign io_out_jmp_code = io_in_valid & io_in__valid ? uop_jmp_code : 4'h0; // @[Decode.scala 79:16]
  assign io_out_mem_code = io_in_valid & io_in__valid ? uop_mem_code : 2'h0; // @[Decode.scala 79:16]
  assign io_out_mem_size = io_in_valid & io_in__valid ? uop_mem_size : 2'h0; // @[Decode.scala 79:16]
  assign io_out_sys_code = io_in_valid & io_in__valid ? uop_sys_code : 3'h0; // @[Decode.scala 79:16]
  assign io_out_w_type = io_in_valid & io_in__valid & uop_w_type; // @[Decode.scala 79:16]
  assign io_out_rs1_src = io_in_valid & io_in__valid ? uop_rs1_src : 2'h0; // @[Decode.scala 79:16]
  assign io_out_rs2_src = io_in_valid & io_in__valid ? uop_rs2_src : 2'h0; // @[Decode.scala 79:16]
  assign io_out_rs1_addr = io_in_valid & io_in__valid ? uop_rs1_addr : 5'h0; // @[Decode.scala 79:16]
  assign io_out_rs2_addr = io_in_valid & io_in__valid ? uop_rs2_addr : 5'h0; // @[Decode.scala 79:16]
  assign io_out_rd_addr = io_in_valid & io_in__valid ? uop_rd_addr : 5'h0; // @[Decode.scala 79:16]
  assign io_out_rd_en = io_in_valid & io_in__valid & uop_rd_en; // @[Decode.scala 79:16]
  assign io_out_imm = io_in_valid & io_in__valid ? uop_imm : 32'h0; // @[Decode.scala 79:16]
  assign io_out_pred_br = io_in_valid & io_in__valid & io_in__pred_br; // @[Decode.scala 79:16]
  assign io_out_pred_bpc = io_in_valid & io_in__valid ? io_in__pred_bpc : 32'h0; // @[Decode.scala 79:16]
endmodule
module ysyx_210128_Decoder_1(
  input  [31:0] io_in__pc,
  input  [31:0] io_in__inst,
  input         io_in__pred_br,
  input  [31:0] io_in__pred_bpc,
  input         io_in__valid,
  input         io_in_valid,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_npc,
  output [31:0] io_out_inst,
  output [2:0]  io_out_fu_code,
  output [3:0]  io_out_alu_code,
  output [3:0]  io_out_jmp_code,
  output [1:0]  io_out_mem_code,
  output [1:0]  io_out_mem_size,
  output [2:0]  io_out_sys_code,
  output        io_out_w_type,
  output [1:0]  io_out_rs1_src,
  output [1:0]  io_out_rs2_src,
  output [4:0]  io_out_rs1_addr,
  output [4:0]  io_out_rs2_addr,
  output [4:0]  io_out_rd_addr,
  output        io_out_rd_en,
  output [31:0] io_out_imm,
  output        io_out_pred_br,
  output [31:0] io_out_pred_bpc
);
  wire [31:0] uop_npc = io_in__pc + 32'h4; // @[Decode.scala 63:23]
  wire [4:0] uop_rs1_addr = io_in__inst[19:15]; // @[Decode.scala 66:23]
  wire [4:0] uop_rs2_addr = io_in__inst[24:20]; // @[Decode.scala 67:23]
  wire [4:0] uop_rd_addr = io_in__inst[11:7]; // @[Decode.scala 68:22]
  wire [31:0] invInputs = ~io_in__inst; // @[pla.scala 77:21]
  wire  andMatrixInput_0 = invInputs[3]; // @[pla.scala 90:29]
  wire  andMatrixInput_1 = io_in__inst[6]; // @[pla.scala 89:45]
  wire  andMatrixInput_2 = invInputs[12]; // @[pla.scala 90:29]
  wire  andMatrixInput_3 = invInputs[14]; // @[pla.scala 90:29]
  wire [3:0] _T_5 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2,andMatrixInput_3}; // @[Cat.scala 30:58]
  wire  _T_6 = &_T_5; // @[pla.scala 97:74]
  wire  andMatrixInput_0_1 = invInputs[2]; // @[pla.scala 90:29]
  wire  andMatrixInput_2_1 = io_in__inst[13]; // @[pla.scala 89:45]
  wire [2:0] _T_7 = {andMatrixInput_0_1,andMatrixInput_2,andMatrixInput_2_1}; // @[Cat.scala 30:58]
  wire  _T_8 = &_T_7; // @[pla.scala 97:74]
  wire  andMatrixInput_0_2 = io_in__inst[0]; // @[pla.scala 89:45]
  wire  andMatrixInput_1_2 = io_in__inst[1]; // @[pla.scala 89:45]
  wire  andMatrixInput_3_1 = io_in__inst[4]; // @[pla.scala 89:45]
  wire  andMatrixInput_4 = invInputs[6]; // @[pla.scala 90:29]
  wire  andMatrixInput_6 = invInputs[13]; // @[pla.scala 90:29]
  wire  andMatrixInput_8 = invInputs[25]; // @[pla.scala 90:29]
  wire  andMatrixInput_9 = invInputs[26]; // @[pla.scala 90:29]
  wire  andMatrixInput_10 = invInputs[27]; // @[pla.scala 90:29]
  wire  andMatrixInput_11 = invInputs[28]; // @[pla.scala 90:29]
  wire  andMatrixInput_12 = invInputs[29]; // @[pla.scala 90:29]
  wire  andMatrixInput_13 = invInputs[31]; // @[pla.scala 90:29]
  wire [6:0] lo_1 = {andMatrixInput_3,andMatrixInput_8,andMatrixInput_9,andMatrixInput_10,andMatrixInput_11,
    andMatrixInput_12,andMatrixInput_13}; // @[Cat.scala 30:58]
  wire [13:0] _T_9 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_3_1,andMatrixInput_4,
    andMatrixInput_2,andMatrixInput_6,lo_1}; // @[Cat.scala 30:58]
  wire  _T_10 = &_T_9; // @[pla.scala 97:74]
  wire  andMatrixInput_5_1 = io_in__inst[12]; // @[pla.scala 89:45]
  wire  andMatrixInput_7_1 = io_in__inst[14]; // @[pla.scala 89:45]
  wire [6:0] lo_2 = {andMatrixInput_7_1,andMatrixInput_8,andMatrixInput_9,andMatrixInput_10,andMatrixInput_11,
    andMatrixInput_12,andMatrixInput_13}; // @[Cat.scala 30:58]
  wire [13:0] _T_11 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_3_1,andMatrixInput_4,
    andMatrixInput_5_1,andMatrixInput_6,lo_2}; // @[Cat.scala 30:58]
  wire  _T_12 = &_T_11; // @[pla.scala 97:74]
  wire  andMatrixInput_3_3 = invInputs[30]; // @[pla.scala 90:29]
  wire [3:0] _T_13 = {andMatrixInput_3_1,andMatrixInput_2,andMatrixInput_3,andMatrixInput_3_3}; // @[Cat.scala 30:58]
  wire  _T_14 = &_T_13; // @[pla.scala 97:74]
  wire  andMatrixInput_3_4 = io_in__inst[3]; // @[pla.scala 89:45]
  wire [6:0] lo_4 = {andMatrixInput_8,andMatrixInput_9,andMatrixInput_10,andMatrixInput_11,andMatrixInput_12,
    andMatrixInput_3_3,andMatrixInput_13}; // @[Cat.scala 30:58]
  wire [1:0] hi_hi_lo_2 = {andMatrixInput_0_1,andMatrixInput_3_4}; // @[Cat.scala 30:58]
  wire [14:0] _T_15 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_3_4,andMatrixInput_3_1,
    andMatrixInput_4,andMatrixInput_5_1,andMatrixInput_6,lo_4}; // @[Cat.scala 30:58]
  wire  _T_16 = &_T_15; // @[pla.scala 97:74]
  wire  andMatrixInput_0_6 = invInputs[5]; // @[pla.scala 90:29]
  wire  _T_17 = &andMatrixInput_0_6; // @[pla.scala 97:74]
  wire  andMatrixInput_5_3 = io_in__inst[5]; // @[pla.scala 89:45]
  wire [7:0] _T_18 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_0,andMatrixInput_3_1,
    andMatrixInput_5_3,andMatrixInput_1,andMatrixInput_2_1}; // @[Cat.scala 30:58]
  wire  _T_19 = &_T_18; // @[pla.scala 97:74]
  wire  andMatrixInput_4_4 = invInputs[4]; // @[pla.scala 90:29]
  wire [7:0] _T_20 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_0,andMatrixInput_4_4,
    andMatrixInput_0_6,andMatrixInput_4,andMatrixInput_3}; // @[Cat.scala 30:58]
  wire  _T_21 = &_T_20; // @[pla.scala 97:74]
  wire  andMatrixInput_2_8 = invInputs[20]; // @[pla.scala 90:29]
  wire [2:0] _T_22 = {andMatrixInput_0,andMatrixInput_1,andMatrixInput_2_8}; // @[Cat.scala 30:58]
  wire  _T_23 = &_T_22; // @[pla.scala 97:74]
  wire  andMatrixInput_7_5 = invInputs[7]; // @[pla.scala 90:29]
  wire  andMatrixInput_8_3 = invInputs[8]; // @[pla.scala 90:29]
  wire  andMatrixInput_9_3 = invInputs[9]; // @[pla.scala 90:29]
  wire  andMatrixInput_10_3 = invInputs[10]; // @[pla.scala 90:29]
  wire  andMatrixInput_11_3 = invInputs[11]; // @[pla.scala 90:29]
  wire  andMatrixInput_13_3 = invInputs[15]; // @[pla.scala 90:29]
  wire  andMatrixInput_14_1 = invInputs[16]; // @[pla.scala 90:29]
  wire  andMatrixInput_15 = invInputs[17]; // @[pla.scala 90:29]
  wire  andMatrixInput_16 = invInputs[18]; // @[pla.scala 90:29]
  wire  andMatrixInput_17 = invInputs[19]; // @[pla.scala 90:29]
  wire  andMatrixInput_18 = io_in__inst[20]; // @[pla.scala 89:45]
  wire  andMatrixInput_19 = invInputs[21]; // @[pla.scala 90:29]
  wire  andMatrixInput_20 = io_in__inst[22]; // @[pla.scala 89:45]
  wire  andMatrixInput_21 = invInputs[23]; // @[pla.scala 90:29]
  wire  andMatrixInput_22 = invInputs[24]; // @[pla.scala 90:29]
  wire  andMatrixInput_26 = io_in__inst[28]; // @[pla.scala 89:45]
  wire [6:0] lo_lo_5 = {andMatrixInput_8,andMatrixInput_9,andMatrixInput_10,andMatrixInput_26,andMatrixInput_12,
    andMatrixInput_3_3,andMatrixInput_13}; // @[Cat.scala 30:58]
  wire [14:0] lo_7 = {andMatrixInput_15,andMatrixInput_16,andMatrixInput_17,andMatrixInput_18,andMatrixInput_19,
    andMatrixInput_20,andMatrixInput_21,andMatrixInput_22,lo_lo_5}; // @[Cat.scala 30:58]
  wire [6:0] hi_lo_5 = {andMatrixInput_8_3,andMatrixInput_9_3,andMatrixInput_10_3,andMatrixInput_11_3,andMatrixInput_3,
    andMatrixInput_13_3,andMatrixInput_14_1}; // @[Cat.scala 30:58]
  wire [29:0] _T_24 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_0,andMatrixInput_3_1,
    andMatrixInput_5_3,andMatrixInput_1,andMatrixInput_7_5,hi_lo_5,lo_7}; // @[Cat.scala 30:58]
  wire  _T_25 = &_T_24; // @[pla.scala 97:74]
  wire  andMatrixInput_2_10 = io_in__inst[2]; // @[pla.scala 89:45]
  wire [5:0] _T_26 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_2_10,andMatrixInput_0,andMatrixInput_3_1,
    andMatrixInput_4}; // @[Cat.scala 30:58]
  wire  _T_27 = &_T_26; // @[pla.scala 97:74]
  wire  andMatrixInput_19_1 = io_in__inst[21]; // @[pla.scala 89:45]
  wire  andMatrixInput_20_1 = invInputs[22]; // @[pla.scala 90:29]
  wire  andMatrixInput_27_1 = io_in__inst[29]; // @[pla.scala 89:45]
  wire [6:0] lo_lo_6 = {andMatrixInput_8,andMatrixInput_9,andMatrixInput_10,andMatrixInput_26,andMatrixInput_27_1,
    andMatrixInput_3_3,andMatrixInput_13}; // @[Cat.scala 30:58]
  wire [14:0] lo_9 = {andMatrixInput_15,andMatrixInput_16,andMatrixInput_17,andMatrixInput_2_8,andMatrixInput_19_1,
    andMatrixInput_20_1,andMatrixInput_21,andMatrixInput_22,lo_lo_6}; // @[Cat.scala 30:58]
  wire [29:0] _T_28 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_0,andMatrixInput_3_1,
    andMatrixInput_5_3,andMatrixInput_1,andMatrixInput_7_5,hi_lo_5,lo_9}; // @[Cat.scala 30:58]
  wire  _T_29 = &_T_28; // @[pla.scala 97:74]
  wire [5:0] lo_10 = {andMatrixInput_9,andMatrixInput_10,andMatrixInput_11,andMatrixInput_12,andMatrixInput_3_3,
    andMatrixInput_13}; // @[Cat.scala 30:58]
  wire [11:0] _T_30 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0,andMatrixInput_3_1,andMatrixInput_4,
    andMatrixInput_8,lo_10}; // @[Cat.scala 30:58]
  wire  _T_31 = &_T_30; // @[pla.scala 97:74]
  wire [6:0] _T_32 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_0,andMatrixInput_0_6,
    andMatrixInput_4,andMatrixInput_2}; // @[Cat.scala 30:58]
  wire  _T_33 = &_T_32; // @[pla.scala 97:74]
  wire [3:0] _T_34 = {andMatrixInput_0_1,andMatrixInput_5_3,andMatrixInput_5_1,andMatrixInput_2_1}; // @[Cat.scala 30:58]
  wire  _T_35 = &_T_34; // @[pla.scala 97:74]
  wire [9:0] _T_36 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_3_4,andMatrixInput_3_1,
    andMatrixInput_0_6,andMatrixInput_4,andMatrixInput_2,andMatrixInput_6,andMatrixInput_3}; // @[Cat.scala 30:58]
  wire  _T_37 = &_T_36; // @[pla.scala 97:74]
  wire [11:0] _T_38 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0,andMatrixInput_3_1,andMatrixInput_0_6,
    andMatrixInput_4,lo_10}; // @[Cat.scala 30:58]
  wire  _T_39 = &_T_38; // @[pla.scala 97:74]
  wire [3:0] _T_40 = {andMatrixInput_0_1,andMatrixInput_5_3,andMatrixInput_5_1,andMatrixInput_6}; // @[Cat.scala 30:58]
  wire  _T_41 = &_T_40; // @[pla.scala 97:74]
  wire [3:0] _T_42 = {andMatrixInput_0_1,andMatrixInput_5_3,andMatrixInput_2,andMatrixInput_2_1}; // @[Cat.scala 30:58]
  wire  _T_43 = &_T_42; // @[pla.scala 97:74]
  wire [4:0] _T_44 = {andMatrixInput_0_1,andMatrixInput_4_4,andMatrixInput_5_1,andMatrixInput_6,andMatrixInput_7_1}; // @[Cat.scala 30:58]
  wire  _T_45 = &_T_44; // @[pla.scala 97:74]
  wire [2:0] _T_46 = {andMatrixInput_0_1,andMatrixInput_2_1,andMatrixInput_7_1}; // @[Cat.scala 30:58]
  wire  _T_47 = &_T_46; // @[pla.scala 97:74]
  wire [9:0] _T_48 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_2_10,andMatrixInput_3_4,andMatrixInput_4_4,
    andMatrixInput_0_6,andMatrixInput_4,andMatrixInput_5_1,andMatrixInput_6,andMatrixInput_3}; // @[Cat.scala 30:58]
  wire  _T_49 = &_T_48; // @[pla.scala 97:74]
  wire [3:0] _T_50 = {andMatrixInput_4_4,andMatrixInput_0_6,andMatrixInput_6,andMatrixInput_3}; // @[Cat.scala 30:58]
  wire  _T_51 = &_T_50; // @[pla.scala 97:74]
  wire  andMatrixInput_2_23 = io_in__inst[30]; // @[pla.scala 89:45]
  wire [2:0] _T_52 = {andMatrixInput_0_1,andMatrixInput_5_3,andMatrixInput_2_23}; // @[Cat.scala 30:58]
  wire  _T_53 = &_T_52; // @[pla.scala 97:74]
  wire [3:0] _T_54 = {andMatrixInput_0_1,andMatrixInput_1,andMatrixInput_2_1,andMatrixInput_3}; // @[Cat.scala 30:58]
  wire  _T_55 = &_T_54; // @[pla.scala 97:74]
  wire [1:0] _T_56 = {andMatrixInput_6,andMatrixInput_19_1}; // @[Cat.scala 30:58]
  wire  _T_57 = &_T_56; // @[pla.scala 97:74]
  wire [2:0] _T_58 = {andMatrixInput_0_1,andMatrixInput_5_1,andMatrixInput_6}; // @[Cat.scala 30:58]
  wire  _T_59 = &_T_58; // @[pla.scala 97:74]
  wire [2:0] _T_60 = {andMatrixInput_0_1,andMatrixInput_3_1,andMatrixInput_4}; // @[Cat.scala 30:58]
  wire  _T_61 = &_T_60; // @[pla.scala 97:74]
  wire [7:0] _T_62 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_0,andMatrixInput_4_4,
    andMatrixInput_5_3,andMatrixInput_1,andMatrixInput_6}; // @[Cat.scala 30:58]
  wire  _T_63 = &_T_62; // @[pla.scala 97:74]
  wire [2:0] _T_64 = {andMatrixInput_0,andMatrixInput_4_4,andMatrixInput_1}; // @[Cat.scala 30:58]
  wire  _T_65 = &_T_64; // @[pla.scala 97:74]
  wire [2:0] _T_66 = {andMatrixInput_5_1,andMatrixInput_2_1,andMatrixInput_7_1}; // @[Cat.scala 30:58]
  wire  _T_67 = &_T_66; // @[pla.scala 97:74]
  wire  _T_69 = &hi_hi_lo_2; // @[pla.scala 97:74]
  wire [1:0] _T_70 = {andMatrixInput_2_10,andMatrixInput_0_6}; // @[Cat.scala 30:58]
  wire  _T_71 = &_T_70; // @[pla.scala 97:74]
  wire [14:0] _T_72 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_3_4,andMatrixInput_3_1,
    andMatrixInput_4,andMatrixInput_5_1,andMatrixInput_6,lo_2}; // @[Cat.scala 30:58]
  wire  _T_73 = &_T_72; // @[pla.scala 97:74]
  wire [14:0] _T_74 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_3_4,andMatrixInput_3_1,
    andMatrixInput_4,andMatrixInput_2,andMatrixInput_6,lo_1}; // @[Cat.scala 30:58]
  wire  _T_75 = &_T_74; // @[pla.scala 97:74]
  wire [5:0] lo_24 = {andMatrixInput_7_1,andMatrixInput_9,andMatrixInput_10,andMatrixInput_11,andMatrixInput_12,
    andMatrixInput_13}; // @[Cat.scala 30:58]
  wire [11:0] _T_76 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0,andMatrixInput_3_1,andMatrixInput_0_6,
    andMatrixInput_4,lo_24}; // @[Cat.scala 30:58]
  wire  _T_77 = &_T_76; // @[pla.scala 97:74]
  wire [3:0] _T_78 = {andMatrixInput_0_1,andMatrixInput_0_6,andMatrixInput_2,andMatrixInput_3}; // @[Cat.scala 30:58]
  wire  _T_79 = &_T_78; // @[pla.scala 97:74]
  wire [3:0] _T_80 = {andMatrixInput_3_1,andMatrixInput_1,andMatrixInput_5_1,andMatrixInput_3}; // @[Cat.scala 30:58]
  wire  _T_81 = &_T_80; // @[pla.scala 97:74]
  wire [6:0] _T_82 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_0,andMatrixInput_4_4,
    andMatrixInput_4,andMatrixInput_3}; // @[Cat.scala 30:58]
  wire  _T_83 = &_T_82; // @[pla.scala 97:74]
  wire [7:0] _T_84 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_0,andMatrixInput_4_4,
    andMatrixInput_0_6,andMatrixInput_4,andMatrixInput_6}; // @[Cat.scala 30:58]
  wire  _T_85 = &_T_84; // @[pla.scala 97:74]
  wire [3:0] _T_86 = {andMatrixInput_0_1,andMatrixInput_0_6,andMatrixInput_5_1,andMatrixInput_2_1}; // @[Cat.scala 30:58]
  wire  _T_87 = &_T_86; // @[pla.scala 97:74]
  wire [1:0] _T_88 = {andMatrixInput_2_10,andMatrixInput_3_4}; // @[Cat.scala 30:58]
  wire  _T_89 = &_T_88; // @[pla.scala 97:74]
  wire [14:0] lo_30 = {andMatrixInput_15,andMatrixInput_16,andMatrixInput_17,andMatrixInput_2_8,andMatrixInput_19,
    andMatrixInput_20_1,andMatrixInput_21,andMatrixInput_22,lo_4}; // @[Cat.scala 30:58]
  wire [6:0] hi_lo_18 = {andMatrixInput_10_3,andMatrixInput_11_3,andMatrixInput_2,andMatrixInput_6,andMatrixInput_3,
    andMatrixInput_13_3,andMatrixInput_14_1}; // @[Cat.scala 30:58]
  wire [29:0] _T_90 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_5_3,andMatrixInput_1,
    andMatrixInput_7_5,andMatrixInput_8_3,andMatrixInput_9_3,hi_lo_18,lo_30}; // @[Cat.scala 30:58]
  wire  _T_91 = &_T_90; // @[pla.scala 97:74]
  wire [7:0] _T_92 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_0,andMatrixInput_3_1,
    andMatrixInput_5_3,andMatrixInput_1,andMatrixInput_5_1}; // @[Cat.scala 30:58]
  wire  _T_93 = &_T_92; // @[pla.scala 97:74]
  wire [3:0] _T_94 = {andMatrixInput_0_1,andMatrixInput_5_1,andMatrixInput_6,andMatrixInput_2_23}; // @[Cat.scala 30:58]
  wire  _T_95 = &_T_94; // @[pla.scala 97:74]
  wire [6:0] _T_96 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0,andMatrixInput_3_1,andMatrixInput_0_6,
    andMatrixInput_4,andMatrixInput_2_1}; // @[Cat.scala 30:58]
  wire  _T_97 = &_T_96; // @[pla.scala 97:74]
  wire [4:0] _T_98 = {andMatrixInput_0_1,andMatrixInput_0,andMatrixInput_3_1,andMatrixInput_5_1,andMatrixInput_6}; // @[Cat.scala 30:58]
  wire  _T_99 = &_T_98; // @[pla.scala 97:74]
  wire [3:0] _T_100 = {andMatrixInput_0_1,andMatrixInput_5_3,andMatrixInput_2,andMatrixInput_6}; // @[Cat.scala 30:58]
  wire  _T_101 = &_T_100; // @[pla.scala 97:74]
  wire [2:0] _T_102 = {andMatrixInput_5_1,andMatrixInput_7_1,andMatrixInput_3_3}; // @[Cat.scala 30:58]
  wire  _T_103 = &_T_102; // @[pla.scala 97:74]
  wire [6:0] _T_104 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_2_10,andMatrixInput_3_4,andMatrixInput_4_4,
    andMatrixInput_5_3,andMatrixInput_1}; // @[Cat.scala 30:58]
  wire  _T_105 = &_T_104; // @[pla.scala 97:74]
  wire [2:0] _T_106 = {andMatrixInput_0_1,andMatrixInput_4_4,andMatrixInput_4}; // @[Cat.scala 30:58]
  wire  _T_107 = &_T_106; // @[pla.scala 97:74]
  wire [7:0] _T_108 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_0_1,andMatrixInput_0,andMatrixInput_4_4,
    andMatrixInput_5_3,andMatrixInput_1,andMatrixInput_7_1}; // @[Cat.scala 30:58]
  wire  _T_109 = &_T_108; // @[pla.scala 97:74]
  wire [2:0] _T_110 = {andMatrixInput_3_1,andMatrixInput_1,andMatrixInput_7_1}; // @[Cat.scala 30:58]
  wire  _T_111 = &_T_110; // @[pla.scala 97:74]
  wire [8:0] _T_112 = {andMatrixInput_0_2,andMatrixInput_1_2,andMatrixInput_2_10,andMatrixInput_4_4,andMatrixInput_5_3,
    andMatrixInput_1,andMatrixInput_2,andMatrixInput_6,andMatrixInput_3}; // @[Cat.scala 30:58]
  wire  _T_113 = &_T_112; // @[pla.scala 97:74]
  wire [3:0] _T_114 = {andMatrixInput_0_1,andMatrixInput_2,andMatrixInput_6,andMatrixInput_7_1}; // @[Cat.scala 30:58]
  wire  _T_115 = &_T_114; // @[pla.scala 97:74]
  wire [1:0] _T_116 = {andMatrixInput_2_10,andMatrixInput_3_1}; // @[Cat.scala 30:58]
  wire  _T_117 = &_T_116; // @[pla.scala 97:74]
  wire [9:0] _orMatrixOutputs_T = {_T_45,_T_47,_T_51,_T_65,_T_69,_T_79,_T_87,_T_89,_T_111,_T_115}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_1 = |_orMatrixOutputs_T; // @[pla.scala 113:41]
  wire [4:0] _orMatrixOutputs_T_2 = {_T_35,_T_41,_T_43,_T_99,_T_101}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_3 = |_orMatrixOutputs_T_2; // @[pla.scala 113:41]
  wire [3:0] _orMatrixOutputs_T_4 = {_T_89,_T_99,_T_111,_T_117}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_5 = |_orMatrixOutputs_T_4; // @[pla.scala 113:41]
  wire [7:0] orMatrixOutputs_lo_3 = {_T_37,_T_39,_T_77,_T_85,_T_93,_T_97,_T_105,_T_113}; // @[Cat.scala 30:58]
  wire [15:0] _orMatrixOutputs_T_6 = {_T_10,_T_12,_T_16,_T_19,_T_21,_T_27,_T_31,_T_33,orMatrixOutputs_lo_3}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_7 = |_orMatrixOutputs_T_6; // @[pla.scala 113:41]
  wire [4:0] _orMatrixOutputs_T_8 = {_T_6,_T_35,_T_41,_T_43,_T_101}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_9 = |_orMatrixOutputs_T_8; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_10 = {_T_17,_T_89,_T_117}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_11 = |_orMatrixOutputs_T_10; // @[pla.scala 113:41]
  wire [6:0] _orMatrixOutputs_T_12 = {_T_55,_T_61,_T_65,_T_71,_T_81,_T_89,_T_107}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_13 = |_orMatrixOutputs_T_12; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_14 = {_T_71,_T_89,_T_111}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_15 = |_orMatrixOutputs_T_14; // @[pla.scala 113:41]
  wire [3:0] _orMatrixOutputs_T_16 = {_T_16,_T_37,_T_73,_T_75}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_17 = |_orMatrixOutputs_T_16; // @[pla.scala 113:41]
  wire [3:0] _orMatrixOutputs_T_18 = {_T_35,_T_41,_T_57,_T_71}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_19 = |_orMatrixOutputs_T_18; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_20 = {_T_35,_T_43,_T_71}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_21 = |_orMatrixOutputs_T_20; // @[pla.scala 113:41]
  wire [1:0] _orMatrixOutputs_T_22 = {_T_71,_T_101}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_23 = |_orMatrixOutputs_T_22; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_24 = {_T_35,_T_59,_T_87}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_25 = |_orMatrixOutputs_T_24; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_26 = {_T_8,_T_35,_T_87}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_27 = |_orMatrixOutputs_T_26; // @[pla.scala 113:41]
  wire [5:0] _orMatrixOutputs_T_28 = {_T_35,_T_41,_T_43,_T_51,_T_79,_T_101}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_29 = |_orMatrixOutputs_T_28; // @[pla.scala 113:41]
  wire [7:0] _orMatrixOutputs_T_30 = {_T_35,_T_41,_T_43,_T_45,_T_47,_T_87,_T_101,_T_115}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_31 = |_orMatrixOutputs_T_30; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_32 = {_T_43,_T_89,_T_101}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_33 = |_orMatrixOutputs_T_32; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_34 = {_T_6,_T_43,_T_45}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_35 = |_orMatrixOutputs_T_34; // @[pla.scala 113:41]
  wire [2:0] _orMatrixOutputs_T_36 = {_T_41,_T_43,_T_115}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_37 = |_orMatrixOutputs_T_36; // @[pla.scala 113:41]
  wire  _orMatrixOutputs_T_38 = |_T_35; // @[pla.scala 113:41]
  wire [5:0] _orMatrixOutputs_T_39 = {_T_14,_T_67,_T_79,_T_103,_T_115,_T_117}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_40 = |_orMatrixOutputs_T_39; // @[pla.scala 113:41]
  wire [3:0] _orMatrixOutputs_T_41 = {_T_8,_T_47,_T_53,_T_95}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_42 = |_orMatrixOutputs_T_41; // @[pla.scala 113:41]
  wire [3:0] _orMatrixOutputs_T_43 = {_T_35,_T_47,_T_87,_T_115}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_44 = |_orMatrixOutputs_T_43; // @[pla.scala 113:41]
  wire  _orMatrixOutputs_T_45 = |_T_59; // @[pla.scala 113:41]
  wire [7:0] _orMatrixOutputs_T_46 = {_T_14,_T_55,_T_61,_T_69,_T_71,_T_81,_T_111,_T_117}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_47 = |_orMatrixOutputs_T_46; // @[pla.scala 113:41]
  wire [5:0] _orMatrixOutputs_T_48 = {_T_23,_T_55,_T_65,_T_81,_T_89,_T_111}; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_49 = |_orMatrixOutputs_T_48; // @[pla.scala 113:41]
  wire  _orMatrixOutputs_T_50 = |_T_107; // @[pla.scala 113:41]
  wire [4:0] orMatrixOutputs_lo_lo_4 = {_T_93,_T_97,_T_105,_T_109,_T_113}; // @[Cat.scala 30:58]
  wire [10:0] orMatrixOutputs_lo_15 = {_T_49,_T_63,_T_77,_T_83,_T_85,_T_91,orMatrixOutputs_lo_lo_4}; // @[Cat.scala 30:58]
  wire [4:0] orMatrixOutputs_hi_lo_5 = {_T_29,_T_31,_T_33,_T_37,_T_39}; // @[Cat.scala 30:58]
  wire [21:0] _orMatrixOutputs_T_51 = {_T_10,_T_12,_T_16,_T_19,_T_25,_T_27,orMatrixOutputs_hi_lo_5,orMatrixOutputs_lo_15
    }; // @[Cat.scala 30:58]
  wire  _orMatrixOutputs_T_52 = |_orMatrixOutputs_T_51; // @[pla.scala 113:41]
  wire [6:0] orMatrixOutputs_lo_lo_5 = {_orMatrixOutputs_T_13,_orMatrixOutputs_T_11,_orMatrixOutputs_T_9,
    _orMatrixOutputs_T_7,_orMatrixOutputs_T_5,_orMatrixOutputs_T_3,_orMatrixOutputs_T_1}; // @[Cat.scala 30:58]
  wire [13:0] orMatrixOutputs_lo_16 = {_orMatrixOutputs_T_27,_orMatrixOutputs_T_25,_orMatrixOutputs_T_23,
    _orMatrixOutputs_T_21,_orMatrixOutputs_T_19,_orMatrixOutputs_T_17,_orMatrixOutputs_T_15,orMatrixOutputs_lo_lo_5}; // @[Cat.scala 30:58]
  wire [6:0] orMatrixOutputs_hi_lo_6 = {_orMatrixOutputs_T_40,_orMatrixOutputs_T_38,_orMatrixOutputs_T_37,
    _orMatrixOutputs_T_35,_orMatrixOutputs_T_33,_orMatrixOutputs_T_31,_orMatrixOutputs_T_29}; // @[Cat.scala 30:58]
  wire [27:0] orMatrixOutputs = {_orMatrixOutputs_T_52,_orMatrixOutputs_T_50,_orMatrixOutputs_T_49,_orMatrixOutputs_T_47
    ,_orMatrixOutputs_T_45,_orMatrixOutputs_T_44,_orMatrixOutputs_T_42,orMatrixOutputs_hi_lo_6,orMatrixOutputs_lo_16}; // @[Cat.scala 30:58]
  wire [6:0] invMatrixOutputs_lo_lo = {orMatrixOutputs[6],orMatrixOutputs[5],orMatrixOutputs[4],orMatrixOutputs[3],
    orMatrixOutputs[2],orMatrixOutputs[1],orMatrixOutputs[0]}; // @[Cat.scala 30:58]
  wire [13:0] invMatrixOutputs_lo = {orMatrixOutputs[13],orMatrixOutputs[12],orMatrixOutputs[11],orMatrixOutputs[10],
    orMatrixOutputs[9],orMatrixOutputs[8],orMatrixOutputs[7],invMatrixOutputs_lo_lo}; // @[Cat.scala 30:58]
  wire [6:0] invMatrixOutputs_hi_lo = {orMatrixOutputs[20],orMatrixOutputs[19],orMatrixOutputs[18],orMatrixOutputs[17],
    orMatrixOutputs[16],orMatrixOutputs[15],orMatrixOutputs[14]}; // @[Cat.scala 30:58]
  wire [27:0] invMatrixOutputs = {orMatrixOutputs[27],orMatrixOutputs[26],orMatrixOutputs[25],orMatrixOutputs[24],
    orMatrixOutputs[23],orMatrixOutputs[22],orMatrixOutputs[21],invMatrixOutputs_hi_lo,invMatrixOutputs_lo}; // @[Cat.scala 30:58]
  wire [1:0] uop_rs2_src = invMatrixOutputs[5:4]; // @[MicroOp.scala 56:20]
  wire [1:0] uop_rs1_src = invMatrixOutputs[7:6]; // @[MicroOp.scala 56:20]
  wire  uop_w_type = invMatrixOutputs[8]; // @[MicroOp.scala 54:20]
  wire [2:0] uop_sys_code = invMatrixOutputs[11:9]; // @[MicroOp.scala 56:20]
  wire [1:0] uop_mem_size = invMatrixOutputs[13:12]; // @[MicroOp.scala 56:20]
  wire [1:0] uop_mem_code = invMatrixOutputs[15:14]; // @[MicroOp.scala 56:20]
  wire [3:0] uop_jmp_code = invMatrixOutputs[19:16]; // @[MicroOp.scala 56:20]
  wire [3:0] uop_alu_code = invMatrixOutputs[23:20]; // @[MicroOp.scala 56:20]
  wire [2:0] uop_fu_code = invMatrixOutputs[26:24]; // @[MicroOp.scala 56:20]
  wire  uop_valid = invMatrixOutputs[27]; // @[MicroOp.scala 54:20]
  wire  uop_rd_en = invMatrixOutputs[3] & uop_rd_addr != 5'h0; // @[MicroOp.scala 61:24]
  wire [20:0] _T_135 = io_in__inst[31] ? 21'h1fffff : 21'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_137 = {_T_135,io_in__inst[30:20]}; // @[Cat.scala 30:58]
  wire [31:0] _T_143 = {_T_135,io_in__inst[30:25],uop_rd_addr}; // @[Cat.scala 30:58]
  wire [19:0] _T_146 = io_in__inst[31] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_150 = {_T_146,io_in__inst[7],io_in__inst[30:25],io_in__inst[11:8],1'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_153 = {io_in__inst[31:12],12'h0}; // @[Cat.scala 30:58]
  wire [11:0] _T_156 = io_in__inst[31] ? 12'hfff : 12'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_160 = {_T_156,io_in__inst[19:12],andMatrixInput_18,io_in__inst[30:21],1'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_163 = {27'h0,uop_rs2_addr}; // @[Cat.scala 30:58]
  wire [31:0] _T_166 = {26'h0,io_in__inst[25:20]}; // @[Cat.scala 30:58]
  wire [31:0] _T_167 = uop_w_type ? _T_163 : _T_166; // @[MicroOp.scala 68:24]
  wire [31:0] _T_170 = {27'h0,uop_rs1_addr}; // @[Cat.scala 30:58]
  wire [31:0] _T_172 = 3'h1 == invMatrixOutputs[2:0] ? _T_137 : 32'h0; // @[Mux.scala 80:57]
  wire [31:0] _T_174 = 3'h2 == invMatrixOutputs[2:0] ? _T_143 : _T_172; // @[Mux.scala 80:57]
  wire [31:0] _T_176 = 3'h3 == invMatrixOutputs[2:0] ? _T_150 : _T_174; // @[Mux.scala 80:57]
  wire [31:0] _T_178 = 3'h4 == invMatrixOutputs[2:0] ? _T_153 : _T_176; // @[Mux.scala 80:57]
  wire [31:0] _T_180 = 3'h5 == invMatrixOutputs[2:0] ? _T_160 : _T_178; // @[Mux.scala 80:57]
  wire [31:0] _T_182 = 3'h6 == invMatrixOutputs[2:0] ? _T_167 : _T_180; // @[Mux.scala 80:57]
  wire [31:0] uop_imm = 3'h7 == invMatrixOutputs[2:0] ? _T_170 : _T_182; // @[Mux.scala 80:57]
  assign io_out_valid = io_in_valid & io_in__valid & uop_valid; // @[Decode.scala 79:16]
  assign io_out_pc = io_in_valid & io_in__valid ? io_in__pc : 32'h0; // @[Decode.scala 79:16]
  assign io_out_npc = io_in_valid & io_in__valid ? uop_npc : 32'h0; // @[Decode.scala 79:16]
  assign io_out_inst = io_in_valid & io_in__valid ? io_in__inst : 32'h0; // @[Decode.scala 79:16]
  assign io_out_fu_code = io_in_valid & io_in__valid ? uop_fu_code : 3'h0; // @[Decode.scala 79:16]
  assign io_out_alu_code = io_in_valid & io_in__valid ? uop_alu_code : 4'h0; // @[Decode.scala 79:16]
  assign io_out_jmp_code = io_in_valid & io_in__valid ? uop_jmp_code : 4'h0; // @[Decode.scala 79:16]
  assign io_out_mem_code = io_in_valid & io_in__valid ? uop_mem_code : 2'h0; // @[Decode.scala 79:16]
  assign io_out_mem_size = io_in_valid & io_in__valid ? uop_mem_size : 2'h0; // @[Decode.scala 79:16]
  assign io_out_sys_code = io_in_valid & io_in__valid ? uop_sys_code : 3'h0; // @[Decode.scala 79:16]
  assign io_out_w_type = io_in_valid & io_in__valid & uop_w_type; // @[Decode.scala 79:16]
  assign io_out_rs1_src = io_in_valid & io_in__valid ? uop_rs1_src : 2'h0; // @[Decode.scala 79:16]
  assign io_out_rs2_src = io_in_valid & io_in__valid ? uop_rs2_src : 2'h0; // @[Decode.scala 79:16]
  assign io_out_rs1_addr = io_in_valid & io_in__valid ? uop_rs1_addr : 5'h0; // @[Decode.scala 79:16]
  assign io_out_rs2_addr = io_in_valid & io_in__valid ? uop_rs2_addr : 5'h0; // @[Decode.scala 79:16]
  assign io_out_rd_addr = io_in_valid & io_in__valid ? uop_rd_addr : 5'h0; // @[Decode.scala 79:16]
  assign io_out_rd_en = io_in_valid & io_in__valid & uop_rd_en; // @[Decode.scala 79:16]
  assign io_out_imm = io_in_valid & io_in__valid ? uop_imm : 32'h0; // @[Decode.scala 79:16]
  assign io_out_pred_br = io_in_valid & io_in__valid & io_in__pred_br; // @[Decode.scala 79:16]
  assign io_out_pred_bpc = io_in_valid & io_in__valid ? io_in__pred_bpc : 32'h0; // @[Decode.scala 79:16]
endmodule
module ysyx_210128_Decode(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_vec_0_pc,
  input  [31:0] io_in_bits_vec_0_inst,
  input         io_in_bits_vec_0_pred_br,
  input  [31:0] io_in_bits_vec_0_pred_bpc,
  input         io_in_bits_vec_0_valid,
  input  [31:0] io_in_bits_vec_1_pc,
  input  [31:0] io_in_bits_vec_1_inst,
  input         io_in_bits_vec_1_pred_br,
  input  [31:0] io_in_bits_vec_1_pred_bpc,
  input         io_in_bits_vec_1_valid,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_vec_0_valid,
  output [31:0] io_out_bits_vec_0_pc,
  output [31:0] io_out_bits_vec_0_npc,
  output [31:0] io_out_bits_vec_0_inst,
  output [2:0]  io_out_bits_vec_0_fu_code,
  output [3:0]  io_out_bits_vec_0_alu_code,
  output [3:0]  io_out_bits_vec_0_jmp_code,
  output [1:0]  io_out_bits_vec_0_mem_code,
  output [1:0]  io_out_bits_vec_0_mem_size,
  output [2:0]  io_out_bits_vec_0_sys_code,
  output        io_out_bits_vec_0_w_type,
  output [1:0]  io_out_bits_vec_0_rs1_src,
  output [1:0]  io_out_bits_vec_0_rs2_src,
  output [4:0]  io_out_bits_vec_0_rs1_addr,
  output [4:0]  io_out_bits_vec_0_rs2_addr,
  output [4:0]  io_out_bits_vec_0_rd_addr,
  output        io_out_bits_vec_0_rd_en,
  output [31:0] io_out_bits_vec_0_imm,
  output        io_out_bits_vec_0_pred_br,
  output [31:0] io_out_bits_vec_0_pred_bpc,
  output        io_out_bits_vec_1_valid,
  output [31:0] io_out_bits_vec_1_pc,
  output [31:0] io_out_bits_vec_1_npc,
  output [31:0] io_out_bits_vec_1_inst,
  output [2:0]  io_out_bits_vec_1_fu_code,
  output [3:0]  io_out_bits_vec_1_alu_code,
  output [3:0]  io_out_bits_vec_1_jmp_code,
  output [1:0]  io_out_bits_vec_1_mem_code,
  output [1:0]  io_out_bits_vec_1_mem_size,
  output [2:0]  io_out_bits_vec_1_sys_code,
  output        io_out_bits_vec_1_w_type,
  output [1:0]  io_out_bits_vec_1_rs1_src,
  output [1:0]  io_out_bits_vec_1_rs2_src,
  output [4:0]  io_out_bits_vec_1_rs1_addr,
  output [4:0]  io_out_bits_vec_1_rs2_addr,
  output [4:0]  io_out_bits_vec_1_rd_addr,
  output        io_out_bits_vec_1_rd_en,
  output [31:0] io_out_bits_vec_1_imm,
  output        io_out_bits_vec_1_pred_br,
  output [31:0] io_out_bits_vec_1_pred_bpc,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] decoder_0_io_in__pc; // @[Decode.scala 27:25]
  wire [31:0] decoder_0_io_in__inst; // @[Decode.scala 27:25]
  wire  decoder_0_io_in__pred_br; // @[Decode.scala 27:25]
  wire [31:0] decoder_0_io_in__pred_bpc; // @[Decode.scala 27:25]
  wire  decoder_0_io_in__valid; // @[Decode.scala 27:25]
  wire  decoder_0_io_in_valid; // @[Decode.scala 27:25]
  wire  decoder_0_io_out_valid; // @[Decode.scala 27:25]
  wire [31:0] decoder_0_io_out_pc; // @[Decode.scala 27:25]
  wire [31:0] decoder_0_io_out_npc; // @[Decode.scala 27:25]
  wire [31:0] decoder_0_io_out_inst; // @[Decode.scala 27:25]
  wire [2:0] decoder_0_io_out_fu_code; // @[Decode.scala 27:25]
  wire [3:0] decoder_0_io_out_alu_code; // @[Decode.scala 27:25]
  wire [3:0] decoder_0_io_out_jmp_code; // @[Decode.scala 27:25]
  wire [1:0] decoder_0_io_out_mem_code; // @[Decode.scala 27:25]
  wire [1:0] decoder_0_io_out_mem_size; // @[Decode.scala 27:25]
  wire [2:0] decoder_0_io_out_sys_code; // @[Decode.scala 27:25]
  wire  decoder_0_io_out_w_type; // @[Decode.scala 27:25]
  wire [1:0] decoder_0_io_out_rs1_src; // @[Decode.scala 27:25]
  wire [1:0] decoder_0_io_out_rs2_src; // @[Decode.scala 27:25]
  wire [4:0] decoder_0_io_out_rs1_addr; // @[Decode.scala 27:25]
  wire [4:0] decoder_0_io_out_rs2_addr; // @[Decode.scala 27:25]
  wire [4:0] decoder_0_io_out_rd_addr; // @[Decode.scala 27:25]
  wire  decoder_0_io_out_rd_en; // @[Decode.scala 27:25]
  wire [31:0] decoder_0_io_out_imm; // @[Decode.scala 27:25]
  wire  decoder_0_io_out_pred_br; // @[Decode.scala 27:25]
  wire [31:0] decoder_0_io_out_pred_bpc; // @[Decode.scala 27:25]
  wire [31:0] decoder_1_io_in__pc; // @[Decode.scala 27:25]
  wire [31:0] decoder_1_io_in__inst; // @[Decode.scala 27:25]
  wire  decoder_1_io_in__pred_br; // @[Decode.scala 27:25]
  wire [31:0] decoder_1_io_in__pred_bpc; // @[Decode.scala 27:25]
  wire  decoder_1_io_in__valid; // @[Decode.scala 27:25]
  wire  decoder_1_io_in_valid; // @[Decode.scala 27:25]
  wire  decoder_1_io_out_valid; // @[Decode.scala 27:25]
  wire [31:0] decoder_1_io_out_pc; // @[Decode.scala 27:25]
  wire [31:0] decoder_1_io_out_npc; // @[Decode.scala 27:25]
  wire [31:0] decoder_1_io_out_inst; // @[Decode.scala 27:25]
  wire [2:0] decoder_1_io_out_fu_code; // @[Decode.scala 27:25]
  wire [3:0] decoder_1_io_out_alu_code; // @[Decode.scala 27:25]
  wire [3:0] decoder_1_io_out_jmp_code; // @[Decode.scala 27:25]
  wire [1:0] decoder_1_io_out_mem_code; // @[Decode.scala 27:25]
  wire [1:0] decoder_1_io_out_mem_size; // @[Decode.scala 27:25]
  wire [2:0] decoder_1_io_out_sys_code; // @[Decode.scala 27:25]
  wire  decoder_1_io_out_w_type; // @[Decode.scala 27:25]
  wire [1:0] decoder_1_io_out_rs1_src; // @[Decode.scala 27:25]
  wire [1:0] decoder_1_io_out_rs2_src; // @[Decode.scala 27:25]
  wire [4:0] decoder_1_io_out_rs1_addr; // @[Decode.scala 27:25]
  wire [4:0] decoder_1_io_out_rs2_addr; // @[Decode.scala 27:25]
  wire [4:0] decoder_1_io_out_rd_addr; // @[Decode.scala 27:25]
  wire  decoder_1_io_out_rd_en; // @[Decode.scala 27:25]
  wire [31:0] decoder_1_io_out_imm; // @[Decode.scala 27:25]
  wire  decoder_1_io_out_pred_br; // @[Decode.scala 27:25]
  wire [31:0] decoder_1_io_out_pred_bpc; // @[Decode.scala 27:25]
  reg [31:0] reg_in_0_pc; // @[Decode.scala 16:23]
  reg [31:0] reg_in_0_inst; // @[Decode.scala 16:23]
  reg  reg_in_0_pred_br; // @[Decode.scala 16:23]
  reg [31:0] reg_in_0_pred_bpc; // @[Decode.scala 16:23]
  reg  reg_in_0_valid; // @[Decode.scala 16:23]
  reg [31:0] reg_in_1_pc; // @[Decode.scala 16:23]
  reg [31:0] reg_in_1_inst; // @[Decode.scala 16:23]
  reg  reg_in_1_pred_br; // @[Decode.scala 16:23]
  reg [31:0] reg_in_1_pred_bpc; // @[Decode.scala 16:23]
  reg  reg_in_1_valid; // @[Decode.scala 16:23]
  reg  reg_in_valid; // @[Decode.scala 17:29]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_10 = io_in_valid & ~io_flush & ~io_out_ready | reg_in_valid; // @[Decode.scala 21:59 23:18 17:29]
  reg  REG; // @[Decode.scala 39:32]
  ysyx_210128_Decoder decoder_0 ( // @[Decode.scala 27:25]
    .io_in__pc(decoder_0_io_in__pc),
    .io_in__inst(decoder_0_io_in__inst),
    .io_in__pred_br(decoder_0_io_in__pred_br),
    .io_in__pred_bpc(decoder_0_io_in__pred_bpc),
    .io_in__valid(decoder_0_io_in__valid),
    .io_in_valid(decoder_0_io_in_valid),
    .io_out_valid(decoder_0_io_out_valid),
    .io_out_pc(decoder_0_io_out_pc),
    .io_out_npc(decoder_0_io_out_npc),
    .io_out_inst(decoder_0_io_out_inst),
    .io_out_fu_code(decoder_0_io_out_fu_code),
    .io_out_alu_code(decoder_0_io_out_alu_code),
    .io_out_jmp_code(decoder_0_io_out_jmp_code),
    .io_out_mem_code(decoder_0_io_out_mem_code),
    .io_out_mem_size(decoder_0_io_out_mem_size),
    .io_out_sys_code(decoder_0_io_out_sys_code),
    .io_out_w_type(decoder_0_io_out_w_type),
    .io_out_rs1_src(decoder_0_io_out_rs1_src),
    .io_out_rs2_src(decoder_0_io_out_rs2_src),
    .io_out_rs1_addr(decoder_0_io_out_rs1_addr),
    .io_out_rs2_addr(decoder_0_io_out_rs2_addr),
    .io_out_rd_addr(decoder_0_io_out_rd_addr),
    .io_out_rd_en(decoder_0_io_out_rd_en),
    .io_out_imm(decoder_0_io_out_imm),
    .io_out_pred_br(decoder_0_io_out_pred_br),
    .io_out_pred_bpc(decoder_0_io_out_pred_bpc)
  );
  ysyx_210128_Decoder_1 decoder_1 ( // @[Decode.scala 27:25]
    .io_in__pc(decoder_1_io_in__pc),
    .io_in__inst(decoder_1_io_in__inst),
    .io_in__pred_br(decoder_1_io_in__pred_br),
    .io_in__pred_bpc(decoder_1_io_in__pred_bpc),
    .io_in__valid(decoder_1_io_in__valid),
    .io_in_valid(decoder_1_io_in_valid),
    .io_out_valid(decoder_1_io_out_valid),
    .io_out_pc(decoder_1_io_out_pc),
    .io_out_npc(decoder_1_io_out_npc),
    .io_out_inst(decoder_1_io_out_inst),
    .io_out_fu_code(decoder_1_io_out_fu_code),
    .io_out_alu_code(decoder_1_io_out_alu_code),
    .io_out_jmp_code(decoder_1_io_out_jmp_code),
    .io_out_mem_code(decoder_1_io_out_mem_code),
    .io_out_mem_size(decoder_1_io_out_mem_size),
    .io_out_sys_code(decoder_1_io_out_sys_code),
    .io_out_w_type(decoder_1_io_out_w_type),
    .io_out_rs1_src(decoder_1_io_out_rs1_src),
    .io_out_rs2_src(decoder_1_io_out_rs2_src),
    .io_out_rs1_addr(decoder_1_io_out_rs1_addr),
    .io_out_rs2_addr(decoder_1_io_out_rs2_addr),
    .io_out_rd_addr(decoder_1_io_out_rd_addr),
    .io_out_rd_en(decoder_1_io_out_rd_en),
    .io_out_imm(decoder_1_io_out_imm),
    .io_out_pred_br(decoder_1_io_out_pred_br),
    .io_out_pred_bpc(decoder_1_io_out_pred_bpc)
  );
  assign io_in_ready = io_out_ready; // @[Decode.scala 37:15]
  assign io_out_valid = io_out_ready & REG & ~io_in_valid ? reg_in_valid : io_in_valid; // @[Decode.scala 39:65 40:18 43:18]
  assign io_out_bits_vec_0_valid = _T & decoder_0_io_out_valid; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_pc = _T ? decoder_0_io_out_pc : 32'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_npc = _T ? decoder_0_io_out_npc : 32'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_inst = _T ? decoder_0_io_out_inst : 32'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_fu_code = _T ? decoder_0_io_out_fu_code : 3'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_alu_code = _T ? decoder_0_io_out_alu_code : 4'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_jmp_code = _T ? decoder_0_io_out_jmp_code : 4'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_mem_code = _T ? decoder_0_io_out_mem_code : 2'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_mem_size = _T ? decoder_0_io_out_mem_size : 2'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_sys_code = _T ? decoder_0_io_out_sys_code : 3'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_w_type = _T & decoder_0_io_out_w_type; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_rs1_src = _T ? decoder_0_io_out_rs1_src : 2'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_rs2_src = _T ? decoder_0_io_out_rs2_src : 2'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_rs1_addr = _T ? decoder_0_io_out_rs1_addr : 5'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_rs2_addr = _T ? decoder_0_io_out_rs2_addr : 5'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_rd_addr = _T ? decoder_0_io_out_rd_addr : 5'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_rd_en = _T & decoder_0_io_out_rd_en; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_imm = _T ? decoder_0_io_out_imm : 32'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_pred_br = _T & decoder_0_io_out_pred_br; // @[Decode.scala 47:30]
  assign io_out_bits_vec_0_pred_bpc = _T ? decoder_0_io_out_pred_bpc : 32'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_valid = _T & decoder_1_io_out_valid; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_pc = _T ? decoder_1_io_out_pc : 32'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_npc = _T ? decoder_1_io_out_npc : 32'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_inst = _T ? decoder_1_io_out_inst : 32'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_fu_code = _T ? decoder_1_io_out_fu_code : 3'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_alu_code = _T ? decoder_1_io_out_alu_code : 4'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_jmp_code = _T ? decoder_1_io_out_jmp_code : 4'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_mem_code = _T ? decoder_1_io_out_mem_code : 2'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_mem_size = _T ? decoder_1_io_out_mem_size : 2'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_sys_code = _T ? decoder_1_io_out_sys_code : 3'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_w_type = _T & decoder_1_io_out_w_type; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_rs1_src = _T ? decoder_1_io_out_rs1_src : 2'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_rs2_src = _T ? decoder_1_io_out_rs2_src : 2'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_rs1_addr = _T ? decoder_1_io_out_rs1_addr : 5'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_rs2_addr = _T ? decoder_1_io_out_rs2_addr : 5'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_rd_addr = _T ? decoder_1_io_out_rd_addr : 5'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_rd_en = _T & decoder_1_io_out_rd_en; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_imm = _T ? decoder_1_io_out_imm : 32'h0; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_pred_br = _T & decoder_1_io_out_pred_br; // @[Decode.scala 47:30]
  assign io_out_bits_vec_1_pred_bpc = _T ? decoder_1_io_out_pred_bpc : 32'h0; // @[Decode.scala 47:30]
  assign decoder_0_io_in__pc = io_in_valid ? io_in_bits_vec_0_pc : reg_in_0_pc; // @[Decode.scala 32:28]
  assign decoder_0_io_in__inst = io_in_valid ? io_in_bits_vec_0_inst : reg_in_0_inst; // @[Decode.scala 32:28]
  assign decoder_0_io_in__pred_br = io_in_valid ? io_in_bits_vec_0_pred_br : reg_in_0_pred_br; // @[Decode.scala 32:28]
  assign decoder_0_io_in__pred_bpc = io_in_valid ? io_in_bits_vec_0_pred_bpc : reg_in_0_pred_bpc; // @[Decode.scala 32:28]
  assign decoder_0_io_in__valid = io_in_valid ? io_in_bits_vec_0_valid : reg_in_0_valid; // @[Decode.scala 32:28]
  assign decoder_0_io_in_valid = io_in_valid | reg_in_valid; // @[Decode.scala 33:43]
  assign decoder_1_io_in__pc = io_in_valid ? io_in_bits_vec_1_pc : reg_in_1_pc; // @[Decode.scala 32:28]
  assign decoder_1_io_in__inst = io_in_valid ? io_in_bits_vec_1_inst : reg_in_1_inst; // @[Decode.scala 32:28]
  assign decoder_1_io_in__pred_br = io_in_valid ? io_in_bits_vec_1_pred_br : reg_in_1_pred_br; // @[Decode.scala 32:28]
  assign decoder_1_io_in__pred_bpc = io_in_valid ? io_in_bits_vec_1_pred_bpc : reg_in_1_pred_bpc; // @[Decode.scala 32:28]
  assign decoder_1_io_in__valid = io_in_valid ? io_in_bits_vec_1_valid : reg_in_1_valid; // @[Decode.scala 32:28]
  assign decoder_1_io_in_valid = io_in_valid | reg_in_valid; // @[Decode.scala 33:43]
  always @(posedge clock) begin
    if (reset) begin // @[Decode.scala 16:23]
      reg_in_0_pc <= 32'h0; // @[Decode.scala 16:23]
    end else if (!(io_flush | _T)) begin // @[Decode.scala 19:36]
      if (io_in_valid & ~io_flush & ~io_out_ready) begin // @[Decode.scala 21:59]
        reg_in_0_pc <= io_in_bits_vec_0_pc; // @[Decode.scala 22:12]
      end
    end
    if (reset) begin // @[Decode.scala 16:23]
      reg_in_0_inst <= 32'h0; // @[Decode.scala 16:23]
    end else if (!(io_flush | _T)) begin // @[Decode.scala 19:36]
      if (io_in_valid & ~io_flush & ~io_out_ready) begin // @[Decode.scala 21:59]
        reg_in_0_inst <= io_in_bits_vec_0_inst; // @[Decode.scala 22:12]
      end
    end
    if (reset) begin // @[Decode.scala 16:23]
      reg_in_0_pred_br <= 1'h0; // @[Decode.scala 16:23]
    end else if (!(io_flush | _T)) begin // @[Decode.scala 19:36]
      if (io_in_valid & ~io_flush & ~io_out_ready) begin // @[Decode.scala 21:59]
        reg_in_0_pred_br <= io_in_bits_vec_0_pred_br; // @[Decode.scala 22:12]
      end
    end
    if (reset) begin // @[Decode.scala 16:23]
      reg_in_0_pred_bpc <= 32'h0; // @[Decode.scala 16:23]
    end else if (!(io_flush | _T)) begin // @[Decode.scala 19:36]
      if (io_in_valid & ~io_flush & ~io_out_ready) begin // @[Decode.scala 21:59]
        reg_in_0_pred_bpc <= io_in_bits_vec_0_pred_bpc; // @[Decode.scala 22:12]
      end
    end
    if (reset) begin // @[Decode.scala 16:23]
      reg_in_0_valid <= 1'h0; // @[Decode.scala 16:23]
    end else if (!(io_flush | _T)) begin // @[Decode.scala 19:36]
      if (io_in_valid & ~io_flush & ~io_out_ready) begin // @[Decode.scala 21:59]
        reg_in_0_valid <= io_in_bits_vec_0_valid; // @[Decode.scala 22:12]
      end
    end
    if (reset) begin // @[Decode.scala 16:23]
      reg_in_1_pc <= 32'h0; // @[Decode.scala 16:23]
    end else if (!(io_flush | _T)) begin // @[Decode.scala 19:36]
      if (io_in_valid & ~io_flush & ~io_out_ready) begin // @[Decode.scala 21:59]
        reg_in_1_pc <= io_in_bits_vec_1_pc; // @[Decode.scala 22:12]
      end
    end
    if (reset) begin // @[Decode.scala 16:23]
      reg_in_1_inst <= 32'h0; // @[Decode.scala 16:23]
    end else if (!(io_flush | _T)) begin // @[Decode.scala 19:36]
      if (io_in_valid & ~io_flush & ~io_out_ready) begin // @[Decode.scala 21:59]
        reg_in_1_inst <= io_in_bits_vec_1_inst; // @[Decode.scala 22:12]
      end
    end
    if (reset) begin // @[Decode.scala 16:23]
      reg_in_1_pred_br <= 1'h0; // @[Decode.scala 16:23]
    end else if (!(io_flush | _T)) begin // @[Decode.scala 19:36]
      if (io_in_valid & ~io_flush & ~io_out_ready) begin // @[Decode.scala 21:59]
        reg_in_1_pred_br <= io_in_bits_vec_1_pred_br; // @[Decode.scala 22:12]
      end
    end
    if (reset) begin // @[Decode.scala 16:23]
      reg_in_1_pred_bpc <= 32'h0; // @[Decode.scala 16:23]
    end else if (!(io_flush | _T)) begin // @[Decode.scala 19:36]
      if (io_in_valid & ~io_flush & ~io_out_ready) begin // @[Decode.scala 21:59]
        reg_in_1_pred_bpc <= io_in_bits_vec_1_pred_bpc; // @[Decode.scala 22:12]
      end
    end
    if (reset) begin // @[Decode.scala 16:23]
      reg_in_1_valid <= 1'h0; // @[Decode.scala 16:23]
    end else if (!(io_flush | _T)) begin // @[Decode.scala 19:36]
      if (io_in_valid & ~io_flush & ~io_out_ready) begin // @[Decode.scala 21:59]
        reg_in_1_valid <= io_in_bits_vec_1_valid; // @[Decode.scala 22:12]
      end
    end
    if (reset) begin // @[Decode.scala 17:29]
      reg_in_valid <= 1'h0; // @[Decode.scala 17:29]
    end else if (io_out_ready & REG & ~io_in_valid) begin // @[Decode.scala 39:65]
      reg_in_valid <= 1'h0; // @[Decode.scala 41:18]
    end else if (io_flush | _T) begin // @[Decode.scala 19:36]
      reg_in_valid <= 1'h0; // @[Decode.scala 20:18]
    end else begin
      reg_in_valid <= _GEN_10;
    end
    REG <= ~io_out_ready; // @[Decode.scala 39:33]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_in_0_pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_in_0_inst = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_in_0_pred_br = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  reg_in_0_pred_bpc = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_in_0_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  reg_in_1_pc = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_in_1_inst = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_in_1_pred_br = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  reg_in_1_pred_bpc = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_in_1_valid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  reg_in_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_PrfStateTable(
  input         clock,
  input         reset,
  input         io_en,
  output        io_allocatable,
  input         io_rd_req_0,
  input         io_rd_req_1,
  output [5:0]  io_rd_paddr_0,
  output [5:0]  io_rd_paddr_1,
  input  [5:0]  io_exe_0,
  input  [5:0]  io_exe_1,
  input  [5:0]  io_exe_2,
  input  [5:0]  io_cm_0,
  input  [5:0]  io_cm_1,
  input  [5:0]  io_free_0,
  input  [5:0]  io_free_1,
  input         io_cm_recover,
  output [63:0] io_avail_list
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] table_1; // @[Rename.scala 186:22]
  reg [1:0] table_2; // @[Rename.scala 186:22]
  reg [1:0] table_3; // @[Rename.scala 186:22]
  reg [1:0] table_4; // @[Rename.scala 186:22]
  reg [1:0] table_5; // @[Rename.scala 186:22]
  reg [1:0] table_6; // @[Rename.scala 186:22]
  reg [1:0] table_7; // @[Rename.scala 186:22]
  reg [1:0] table_8; // @[Rename.scala 186:22]
  reg [1:0] table_9; // @[Rename.scala 186:22]
  reg [1:0] table_10; // @[Rename.scala 186:22]
  reg [1:0] table_11; // @[Rename.scala 186:22]
  reg [1:0] table_12; // @[Rename.scala 186:22]
  reg [1:0] table_13; // @[Rename.scala 186:22]
  reg [1:0] table_14; // @[Rename.scala 186:22]
  reg [1:0] table_15; // @[Rename.scala 186:22]
  reg [1:0] table_16; // @[Rename.scala 186:22]
  reg [1:0] table_17; // @[Rename.scala 186:22]
  reg [1:0] table_18; // @[Rename.scala 186:22]
  reg [1:0] table_19; // @[Rename.scala 186:22]
  reg [1:0] table_20; // @[Rename.scala 186:22]
  reg [1:0] table_21; // @[Rename.scala 186:22]
  reg [1:0] table_22; // @[Rename.scala 186:22]
  reg [1:0] table_23; // @[Rename.scala 186:22]
  reg [1:0] table_24; // @[Rename.scala 186:22]
  reg [1:0] table_25; // @[Rename.scala 186:22]
  reg [1:0] table_26; // @[Rename.scala 186:22]
  reg [1:0] table_27; // @[Rename.scala 186:22]
  reg [1:0] table_28; // @[Rename.scala 186:22]
  reg [1:0] table_29; // @[Rename.scala 186:22]
  reg [1:0] table_30; // @[Rename.scala 186:22]
  reg [1:0] table_31; // @[Rename.scala 186:22]
  reg [1:0] table_32; // @[Rename.scala 186:22]
  reg [1:0] table_33; // @[Rename.scala 186:22]
  reg [1:0] table_34; // @[Rename.scala 186:22]
  reg [1:0] table_35; // @[Rename.scala 186:22]
  reg [1:0] table_36; // @[Rename.scala 186:22]
  reg [1:0] table_37; // @[Rename.scala 186:22]
  reg [1:0] table_38; // @[Rename.scala 186:22]
  reg [1:0] table_39; // @[Rename.scala 186:22]
  reg [1:0] table_40; // @[Rename.scala 186:22]
  reg [1:0] table_41; // @[Rename.scala 186:22]
  reg [1:0] table_42; // @[Rename.scala 186:22]
  reg [1:0] table_43; // @[Rename.scala 186:22]
  reg [1:0] table_44; // @[Rename.scala 186:22]
  reg [1:0] table_45; // @[Rename.scala 186:22]
  reg [1:0] table_46; // @[Rename.scala 186:22]
  reg [1:0] table_47; // @[Rename.scala 186:22]
  reg [1:0] table_48; // @[Rename.scala 186:22]
  reg [1:0] table_49; // @[Rename.scala 186:22]
  reg [1:0] table_50; // @[Rename.scala 186:22]
  reg [1:0] table_51; // @[Rename.scala 186:22]
  reg [1:0] table_52; // @[Rename.scala 186:22]
  reg [1:0] table_53; // @[Rename.scala 186:22]
  reg [1:0] table_54; // @[Rename.scala 186:22]
  reg [1:0] table_55; // @[Rename.scala 186:22]
  reg [1:0] table_56; // @[Rename.scala 186:22]
  reg [1:0] table_57; // @[Rename.scala 186:22]
  reg [1:0] table_58; // @[Rename.scala 186:22]
  reg [1:0] table_59; // @[Rename.scala 186:22]
  reg [1:0] table_60; // @[Rename.scala 186:22]
  reg [1:0] table_61; // @[Rename.scala 186:22]
  reg [1:0] table_62; // @[Rename.scala 186:22]
  reg [1:0] table_63; // @[Rename.scala 186:22]
  wire  _T_1 = table_1 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_2 = table_2 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_3 = table_3 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_4 = table_4 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_5 = table_5 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_6 = table_6 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_7 = table_7 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_8 = table_8 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_9 = table_9 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_10 = table_10 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_11 = table_11 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_12 = table_12 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_13 = table_13 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_14 = table_14 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_15 = table_15 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_16 = table_16 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_17 = table_17 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_18 = table_18 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_19 = table_19 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_20 = table_20 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_21 = table_21 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_22 = table_22 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_23 = table_23 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_24 = table_24 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_25 = table_25 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_26 = table_26 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_27 = table_27 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_28 = table_28 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_29 = table_29 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_30 = table_30 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_31 = table_31 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_32 = table_32 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_33 = table_33 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_34 = table_34 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_35 = table_35 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_36 = table_36 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_37 = table_37 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_38 = table_38 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_39 = table_39 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_40 = table_40 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_41 = table_41 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_42 = table_42 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_43 = table_43 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_44 = table_44 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_45 = table_45 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_46 = table_46 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_47 = table_47 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_48 = table_48 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_49 = table_49 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_50 = table_50 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_51 = table_51 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_52 = table_52 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_53 = table_53 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_54 = table_54 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_55 = table_55 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_56 = table_56 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_57 = table_57 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_58 = table_58 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_59 = table_59 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_60 = table_60 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_61 = table_61 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_62 = table_62 == 2'h0; // @[Rename.scala 188:35]
  wire  _T_63 = table_63 == 2'h0; // @[Rename.scala 188:35]
  wire [7:0] lo_lo_lo = {_T_7,_T_6,_T_5,_T_4,_T_3,_T_2,_T_1,1'h0}; // @[Cat.scala 30:58]
  wire [15:0] lo_lo = {_T_15,_T_14,_T_13,_T_12,_T_11,_T_10,_T_9,_T_8,lo_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] lo_hi_lo = {_T_23,_T_22,_T_21,_T_20,_T_19,_T_18,_T_17,_T_16}; // @[Cat.scala 30:58]
  wire [31:0] lo = {_T_31,_T_30,_T_29,_T_28,_T_27,_T_26,_T_25,_T_24,lo_hi_lo,lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_lo_lo = {_T_39,_T_38,_T_37,_T_36,_T_35,_T_34,_T_33,_T_32}; // @[Cat.scala 30:58]
  wire [15:0] hi_lo = {_T_47,_T_46,_T_45,_T_44,_T_43,_T_42,_T_41,_T_40,hi_lo_lo}; // @[Cat.scala 30:58]
  wire [7:0] hi_hi_lo = {_T_55,_T_54,_T_53,_T_52,_T_51,_T_50,_T_49,_T_48}; // @[Cat.scala 30:58]
  wire [31:0] hi = {_T_63,_T_62,_T_61,_T_60,_T_59,_T_58,_T_57,_T_56,hi_hi_lo,hi_lo}; // @[Cat.scala 30:58]
  wire [63:0] fl0 = {hi,lo}; // @[Cat.scala 30:58]
  wire [1:0] _T_128 = fl0[0] + fl0[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_130 = fl0[2] + fl0[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_132 = _T_128 + _T_130; // @[Bitwise.scala 47:55]
  wire [1:0] _T_134 = fl0[4] + fl0[5]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_136 = fl0[6] + fl0[7]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_138 = _T_134 + _T_136; // @[Bitwise.scala 47:55]
  wire [3:0] _T_140 = _T_132 + _T_138; // @[Bitwise.scala 47:55]
  wire [1:0] _T_142 = fl0[8] + fl0[9]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_144 = fl0[10] + fl0[11]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_146 = _T_142 + _T_144; // @[Bitwise.scala 47:55]
  wire [1:0] _T_148 = fl0[12] + fl0[13]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_150 = fl0[14] + fl0[15]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_152 = _T_148 + _T_150; // @[Bitwise.scala 47:55]
  wire [3:0] _T_154 = _T_146 + _T_152; // @[Bitwise.scala 47:55]
  wire [4:0] _T_156 = _T_140 + _T_154; // @[Bitwise.scala 47:55]
  wire [1:0] _T_158 = fl0[16] + fl0[17]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_160 = fl0[18] + fl0[19]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_162 = _T_158 + _T_160; // @[Bitwise.scala 47:55]
  wire [1:0] _T_164 = fl0[20] + fl0[21]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_166 = fl0[22] + fl0[23]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_168 = _T_164 + _T_166; // @[Bitwise.scala 47:55]
  wire [3:0] _T_170 = _T_162 + _T_168; // @[Bitwise.scala 47:55]
  wire [1:0] _T_172 = fl0[24] + fl0[25]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_174 = fl0[26] + fl0[27]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_176 = _T_172 + _T_174; // @[Bitwise.scala 47:55]
  wire [1:0] _T_178 = fl0[28] + fl0[29]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_180 = fl0[30] + fl0[31]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_182 = _T_178 + _T_180; // @[Bitwise.scala 47:55]
  wire [3:0] _T_184 = _T_176 + _T_182; // @[Bitwise.scala 47:55]
  wire [4:0] _T_186 = _T_170 + _T_184; // @[Bitwise.scala 47:55]
  wire [5:0] _T_188 = _T_156 + _T_186; // @[Bitwise.scala 47:55]
  wire [1:0] _T_190 = fl0[32] + fl0[33]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_192 = fl0[34] + fl0[35]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_194 = _T_190 + _T_192; // @[Bitwise.scala 47:55]
  wire [1:0] _T_196 = fl0[36] + fl0[37]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_198 = fl0[38] + fl0[39]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_200 = _T_196 + _T_198; // @[Bitwise.scala 47:55]
  wire [3:0] _T_202 = _T_194 + _T_200; // @[Bitwise.scala 47:55]
  wire [1:0] _T_204 = fl0[40] + fl0[41]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_206 = fl0[42] + fl0[43]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_208 = _T_204 + _T_206; // @[Bitwise.scala 47:55]
  wire [1:0] _T_210 = fl0[44] + fl0[45]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_212 = fl0[46] + fl0[47]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_214 = _T_210 + _T_212; // @[Bitwise.scala 47:55]
  wire [3:0] _T_216 = _T_208 + _T_214; // @[Bitwise.scala 47:55]
  wire [4:0] _T_218 = _T_202 + _T_216; // @[Bitwise.scala 47:55]
  wire [1:0] _T_220 = fl0[48] + fl0[49]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_222 = fl0[50] + fl0[51]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_224 = _T_220 + _T_222; // @[Bitwise.scala 47:55]
  wire [1:0] _T_226 = fl0[52] + fl0[53]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_228 = fl0[54] + fl0[55]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_230 = _T_226 + _T_228; // @[Bitwise.scala 47:55]
  wire [3:0] _T_232 = _T_224 + _T_230; // @[Bitwise.scala 47:55]
  wire [1:0] _T_234 = fl0[56] + fl0[57]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_236 = fl0[58] + fl0[59]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_238 = _T_234 + _T_236; // @[Bitwise.scala 47:55]
  wire [1:0] _T_240 = fl0[60] + fl0[61]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_242 = fl0[62] + fl0[63]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_244 = _T_240 + _T_242; // @[Bitwise.scala 47:55]
  wire [3:0] _T_246 = _T_238 + _T_244; // @[Bitwise.scala 47:55]
  wire [4:0] _T_248 = _T_232 + _T_246; // @[Bitwise.scala 47:55]
  wire [5:0] _T_250 = _T_218 + _T_248; // @[Bitwise.scala 47:55]
  wire [6:0] free_count = _T_188 + _T_250; // @[Bitwise.scala 47:55]
  wire  _T_255 = table_1 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_256 = table_2 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_257 = table_3 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_258 = table_4 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_259 = table_5 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_260 = table_6 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_261 = table_7 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_262 = table_8 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_263 = table_9 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_264 = table_10 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_265 = table_11 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_266 = table_12 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_267 = table_13 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_268 = table_14 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_269 = table_15 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_270 = table_16 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_271 = table_17 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_272 = table_18 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_273 = table_19 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_274 = table_20 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_275 = table_21 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_276 = table_22 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_277 = table_23 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_278 = table_24 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_279 = table_25 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_280 = table_26 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_281 = table_27 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_282 = table_28 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_283 = table_29 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_284 = table_30 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_285 = table_31 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_286 = table_32 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_287 = table_33 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_288 = table_34 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_289 = table_35 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_290 = table_36 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_291 = table_37 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_292 = table_38 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_293 = table_39 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_294 = table_40 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_295 = table_41 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_296 = table_42 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_297 = table_43 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_298 = table_44 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_299 = table_45 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_300 = table_46 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_301 = table_47 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_302 = table_48 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_303 = table_49 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_304 = table_50 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_305 = table_51 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_306 = table_52 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_307 = table_53 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_308 = table_54 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_309 = table_55 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_310 = table_56 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_311 = table_57 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_312 = table_58 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_313 = table_59 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_314 = table_60 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_315 = table_61 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_316 = table_62 == 2'h2; // @[Rename.scala 192:36]
  wire  _T_317 = table_63 == 2'h2; // @[Rename.scala 192:36]
  wire [7:0] lo_lo_lo_1 = {_T_261,_T_260,_T_259,_T_258,_T_257,_T_256,_T_255,1'h0}; // @[Cat.scala 30:58]
  wire [15:0] lo_lo_1 = {_T_269,_T_268,_T_267,_T_266,_T_265,_T_264,_T_263,_T_262,lo_lo_lo_1}; // @[Cat.scala 30:58]
  wire [7:0] lo_hi_lo_1 = {_T_277,_T_276,_T_275,_T_274,_T_273,_T_272,_T_271,_T_270}; // @[Cat.scala 30:58]
  wire [31:0] lo_1 = {_T_285,_T_284,_T_283,_T_282,_T_281,_T_280,_T_279,_T_278,lo_hi_lo_1,lo_lo_1}; // @[Cat.scala 30:58]
  wire [7:0] hi_lo_lo_1 = {_T_293,_T_292,_T_291,_T_290,_T_289,_T_288,_T_287,_T_286}; // @[Cat.scala 30:58]
  wire [15:0] hi_lo_1 = {_T_301,_T_300,_T_299,_T_298,_T_297,_T_296,_T_295,_T_294,hi_lo_lo_1}; // @[Cat.scala 30:58]
  wire [7:0] hi_hi_lo_1 = {_T_309,_T_308,_T_307,_T_306,_T_305,_T_304,_T_303,_T_302}; // @[Cat.scala 30:58]
  wire [31:0] hi_1 = {_T_317,_T_316,_T_315,_T_314,_T_313,_T_312,_T_311,_T_310,hi_hi_lo_1,hi_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _T_318 = {hi_1,lo_1}; // @[Cat.scala 30:58]
  wire  _T_320 = table_1 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_321 = table_2 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_322 = table_3 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_323 = table_4 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_324 = table_5 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_325 = table_6 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_326 = table_7 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_327 = table_8 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_328 = table_9 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_329 = table_10 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_330 = table_11 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_331 = table_12 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_332 = table_13 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_333 = table_14 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_334 = table_15 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_335 = table_16 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_336 = table_17 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_337 = table_18 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_338 = table_19 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_339 = table_20 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_340 = table_21 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_341 = table_22 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_342 = table_23 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_343 = table_24 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_344 = table_25 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_345 = table_26 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_346 = table_27 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_347 = table_28 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_348 = table_29 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_349 = table_30 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_350 = table_31 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_351 = table_32 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_352 = table_33 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_353 = table_34 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_354 = table_35 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_355 = table_36 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_356 = table_37 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_357 = table_38 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_358 = table_39 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_359 = table_40 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_360 = table_41 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_361 = table_42 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_362 = table_43 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_363 = table_44 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_364 = table_45 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_365 = table_46 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_366 = table_47 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_367 = table_48 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_368 = table_49 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_369 = table_50 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_370 = table_51 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_371 = table_52 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_372 = table_53 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_373 = table_54 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_374 = table_55 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_375 = table_56 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_376 = table_57 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_377 = table_58 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_378 = table_59 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_379 = table_60 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_380 = table_61 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_381 = table_62 == 2'h3; // @[Rename.scala 192:77]
  wire  _T_382 = table_63 == 2'h3; // @[Rename.scala 192:77]
  wire [7:0] lo_lo_lo_2 = {_T_326,_T_325,_T_324,_T_323,_T_322,_T_321,_T_320,1'h1}; // @[Cat.scala 30:58]
  wire [15:0] lo_lo_2 = {_T_334,_T_333,_T_332,_T_331,_T_330,_T_329,_T_328,_T_327,lo_lo_lo_2}; // @[Cat.scala 30:58]
  wire [7:0] lo_hi_lo_2 = {_T_342,_T_341,_T_340,_T_339,_T_338,_T_337,_T_336,_T_335}; // @[Cat.scala 30:58]
  wire [31:0] lo_2 = {_T_350,_T_349,_T_348,_T_347,_T_346,_T_345,_T_344,_T_343,lo_hi_lo_2,lo_lo_2}; // @[Cat.scala 30:58]
  wire [7:0] hi_lo_lo_2 = {_T_358,_T_357,_T_356,_T_355,_T_354,_T_353,_T_352,_T_351}; // @[Cat.scala 30:58]
  wire [15:0] hi_lo_2 = {_T_366,_T_365,_T_364,_T_363,_T_362,_T_361,_T_360,_T_359,hi_lo_lo_2}; // @[Cat.scala 30:58]
  wire [7:0] hi_hi_lo_2 = {_T_374,_T_373,_T_372,_T_371,_T_370,_T_369,_T_368,_T_367}; // @[Cat.scala 30:58]
  wire [31:0] hi_2 = {_T_382,_T_381,_T_380,_T_379,_T_378,_T_377,_T_376,_T_375,hi_hi_lo_2,hi_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _T_383 = {hi_2,lo_2}; // @[Cat.scala 30:58]
  wire  _T_384 = io_en & io_rd_req_0; // @[Rename.scala 196:31]
  wire [5:0] _T_449 = fl0[62] ? 6'h3e : 6'h3f; // @[Mux.scala 47:69]
  wire [5:0] _T_450 = fl0[61] ? 6'h3d : _T_449; // @[Mux.scala 47:69]
  wire [5:0] _T_451 = fl0[60] ? 6'h3c : _T_450; // @[Mux.scala 47:69]
  wire [5:0] _T_452 = fl0[59] ? 6'h3b : _T_451; // @[Mux.scala 47:69]
  wire [5:0] _T_453 = fl0[58] ? 6'h3a : _T_452; // @[Mux.scala 47:69]
  wire [5:0] _T_454 = fl0[57] ? 6'h39 : _T_453; // @[Mux.scala 47:69]
  wire [5:0] _T_455 = fl0[56] ? 6'h38 : _T_454; // @[Mux.scala 47:69]
  wire [5:0] _T_456 = fl0[55] ? 6'h37 : _T_455; // @[Mux.scala 47:69]
  wire [5:0] _T_457 = fl0[54] ? 6'h36 : _T_456; // @[Mux.scala 47:69]
  wire [5:0] _T_458 = fl0[53] ? 6'h35 : _T_457; // @[Mux.scala 47:69]
  wire [5:0] _T_459 = fl0[52] ? 6'h34 : _T_458; // @[Mux.scala 47:69]
  wire [5:0] _T_460 = fl0[51] ? 6'h33 : _T_459; // @[Mux.scala 47:69]
  wire [5:0] _T_461 = fl0[50] ? 6'h32 : _T_460; // @[Mux.scala 47:69]
  wire [5:0] _T_462 = fl0[49] ? 6'h31 : _T_461; // @[Mux.scala 47:69]
  wire [5:0] _T_463 = fl0[48] ? 6'h30 : _T_462; // @[Mux.scala 47:69]
  wire [5:0] _T_464 = fl0[47] ? 6'h2f : _T_463; // @[Mux.scala 47:69]
  wire [5:0] _T_465 = fl0[46] ? 6'h2e : _T_464; // @[Mux.scala 47:69]
  wire [5:0] _T_466 = fl0[45] ? 6'h2d : _T_465; // @[Mux.scala 47:69]
  wire [5:0] _T_467 = fl0[44] ? 6'h2c : _T_466; // @[Mux.scala 47:69]
  wire [5:0] _T_468 = fl0[43] ? 6'h2b : _T_467; // @[Mux.scala 47:69]
  wire [5:0] _T_469 = fl0[42] ? 6'h2a : _T_468; // @[Mux.scala 47:69]
  wire [5:0] _T_470 = fl0[41] ? 6'h29 : _T_469; // @[Mux.scala 47:69]
  wire [5:0] _T_471 = fl0[40] ? 6'h28 : _T_470; // @[Mux.scala 47:69]
  wire [5:0] _T_472 = fl0[39] ? 6'h27 : _T_471; // @[Mux.scala 47:69]
  wire [5:0] _T_473 = fl0[38] ? 6'h26 : _T_472; // @[Mux.scala 47:69]
  wire [5:0] _T_474 = fl0[37] ? 6'h25 : _T_473; // @[Mux.scala 47:69]
  wire [5:0] _T_475 = fl0[36] ? 6'h24 : _T_474; // @[Mux.scala 47:69]
  wire [5:0] _T_476 = fl0[35] ? 6'h23 : _T_475; // @[Mux.scala 47:69]
  wire [5:0] _T_477 = fl0[34] ? 6'h22 : _T_476; // @[Mux.scala 47:69]
  wire [5:0] _T_478 = fl0[33] ? 6'h21 : _T_477; // @[Mux.scala 47:69]
  wire [5:0] _T_479 = fl0[32] ? 6'h20 : _T_478; // @[Mux.scala 47:69]
  wire [5:0] _T_480 = fl0[31] ? 6'h1f : _T_479; // @[Mux.scala 47:69]
  wire [5:0] _T_481 = fl0[30] ? 6'h1e : _T_480; // @[Mux.scala 47:69]
  wire [5:0] _T_482 = fl0[29] ? 6'h1d : _T_481; // @[Mux.scala 47:69]
  wire [5:0] _T_483 = fl0[28] ? 6'h1c : _T_482; // @[Mux.scala 47:69]
  wire [5:0] _T_484 = fl0[27] ? 6'h1b : _T_483; // @[Mux.scala 47:69]
  wire [5:0] _T_485 = fl0[26] ? 6'h1a : _T_484; // @[Mux.scala 47:69]
  wire [5:0] _T_486 = fl0[25] ? 6'h19 : _T_485; // @[Mux.scala 47:69]
  wire [5:0] _T_487 = fl0[24] ? 6'h18 : _T_486; // @[Mux.scala 47:69]
  wire [5:0] _T_488 = fl0[23] ? 6'h17 : _T_487; // @[Mux.scala 47:69]
  wire [5:0] _T_489 = fl0[22] ? 6'h16 : _T_488; // @[Mux.scala 47:69]
  wire [5:0] _T_490 = fl0[21] ? 6'h15 : _T_489; // @[Mux.scala 47:69]
  wire [5:0] _T_491 = fl0[20] ? 6'h14 : _T_490; // @[Mux.scala 47:69]
  wire [5:0] _T_492 = fl0[19] ? 6'h13 : _T_491; // @[Mux.scala 47:69]
  wire [5:0] _T_493 = fl0[18] ? 6'h12 : _T_492; // @[Mux.scala 47:69]
  wire [5:0] _T_494 = fl0[17] ? 6'h11 : _T_493; // @[Mux.scala 47:69]
  wire [5:0] _T_495 = fl0[16] ? 6'h10 : _T_494; // @[Mux.scala 47:69]
  wire [5:0] _T_496 = fl0[15] ? 6'hf : _T_495; // @[Mux.scala 47:69]
  wire [5:0] _T_497 = fl0[14] ? 6'he : _T_496; // @[Mux.scala 47:69]
  wire [5:0] _T_498 = fl0[13] ? 6'hd : _T_497; // @[Mux.scala 47:69]
  wire [5:0] _T_499 = fl0[12] ? 6'hc : _T_498; // @[Mux.scala 47:69]
  wire [5:0] _T_500 = fl0[11] ? 6'hb : _T_499; // @[Mux.scala 47:69]
  wire [5:0] _T_501 = fl0[10] ? 6'ha : _T_500; // @[Mux.scala 47:69]
  wire [5:0] _T_502 = fl0[9] ? 6'h9 : _T_501; // @[Mux.scala 47:69]
  wire [5:0] _T_503 = fl0[8] ? 6'h8 : _T_502; // @[Mux.scala 47:69]
  wire [5:0] _T_504 = fl0[7] ? 6'h7 : _T_503; // @[Mux.scala 47:69]
  wire [5:0] _T_505 = fl0[6] ? 6'h6 : _T_504; // @[Mux.scala 47:69]
  wire [5:0] _T_506 = fl0[5] ? 6'h5 : _T_505; // @[Mux.scala 47:69]
  wire [5:0] _T_507 = fl0[4] ? 6'h4 : _T_506; // @[Mux.scala 47:69]
  wire [5:0] _T_508 = fl0[3] ? 6'h3 : _T_507; // @[Mux.scala 47:69]
  wire [5:0] _T_509 = fl0[2] ? 6'h2 : _T_508; // @[Mux.scala 47:69]
  wire [5:0] _T_510 = fl0[1] ? 6'h1 : _T_509; // @[Mux.scala 47:69]
  wire [5:0] _T_511 = fl0[0] ? 6'h0 : _T_510; // @[Mux.scala 47:69]
  wire [63:0] _T_513 = 64'h1 << io_rd_paddr_0; // @[OneHot.scala 65:12]
  wire [63:0] _T_515 = ~_T_513; // @[Rename.scala 198:19]
  wire [63:0] fl1 = fl0 & _T_515; // @[Rename.scala 198:17]
  wire  _T_516 = io_en & io_rd_req_1; // @[Rename.scala 199:31]
  wire [5:0] _T_581 = fl1[62] ? 6'h3e : 6'h3f; // @[Mux.scala 47:69]
  wire [5:0] _T_582 = fl1[61] ? 6'h3d : _T_581; // @[Mux.scala 47:69]
  wire [5:0] _T_583 = fl1[60] ? 6'h3c : _T_582; // @[Mux.scala 47:69]
  wire [5:0] _T_584 = fl1[59] ? 6'h3b : _T_583; // @[Mux.scala 47:69]
  wire [5:0] _T_585 = fl1[58] ? 6'h3a : _T_584; // @[Mux.scala 47:69]
  wire [5:0] _T_586 = fl1[57] ? 6'h39 : _T_585; // @[Mux.scala 47:69]
  wire [5:0] _T_587 = fl1[56] ? 6'h38 : _T_586; // @[Mux.scala 47:69]
  wire [5:0] _T_588 = fl1[55] ? 6'h37 : _T_587; // @[Mux.scala 47:69]
  wire [5:0] _T_589 = fl1[54] ? 6'h36 : _T_588; // @[Mux.scala 47:69]
  wire [5:0] _T_590 = fl1[53] ? 6'h35 : _T_589; // @[Mux.scala 47:69]
  wire [5:0] _T_591 = fl1[52] ? 6'h34 : _T_590; // @[Mux.scala 47:69]
  wire [5:0] _T_592 = fl1[51] ? 6'h33 : _T_591; // @[Mux.scala 47:69]
  wire [5:0] _T_593 = fl1[50] ? 6'h32 : _T_592; // @[Mux.scala 47:69]
  wire [5:0] _T_594 = fl1[49] ? 6'h31 : _T_593; // @[Mux.scala 47:69]
  wire [5:0] _T_595 = fl1[48] ? 6'h30 : _T_594; // @[Mux.scala 47:69]
  wire [5:0] _T_596 = fl1[47] ? 6'h2f : _T_595; // @[Mux.scala 47:69]
  wire [5:0] _T_597 = fl1[46] ? 6'h2e : _T_596; // @[Mux.scala 47:69]
  wire [5:0] _T_598 = fl1[45] ? 6'h2d : _T_597; // @[Mux.scala 47:69]
  wire [5:0] _T_599 = fl1[44] ? 6'h2c : _T_598; // @[Mux.scala 47:69]
  wire [5:0] _T_600 = fl1[43] ? 6'h2b : _T_599; // @[Mux.scala 47:69]
  wire [5:0] _T_601 = fl1[42] ? 6'h2a : _T_600; // @[Mux.scala 47:69]
  wire [5:0] _T_602 = fl1[41] ? 6'h29 : _T_601; // @[Mux.scala 47:69]
  wire [5:0] _T_603 = fl1[40] ? 6'h28 : _T_602; // @[Mux.scala 47:69]
  wire [5:0] _T_604 = fl1[39] ? 6'h27 : _T_603; // @[Mux.scala 47:69]
  wire [5:0] _T_605 = fl1[38] ? 6'h26 : _T_604; // @[Mux.scala 47:69]
  wire [5:0] _T_606 = fl1[37] ? 6'h25 : _T_605; // @[Mux.scala 47:69]
  wire [5:0] _T_607 = fl1[36] ? 6'h24 : _T_606; // @[Mux.scala 47:69]
  wire [5:0] _T_608 = fl1[35] ? 6'h23 : _T_607; // @[Mux.scala 47:69]
  wire [5:0] _T_609 = fl1[34] ? 6'h22 : _T_608; // @[Mux.scala 47:69]
  wire [5:0] _T_610 = fl1[33] ? 6'h21 : _T_609; // @[Mux.scala 47:69]
  wire [5:0] _T_611 = fl1[32] ? 6'h20 : _T_610; // @[Mux.scala 47:69]
  wire [5:0] _T_612 = fl1[31] ? 6'h1f : _T_611; // @[Mux.scala 47:69]
  wire [5:0] _T_613 = fl1[30] ? 6'h1e : _T_612; // @[Mux.scala 47:69]
  wire [5:0] _T_614 = fl1[29] ? 6'h1d : _T_613; // @[Mux.scala 47:69]
  wire [5:0] _T_615 = fl1[28] ? 6'h1c : _T_614; // @[Mux.scala 47:69]
  wire [5:0] _T_616 = fl1[27] ? 6'h1b : _T_615; // @[Mux.scala 47:69]
  wire [5:0] _T_617 = fl1[26] ? 6'h1a : _T_616; // @[Mux.scala 47:69]
  wire [5:0] _T_618 = fl1[25] ? 6'h19 : _T_617; // @[Mux.scala 47:69]
  wire [5:0] _T_619 = fl1[24] ? 6'h18 : _T_618; // @[Mux.scala 47:69]
  wire [5:0] _T_620 = fl1[23] ? 6'h17 : _T_619; // @[Mux.scala 47:69]
  wire [5:0] _T_621 = fl1[22] ? 6'h16 : _T_620; // @[Mux.scala 47:69]
  wire [5:0] _T_622 = fl1[21] ? 6'h15 : _T_621; // @[Mux.scala 47:69]
  wire [5:0] _T_623 = fl1[20] ? 6'h14 : _T_622; // @[Mux.scala 47:69]
  wire [5:0] _T_624 = fl1[19] ? 6'h13 : _T_623; // @[Mux.scala 47:69]
  wire [5:0] _T_625 = fl1[18] ? 6'h12 : _T_624; // @[Mux.scala 47:69]
  wire [5:0] _T_626 = fl1[17] ? 6'h11 : _T_625; // @[Mux.scala 47:69]
  wire [5:0] _T_627 = fl1[16] ? 6'h10 : _T_626; // @[Mux.scala 47:69]
  wire [5:0] _T_628 = fl1[15] ? 6'hf : _T_627; // @[Mux.scala 47:69]
  wire [5:0] _T_629 = fl1[14] ? 6'he : _T_628; // @[Mux.scala 47:69]
  wire [5:0] _T_630 = fl1[13] ? 6'hd : _T_629; // @[Mux.scala 47:69]
  wire [5:0] _T_631 = fl1[12] ? 6'hc : _T_630; // @[Mux.scala 47:69]
  wire [5:0] _T_632 = fl1[11] ? 6'hb : _T_631; // @[Mux.scala 47:69]
  wire [5:0] _T_633 = fl1[10] ? 6'ha : _T_632; // @[Mux.scala 47:69]
  wire [5:0] _T_634 = fl1[9] ? 6'h9 : _T_633; // @[Mux.scala 47:69]
  wire [5:0] _T_635 = fl1[8] ? 6'h8 : _T_634; // @[Mux.scala 47:69]
  wire [5:0] _T_636 = fl1[7] ? 6'h7 : _T_635; // @[Mux.scala 47:69]
  wire [5:0] _T_637 = fl1[6] ? 6'h6 : _T_636; // @[Mux.scala 47:69]
  wire [5:0] _T_638 = fl1[5] ? 6'h5 : _T_637; // @[Mux.scala 47:69]
  wire [5:0] _T_639 = fl1[4] ? 6'h4 : _T_638; // @[Mux.scala 47:69]
  wire [5:0] _T_640 = fl1[3] ? 6'h3 : _T_639; // @[Mux.scala 47:69]
  wire [5:0] _T_641 = fl1[2] ? 6'h2 : _T_640; // @[Mux.scala 47:69]
  wire [5:0] _T_642 = fl1[1] ? 6'h1 : _T_641; // @[Mux.scala 47:69]
  wire [5:0] _T_643 = fl1[0] ? 6'h0 : _T_642; // @[Mux.scala 47:69]
  wire [1:0] _GEN_1 = 6'h1 == io_rd_paddr_0 ? 2'h1 : table_1; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_2 = 6'h2 == io_rd_paddr_0 ? 2'h1 : table_2; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_3 = 6'h3 == io_rd_paddr_0 ? 2'h1 : table_3; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_4 = 6'h4 == io_rd_paddr_0 ? 2'h1 : table_4; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_5 = 6'h5 == io_rd_paddr_0 ? 2'h1 : table_5; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_6 = 6'h6 == io_rd_paddr_0 ? 2'h1 : table_6; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_7 = 6'h7 == io_rd_paddr_0 ? 2'h1 : table_7; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_8 = 6'h8 == io_rd_paddr_0 ? 2'h1 : table_8; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_9 = 6'h9 == io_rd_paddr_0 ? 2'h1 : table_9; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_10 = 6'ha == io_rd_paddr_0 ? 2'h1 : table_10; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_11 = 6'hb == io_rd_paddr_0 ? 2'h1 : table_11; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_12 = 6'hc == io_rd_paddr_0 ? 2'h1 : table_12; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_13 = 6'hd == io_rd_paddr_0 ? 2'h1 : table_13; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_14 = 6'he == io_rd_paddr_0 ? 2'h1 : table_14; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_15 = 6'hf == io_rd_paddr_0 ? 2'h1 : table_15; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_16 = 6'h10 == io_rd_paddr_0 ? 2'h1 : table_16; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_17 = 6'h11 == io_rd_paddr_0 ? 2'h1 : table_17; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_18 = 6'h12 == io_rd_paddr_0 ? 2'h1 : table_18; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_19 = 6'h13 == io_rd_paddr_0 ? 2'h1 : table_19; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_20 = 6'h14 == io_rd_paddr_0 ? 2'h1 : table_20; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_21 = 6'h15 == io_rd_paddr_0 ? 2'h1 : table_21; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_22 = 6'h16 == io_rd_paddr_0 ? 2'h1 : table_22; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_23 = 6'h17 == io_rd_paddr_0 ? 2'h1 : table_23; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_24 = 6'h18 == io_rd_paddr_0 ? 2'h1 : table_24; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_25 = 6'h19 == io_rd_paddr_0 ? 2'h1 : table_25; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_26 = 6'h1a == io_rd_paddr_0 ? 2'h1 : table_26; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_27 = 6'h1b == io_rd_paddr_0 ? 2'h1 : table_27; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_28 = 6'h1c == io_rd_paddr_0 ? 2'h1 : table_28; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_29 = 6'h1d == io_rd_paddr_0 ? 2'h1 : table_29; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_30 = 6'h1e == io_rd_paddr_0 ? 2'h1 : table_30; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_31 = 6'h1f == io_rd_paddr_0 ? 2'h1 : table_31; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_32 = 6'h20 == io_rd_paddr_0 ? 2'h1 : table_32; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_33 = 6'h21 == io_rd_paddr_0 ? 2'h1 : table_33; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_34 = 6'h22 == io_rd_paddr_0 ? 2'h1 : table_34; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_35 = 6'h23 == io_rd_paddr_0 ? 2'h1 : table_35; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_36 = 6'h24 == io_rd_paddr_0 ? 2'h1 : table_36; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_37 = 6'h25 == io_rd_paddr_0 ? 2'h1 : table_37; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_38 = 6'h26 == io_rd_paddr_0 ? 2'h1 : table_38; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_39 = 6'h27 == io_rd_paddr_0 ? 2'h1 : table_39; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_40 = 6'h28 == io_rd_paddr_0 ? 2'h1 : table_40; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_41 = 6'h29 == io_rd_paddr_0 ? 2'h1 : table_41; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_42 = 6'h2a == io_rd_paddr_0 ? 2'h1 : table_42; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_43 = 6'h2b == io_rd_paddr_0 ? 2'h1 : table_43; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_44 = 6'h2c == io_rd_paddr_0 ? 2'h1 : table_44; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_45 = 6'h2d == io_rd_paddr_0 ? 2'h1 : table_45; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_46 = 6'h2e == io_rd_paddr_0 ? 2'h1 : table_46; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_47 = 6'h2f == io_rd_paddr_0 ? 2'h1 : table_47; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_48 = 6'h30 == io_rd_paddr_0 ? 2'h1 : table_48; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_49 = 6'h31 == io_rd_paddr_0 ? 2'h1 : table_49; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_50 = 6'h32 == io_rd_paddr_0 ? 2'h1 : table_50; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_51 = 6'h33 == io_rd_paddr_0 ? 2'h1 : table_51; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_52 = 6'h34 == io_rd_paddr_0 ? 2'h1 : table_52; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_53 = 6'h35 == io_rd_paddr_0 ? 2'h1 : table_53; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_54 = 6'h36 == io_rd_paddr_0 ? 2'h1 : table_54; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_55 = 6'h37 == io_rd_paddr_0 ? 2'h1 : table_55; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_56 = 6'h38 == io_rd_paddr_0 ? 2'h1 : table_56; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_57 = 6'h39 == io_rd_paddr_0 ? 2'h1 : table_57; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_58 = 6'h3a == io_rd_paddr_0 ? 2'h1 : table_58; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_59 = 6'h3b == io_rd_paddr_0 ? 2'h1 : table_59; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_60 = 6'h3c == io_rd_paddr_0 ? 2'h1 : table_60; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_61 = 6'h3d == io_rd_paddr_0 ? 2'h1 : table_61; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_62 = 6'h3e == io_rd_paddr_0 ? 2'h1 : table_62; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_63 = 6'h3f == io_rd_paddr_0 ? 2'h1 : table_63; // @[Rename.scala 186:22 203:{29,29}]
  wire [1:0] _GEN_65 = _T_384 ? _GEN_1 : table_1; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_66 = _T_384 ? _GEN_2 : table_2; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_67 = _T_384 ? _GEN_3 : table_3; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_68 = _T_384 ? _GEN_4 : table_4; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_69 = _T_384 ? _GEN_5 : table_5; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_70 = _T_384 ? _GEN_6 : table_6; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_71 = _T_384 ? _GEN_7 : table_7; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_72 = _T_384 ? _GEN_8 : table_8; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_73 = _T_384 ? _GEN_9 : table_9; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_74 = _T_384 ? _GEN_10 : table_10; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_75 = _T_384 ? _GEN_11 : table_11; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_76 = _T_384 ? _GEN_12 : table_12; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_77 = _T_384 ? _GEN_13 : table_13; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_78 = _T_384 ? _GEN_14 : table_14; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_79 = _T_384 ? _GEN_15 : table_15; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_80 = _T_384 ? _GEN_16 : table_16; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_81 = _T_384 ? _GEN_17 : table_17; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_82 = _T_384 ? _GEN_18 : table_18; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_83 = _T_384 ? _GEN_19 : table_19; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_84 = _T_384 ? _GEN_20 : table_20; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_85 = _T_384 ? _GEN_21 : table_21; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_86 = _T_384 ? _GEN_22 : table_22; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_87 = _T_384 ? _GEN_23 : table_23; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_88 = _T_384 ? _GEN_24 : table_24; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_89 = _T_384 ? _GEN_25 : table_25; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_90 = _T_384 ? _GEN_26 : table_26; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_91 = _T_384 ? _GEN_27 : table_27; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_92 = _T_384 ? _GEN_28 : table_28; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_93 = _T_384 ? _GEN_29 : table_29; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_94 = _T_384 ? _GEN_30 : table_30; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_95 = _T_384 ? _GEN_31 : table_31; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_96 = _T_384 ? _GEN_32 : table_32; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_97 = _T_384 ? _GEN_33 : table_33; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_98 = _T_384 ? _GEN_34 : table_34; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_99 = _T_384 ? _GEN_35 : table_35; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_100 = _T_384 ? _GEN_36 : table_36; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_101 = _T_384 ? _GEN_37 : table_37; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_102 = _T_384 ? _GEN_38 : table_38; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_103 = _T_384 ? _GEN_39 : table_39; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_104 = _T_384 ? _GEN_40 : table_40; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_105 = _T_384 ? _GEN_41 : table_41; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_106 = _T_384 ? _GEN_42 : table_42; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_107 = _T_384 ? _GEN_43 : table_43; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_108 = _T_384 ? _GEN_44 : table_44; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_109 = _T_384 ? _GEN_45 : table_45; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_110 = _T_384 ? _GEN_46 : table_46; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_111 = _T_384 ? _GEN_47 : table_47; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_112 = _T_384 ? _GEN_48 : table_48; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_113 = _T_384 ? _GEN_49 : table_49; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_114 = _T_384 ? _GEN_50 : table_50; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_115 = _T_384 ? _GEN_51 : table_51; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_116 = _T_384 ? _GEN_52 : table_52; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_117 = _T_384 ? _GEN_53 : table_53; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_118 = _T_384 ? _GEN_54 : table_54; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_119 = _T_384 ? _GEN_55 : table_55; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_120 = _T_384 ? _GEN_56 : table_56; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_121 = _T_384 ? _GEN_57 : table_57; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_122 = _T_384 ? _GEN_58 : table_58; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_123 = _T_384 ? _GEN_59 : table_59; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_124 = _T_384 ? _GEN_60 : table_60; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_125 = _T_384 ? _GEN_61 : table_61; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_126 = _T_384 ? _GEN_62 : table_62; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_127 = _T_384 ? _GEN_63 : table_63; // @[Rename.scala 186:22 202:34]
  wire [1:0] _GEN_129 = 6'h1 == io_rd_paddr_1 ? 2'h1 : _GEN_65; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_130 = 6'h2 == io_rd_paddr_1 ? 2'h1 : _GEN_66; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_131 = 6'h3 == io_rd_paddr_1 ? 2'h1 : _GEN_67; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_132 = 6'h4 == io_rd_paddr_1 ? 2'h1 : _GEN_68; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_133 = 6'h5 == io_rd_paddr_1 ? 2'h1 : _GEN_69; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_134 = 6'h6 == io_rd_paddr_1 ? 2'h1 : _GEN_70; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_135 = 6'h7 == io_rd_paddr_1 ? 2'h1 : _GEN_71; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_136 = 6'h8 == io_rd_paddr_1 ? 2'h1 : _GEN_72; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_137 = 6'h9 == io_rd_paddr_1 ? 2'h1 : _GEN_73; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_138 = 6'ha == io_rd_paddr_1 ? 2'h1 : _GEN_74; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_139 = 6'hb == io_rd_paddr_1 ? 2'h1 : _GEN_75; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_140 = 6'hc == io_rd_paddr_1 ? 2'h1 : _GEN_76; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_141 = 6'hd == io_rd_paddr_1 ? 2'h1 : _GEN_77; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_142 = 6'he == io_rd_paddr_1 ? 2'h1 : _GEN_78; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_143 = 6'hf == io_rd_paddr_1 ? 2'h1 : _GEN_79; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_144 = 6'h10 == io_rd_paddr_1 ? 2'h1 : _GEN_80; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_145 = 6'h11 == io_rd_paddr_1 ? 2'h1 : _GEN_81; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_146 = 6'h12 == io_rd_paddr_1 ? 2'h1 : _GEN_82; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_147 = 6'h13 == io_rd_paddr_1 ? 2'h1 : _GEN_83; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_148 = 6'h14 == io_rd_paddr_1 ? 2'h1 : _GEN_84; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_149 = 6'h15 == io_rd_paddr_1 ? 2'h1 : _GEN_85; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_150 = 6'h16 == io_rd_paddr_1 ? 2'h1 : _GEN_86; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_151 = 6'h17 == io_rd_paddr_1 ? 2'h1 : _GEN_87; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_152 = 6'h18 == io_rd_paddr_1 ? 2'h1 : _GEN_88; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_153 = 6'h19 == io_rd_paddr_1 ? 2'h1 : _GEN_89; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_154 = 6'h1a == io_rd_paddr_1 ? 2'h1 : _GEN_90; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_155 = 6'h1b == io_rd_paddr_1 ? 2'h1 : _GEN_91; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_156 = 6'h1c == io_rd_paddr_1 ? 2'h1 : _GEN_92; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_157 = 6'h1d == io_rd_paddr_1 ? 2'h1 : _GEN_93; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_158 = 6'h1e == io_rd_paddr_1 ? 2'h1 : _GEN_94; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_159 = 6'h1f == io_rd_paddr_1 ? 2'h1 : _GEN_95; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_160 = 6'h20 == io_rd_paddr_1 ? 2'h1 : _GEN_96; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_161 = 6'h21 == io_rd_paddr_1 ? 2'h1 : _GEN_97; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_162 = 6'h22 == io_rd_paddr_1 ? 2'h1 : _GEN_98; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_163 = 6'h23 == io_rd_paddr_1 ? 2'h1 : _GEN_99; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_164 = 6'h24 == io_rd_paddr_1 ? 2'h1 : _GEN_100; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_165 = 6'h25 == io_rd_paddr_1 ? 2'h1 : _GEN_101; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_166 = 6'h26 == io_rd_paddr_1 ? 2'h1 : _GEN_102; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_167 = 6'h27 == io_rd_paddr_1 ? 2'h1 : _GEN_103; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_168 = 6'h28 == io_rd_paddr_1 ? 2'h1 : _GEN_104; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_169 = 6'h29 == io_rd_paddr_1 ? 2'h1 : _GEN_105; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_170 = 6'h2a == io_rd_paddr_1 ? 2'h1 : _GEN_106; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_171 = 6'h2b == io_rd_paddr_1 ? 2'h1 : _GEN_107; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_172 = 6'h2c == io_rd_paddr_1 ? 2'h1 : _GEN_108; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_173 = 6'h2d == io_rd_paddr_1 ? 2'h1 : _GEN_109; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_174 = 6'h2e == io_rd_paddr_1 ? 2'h1 : _GEN_110; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_175 = 6'h2f == io_rd_paddr_1 ? 2'h1 : _GEN_111; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_176 = 6'h30 == io_rd_paddr_1 ? 2'h1 : _GEN_112; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_177 = 6'h31 == io_rd_paddr_1 ? 2'h1 : _GEN_113; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_178 = 6'h32 == io_rd_paddr_1 ? 2'h1 : _GEN_114; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_179 = 6'h33 == io_rd_paddr_1 ? 2'h1 : _GEN_115; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_180 = 6'h34 == io_rd_paddr_1 ? 2'h1 : _GEN_116; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_181 = 6'h35 == io_rd_paddr_1 ? 2'h1 : _GEN_117; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_182 = 6'h36 == io_rd_paddr_1 ? 2'h1 : _GEN_118; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_183 = 6'h37 == io_rd_paddr_1 ? 2'h1 : _GEN_119; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_184 = 6'h38 == io_rd_paddr_1 ? 2'h1 : _GEN_120; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_185 = 6'h39 == io_rd_paddr_1 ? 2'h1 : _GEN_121; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_186 = 6'h3a == io_rd_paddr_1 ? 2'h1 : _GEN_122; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_187 = 6'h3b == io_rd_paddr_1 ? 2'h1 : _GEN_123; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_188 = 6'h3c == io_rd_paddr_1 ? 2'h1 : _GEN_124; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_189 = 6'h3d == io_rd_paddr_1 ? 2'h1 : _GEN_125; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_190 = 6'h3e == io_rd_paddr_1 ? 2'h1 : _GEN_126; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_191 = 6'h3f == io_rd_paddr_1 ? 2'h1 : _GEN_127; // @[Rename.scala 203:{29,29}]
  wire [1:0] _GEN_193 = _T_516 ? _GEN_129 : _GEN_65; // @[Rename.scala 202:34]
  wire [1:0] _GEN_194 = _T_516 ? _GEN_130 : _GEN_66; // @[Rename.scala 202:34]
  wire [1:0] _GEN_195 = _T_516 ? _GEN_131 : _GEN_67; // @[Rename.scala 202:34]
  wire [1:0] _GEN_196 = _T_516 ? _GEN_132 : _GEN_68; // @[Rename.scala 202:34]
  wire [1:0] _GEN_197 = _T_516 ? _GEN_133 : _GEN_69; // @[Rename.scala 202:34]
  wire [1:0] _GEN_198 = _T_516 ? _GEN_134 : _GEN_70; // @[Rename.scala 202:34]
  wire [1:0] _GEN_199 = _T_516 ? _GEN_135 : _GEN_71; // @[Rename.scala 202:34]
  wire [1:0] _GEN_200 = _T_516 ? _GEN_136 : _GEN_72; // @[Rename.scala 202:34]
  wire [1:0] _GEN_201 = _T_516 ? _GEN_137 : _GEN_73; // @[Rename.scala 202:34]
  wire [1:0] _GEN_202 = _T_516 ? _GEN_138 : _GEN_74; // @[Rename.scala 202:34]
  wire [1:0] _GEN_203 = _T_516 ? _GEN_139 : _GEN_75; // @[Rename.scala 202:34]
  wire [1:0] _GEN_204 = _T_516 ? _GEN_140 : _GEN_76; // @[Rename.scala 202:34]
  wire [1:0] _GEN_205 = _T_516 ? _GEN_141 : _GEN_77; // @[Rename.scala 202:34]
  wire [1:0] _GEN_206 = _T_516 ? _GEN_142 : _GEN_78; // @[Rename.scala 202:34]
  wire [1:0] _GEN_207 = _T_516 ? _GEN_143 : _GEN_79; // @[Rename.scala 202:34]
  wire [1:0] _GEN_208 = _T_516 ? _GEN_144 : _GEN_80; // @[Rename.scala 202:34]
  wire [1:0] _GEN_209 = _T_516 ? _GEN_145 : _GEN_81; // @[Rename.scala 202:34]
  wire [1:0] _GEN_210 = _T_516 ? _GEN_146 : _GEN_82; // @[Rename.scala 202:34]
  wire [1:0] _GEN_211 = _T_516 ? _GEN_147 : _GEN_83; // @[Rename.scala 202:34]
  wire [1:0] _GEN_212 = _T_516 ? _GEN_148 : _GEN_84; // @[Rename.scala 202:34]
  wire [1:0] _GEN_213 = _T_516 ? _GEN_149 : _GEN_85; // @[Rename.scala 202:34]
  wire [1:0] _GEN_214 = _T_516 ? _GEN_150 : _GEN_86; // @[Rename.scala 202:34]
  wire [1:0] _GEN_215 = _T_516 ? _GEN_151 : _GEN_87; // @[Rename.scala 202:34]
  wire [1:0] _GEN_216 = _T_516 ? _GEN_152 : _GEN_88; // @[Rename.scala 202:34]
  wire [1:0] _GEN_217 = _T_516 ? _GEN_153 : _GEN_89; // @[Rename.scala 202:34]
  wire [1:0] _GEN_218 = _T_516 ? _GEN_154 : _GEN_90; // @[Rename.scala 202:34]
  wire [1:0] _GEN_219 = _T_516 ? _GEN_155 : _GEN_91; // @[Rename.scala 202:34]
  wire [1:0] _GEN_220 = _T_516 ? _GEN_156 : _GEN_92; // @[Rename.scala 202:34]
  wire [1:0] _GEN_221 = _T_516 ? _GEN_157 : _GEN_93; // @[Rename.scala 202:34]
  wire [1:0] _GEN_222 = _T_516 ? _GEN_158 : _GEN_94; // @[Rename.scala 202:34]
  wire [1:0] _GEN_223 = _T_516 ? _GEN_159 : _GEN_95; // @[Rename.scala 202:34]
  wire [1:0] _GEN_224 = _T_516 ? _GEN_160 : _GEN_96; // @[Rename.scala 202:34]
  wire [1:0] _GEN_225 = _T_516 ? _GEN_161 : _GEN_97; // @[Rename.scala 202:34]
  wire [1:0] _GEN_226 = _T_516 ? _GEN_162 : _GEN_98; // @[Rename.scala 202:34]
  wire [1:0] _GEN_227 = _T_516 ? _GEN_163 : _GEN_99; // @[Rename.scala 202:34]
  wire [1:0] _GEN_228 = _T_516 ? _GEN_164 : _GEN_100; // @[Rename.scala 202:34]
  wire [1:0] _GEN_229 = _T_516 ? _GEN_165 : _GEN_101; // @[Rename.scala 202:34]
  wire [1:0] _GEN_230 = _T_516 ? _GEN_166 : _GEN_102; // @[Rename.scala 202:34]
  wire [1:0] _GEN_231 = _T_516 ? _GEN_167 : _GEN_103; // @[Rename.scala 202:34]
  wire [1:0] _GEN_232 = _T_516 ? _GEN_168 : _GEN_104; // @[Rename.scala 202:34]
  wire [1:0] _GEN_233 = _T_516 ? _GEN_169 : _GEN_105; // @[Rename.scala 202:34]
  wire [1:0] _GEN_234 = _T_516 ? _GEN_170 : _GEN_106; // @[Rename.scala 202:34]
  wire [1:0] _GEN_235 = _T_516 ? _GEN_171 : _GEN_107; // @[Rename.scala 202:34]
  wire [1:0] _GEN_236 = _T_516 ? _GEN_172 : _GEN_108; // @[Rename.scala 202:34]
  wire [1:0] _GEN_237 = _T_516 ? _GEN_173 : _GEN_109; // @[Rename.scala 202:34]
  wire [1:0] _GEN_238 = _T_516 ? _GEN_174 : _GEN_110; // @[Rename.scala 202:34]
  wire [1:0] _GEN_239 = _T_516 ? _GEN_175 : _GEN_111; // @[Rename.scala 202:34]
  wire [1:0] _GEN_240 = _T_516 ? _GEN_176 : _GEN_112; // @[Rename.scala 202:34]
  wire [1:0] _GEN_241 = _T_516 ? _GEN_177 : _GEN_113; // @[Rename.scala 202:34]
  wire [1:0] _GEN_242 = _T_516 ? _GEN_178 : _GEN_114; // @[Rename.scala 202:34]
  wire [1:0] _GEN_243 = _T_516 ? _GEN_179 : _GEN_115; // @[Rename.scala 202:34]
  wire [1:0] _GEN_244 = _T_516 ? _GEN_180 : _GEN_116; // @[Rename.scala 202:34]
  wire [1:0] _GEN_245 = _T_516 ? _GEN_181 : _GEN_117; // @[Rename.scala 202:34]
  wire [1:0] _GEN_246 = _T_516 ? _GEN_182 : _GEN_118; // @[Rename.scala 202:34]
  wire [1:0] _GEN_247 = _T_516 ? _GEN_183 : _GEN_119; // @[Rename.scala 202:34]
  wire [1:0] _GEN_248 = _T_516 ? _GEN_184 : _GEN_120; // @[Rename.scala 202:34]
  wire [1:0] _GEN_249 = _T_516 ? _GEN_185 : _GEN_121; // @[Rename.scala 202:34]
  wire [1:0] _GEN_250 = _T_516 ? _GEN_186 : _GEN_122; // @[Rename.scala 202:34]
  wire [1:0] _GEN_251 = _T_516 ? _GEN_187 : _GEN_123; // @[Rename.scala 202:34]
  wire [1:0] _GEN_252 = _T_516 ? _GEN_188 : _GEN_124; // @[Rename.scala 202:34]
  wire [1:0] _GEN_253 = _T_516 ? _GEN_189 : _GEN_125; // @[Rename.scala 202:34]
  wire [1:0] _GEN_254 = _T_516 ? _GEN_190 : _GEN_126; // @[Rename.scala 202:34]
  wire [1:0] _GEN_255 = _T_516 ? _GEN_191 : _GEN_127; // @[Rename.scala 202:34]
  wire [1:0] _GEN_257 = 6'h1 == io_exe_0 ? 2'h2 : _GEN_193; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_258 = 6'h2 == io_exe_0 ? 2'h2 : _GEN_194; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_259 = 6'h3 == io_exe_0 ? 2'h2 : _GEN_195; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_260 = 6'h4 == io_exe_0 ? 2'h2 : _GEN_196; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_261 = 6'h5 == io_exe_0 ? 2'h2 : _GEN_197; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_262 = 6'h6 == io_exe_0 ? 2'h2 : _GEN_198; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_263 = 6'h7 == io_exe_0 ? 2'h2 : _GEN_199; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_264 = 6'h8 == io_exe_0 ? 2'h2 : _GEN_200; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_265 = 6'h9 == io_exe_0 ? 2'h2 : _GEN_201; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_266 = 6'ha == io_exe_0 ? 2'h2 : _GEN_202; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_267 = 6'hb == io_exe_0 ? 2'h2 : _GEN_203; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_268 = 6'hc == io_exe_0 ? 2'h2 : _GEN_204; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_269 = 6'hd == io_exe_0 ? 2'h2 : _GEN_205; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_270 = 6'he == io_exe_0 ? 2'h2 : _GEN_206; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_271 = 6'hf == io_exe_0 ? 2'h2 : _GEN_207; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_272 = 6'h10 == io_exe_0 ? 2'h2 : _GEN_208; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_273 = 6'h11 == io_exe_0 ? 2'h2 : _GEN_209; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_274 = 6'h12 == io_exe_0 ? 2'h2 : _GEN_210; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_275 = 6'h13 == io_exe_0 ? 2'h2 : _GEN_211; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_276 = 6'h14 == io_exe_0 ? 2'h2 : _GEN_212; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_277 = 6'h15 == io_exe_0 ? 2'h2 : _GEN_213; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_278 = 6'h16 == io_exe_0 ? 2'h2 : _GEN_214; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_279 = 6'h17 == io_exe_0 ? 2'h2 : _GEN_215; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_280 = 6'h18 == io_exe_0 ? 2'h2 : _GEN_216; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_281 = 6'h19 == io_exe_0 ? 2'h2 : _GEN_217; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_282 = 6'h1a == io_exe_0 ? 2'h2 : _GEN_218; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_283 = 6'h1b == io_exe_0 ? 2'h2 : _GEN_219; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_284 = 6'h1c == io_exe_0 ? 2'h2 : _GEN_220; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_285 = 6'h1d == io_exe_0 ? 2'h2 : _GEN_221; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_286 = 6'h1e == io_exe_0 ? 2'h2 : _GEN_222; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_287 = 6'h1f == io_exe_0 ? 2'h2 : _GEN_223; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_288 = 6'h20 == io_exe_0 ? 2'h2 : _GEN_224; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_289 = 6'h21 == io_exe_0 ? 2'h2 : _GEN_225; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_290 = 6'h22 == io_exe_0 ? 2'h2 : _GEN_226; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_291 = 6'h23 == io_exe_0 ? 2'h2 : _GEN_227; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_292 = 6'h24 == io_exe_0 ? 2'h2 : _GEN_228; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_293 = 6'h25 == io_exe_0 ? 2'h2 : _GEN_229; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_294 = 6'h26 == io_exe_0 ? 2'h2 : _GEN_230; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_295 = 6'h27 == io_exe_0 ? 2'h2 : _GEN_231; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_296 = 6'h28 == io_exe_0 ? 2'h2 : _GEN_232; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_297 = 6'h29 == io_exe_0 ? 2'h2 : _GEN_233; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_298 = 6'h2a == io_exe_0 ? 2'h2 : _GEN_234; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_299 = 6'h2b == io_exe_0 ? 2'h2 : _GEN_235; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_300 = 6'h2c == io_exe_0 ? 2'h2 : _GEN_236; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_301 = 6'h2d == io_exe_0 ? 2'h2 : _GEN_237; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_302 = 6'h2e == io_exe_0 ? 2'h2 : _GEN_238; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_303 = 6'h2f == io_exe_0 ? 2'h2 : _GEN_239; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_304 = 6'h30 == io_exe_0 ? 2'h2 : _GEN_240; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_305 = 6'h31 == io_exe_0 ? 2'h2 : _GEN_241; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_306 = 6'h32 == io_exe_0 ? 2'h2 : _GEN_242; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_307 = 6'h33 == io_exe_0 ? 2'h2 : _GEN_243; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_308 = 6'h34 == io_exe_0 ? 2'h2 : _GEN_244; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_309 = 6'h35 == io_exe_0 ? 2'h2 : _GEN_245; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_310 = 6'h36 == io_exe_0 ? 2'h2 : _GEN_246; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_311 = 6'h37 == io_exe_0 ? 2'h2 : _GEN_247; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_312 = 6'h38 == io_exe_0 ? 2'h2 : _GEN_248; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_313 = 6'h39 == io_exe_0 ? 2'h2 : _GEN_249; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_314 = 6'h3a == io_exe_0 ? 2'h2 : _GEN_250; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_315 = 6'h3b == io_exe_0 ? 2'h2 : _GEN_251; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_316 = 6'h3c == io_exe_0 ? 2'h2 : _GEN_252; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_317 = 6'h3d == io_exe_0 ? 2'h2 : _GEN_253; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_318 = 6'h3e == io_exe_0 ? 2'h2 : _GEN_254; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_319 = 6'h3f == io_exe_0 ? 2'h2 : _GEN_255; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_321 = io_exe_0 != 6'h0 ? _GEN_257 : _GEN_193; // @[Rename.scala 208:30]
  wire [1:0] _GEN_322 = io_exe_0 != 6'h0 ? _GEN_258 : _GEN_194; // @[Rename.scala 208:30]
  wire [1:0] _GEN_323 = io_exe_0 != 6'h0 ? _GEN_259 : _GEN_195; // @[Rename.scala 208:30]
  wire [1:0] _GEN_324 = io_exe_0 != 6'h0 ? _GEN_260 : _GEN_196; // @[Rename.scala 208:30]
  wire [1:0] _GEN_325 = io_exe_0 != 6'h0 ? _GEN_261 : _GEN_197; // @[Rename.scala 208:30]
  wire [1:0] _GEN_326 = io_exe_0 != 6'h0 ? _GEN_262 : _GEN_198; // @[Rename.scala 208:30]
  wire [1:0] _GEN_327 = io_exe_0 != 6'h0 ? _GEN_263 : _GEN_199; // @[Rename.scala 208:30]
  wire [1:0] _GEN_328 = io_exe_0 != 6'h0 ? _GEN_264 : _GEN_200; // @[Rename.scala 208:30]
  wire [1:0] _GEN_329 = io_exe_0 != 6'h0 ? _GEN_265 : _GEN_201; // @[Rename.scala 208:30]
  wire [1:0] _GEN_330 = io_exe_0 != 6'h0 ? _GEN_266 : _GEN_202; // @[Rename.scala 208:30]
  wire [1:0] _GEN_331 = io_exe_0 != 6'h0 ? _GEN_267 : _GEN_203; // @[Rename.scala 208:30]
  wire [1:0] _GEN_332 = io_exe_0 != 6'h0 ? _GEN_268 : _GEN_204; // @[Rename.scala 208:30]
  wire [1:0] _GEN_333 = io_exe_0 != 6'h0 ? _GEN_269 : _GEN_205; // @[Rename.scala 208:30]
  wire [1:0] _GEN_334 = io_exe_0 != 6'h0 ? _GEN_270 : _GEN_206; // @[Rename.scala 208:30]
  wire [1:0] _GEN_335 = io_exe_0 != 6'h0 ? _GEN_271 : _GEN_207; // @[Rename.scala 208:30]
  wire [1:0] _GEN_336 = io_exe_0 != 6'h0 ? _GEN_272 : _GEN_208; // @[Rename.scala 208:30]
  wire [1:0] _GEN_337 = io_exe_0 != 6'h0 ? _GEN_273 : _GEN_209; // @[Rename.scala 208:30]
  wire [1:0] _GEN_338 = io_exe_0 != 6'h0 ? _GEN_274 : _GEN_210; // @[Rename.scala 208:30]
  wire [1:0] _GEN_339 = io_exe_0 != 6'h0 ? _GEN_275 : _GEN_211; // @[Rename.scala 208:30]
  wire [1:0] _GEN_340 = io_exe_0 != 6'h0 ? _GEN_276 : _GEN_212; // @[Rename.scala 208:30]
  wire [1:0] _GEN_341 = io_exe_0 != 6'h0 ? _GEN_277 : _GEN_213; // @[Rename.scala 208:30]
  wire [1:0] _GEN_342 = io_exe_0 != 6'h0 ? _GEN_278 : _GEN_214; // @[Rename.scala 208:30]
  wire [1:0] _GEN_343 = io_exe_0 != 6'h0 ? _GEN_279 : _GEN_215; // @[Rename.scala 208:30]
  wire [1:0] _GEN_344 = io_exe_0 != 6'h0 ? _GEN_280 : _GEN_216; // @[Rename.scala 208:30]
  wire [1:0] _GEN_345 = io_exe_0 != 6'h0 ? _GEN_281 : _GEN_217; // @[Rename.scala 208:30]
  wire [1:0] _GEN_346 = io_exe_0 != 6'h0 ? _GEN_282 : _GEN_218; // @[Rename.scala 208:30]
  wire [1:0] _GEN_347 = io_exe_0 != 6'h0 ? _GEN_283 : _GEN_219; // @[Rename.scala 208:30]
  wire [1:0] _GEN_348 = io_exe_0 != 6'h0 ? _GEN_284 : _GEN_220; // @[Rename.scala 208:30]
  wire [1:0] _GEN_349 = io_exe_0 != 6'h0 ? _GEN_285 : _GEN_221; // @[Rename.scala 208:30]
  wire [1:0] _GEN_350 = io_exe_0 != 6'h0 ? _GEN_286 : _GEN_222; // @[Rename.scala 208:30]
  wire [1:0] _GEN_351 = io_exe_0 != 6'h0 ? _GEN_287 : _GEN_223; // @[Rename.scala 208:30]
  wire [1:0] _GEN_352 = io_exe_0 != 6'h0 ? _GEN_288 : _GEN_224; // @[Rename.scala 208:30]
  wire [1:0] _GEN_353 = io_exe_0 != 6'h0 ? _GEN_289 : _GEN_225; // @[Rename.scala 208:30]
  wire [1:0] _GEN_354 = io_exe_0 != 6'h0 ? _GEN_290 : _GEN_226; // @[Rename.scala 208:30]
  wire [1:0] _GEN_355 = io_exe_0 != 6'h0 ? _GEN_291 : _GEN_227; // @[Rename.scala 208:30]
  wire [1:0] _GEN_356 = io_exe_0 != 6'h0 ? _GEN_292 : _GEN_228; // @[Rename.scala 208:30]
  wire [1:0] _GEN_357 = io_exe_0 != 6'h0 ? _GEN_293 : _GEN_229; // @[Rename.scala 208:30]
  wire [1:0] _GEN_358 = io_exe_0 != 6'h0 ? _GEN_294 : _GEN_230; // @[Rename.scala 208:30]
  wire [1:0] _GEN_359 = io_exe_0 != 6'h0 ? _GEN_295 : _GEN_231; // @[Rename.scala 208:30]
  wire [1:0] _GEN_360 = io_exe_0 != 6'h0 ? _GEN_296 : _GEN_232; // @[Rename.scala 208:30]
  wire [1:0] _GEN_361 = io_exe_0 != 6'h0 ? _GEN_297 : _GEN_233; // @[Rename.scala 208:30]
  wire [1:0] _GEN_362 = io_exe_0 != 6'h0 ? _GEN_298 : _GEN_234; // @[Rename.scala 208:30]
  wire [1:0] _GEN_363 = io_exe_0 != 6'h0 ? _GEN_299 : _GEN_235; // @[Rename.scala 208:30]
  wire [1:0] _GEN_364 = io_exe_0 != 6'h0 ? _GEN_300 : _GEN_236; // @[Rename.scala 208:30]
  wire [1:0] _GEN_365 = io_exe_0 != 6'h0 ? _GEN_301 : _GEN_237; // @[Rename.scala 208:30]
  wire [1:0] _GEN_366 = io_exe_0 != 6'h0 ? _GEN_302 : _GEN_238; // @[Rename.scala 208:30]
  wire [1:0] _GEN_367 = io_exe_0 != 6'h0 ? _GEN_303 : _GEN_239; // @[Rename.scala 208:30]
  wire [1:0] _GEN_368 = io_exe_0 != 6'h0 ? _GEN_304 : _GEN_240; // @[Rename.scala 208:30]
  wire [1:0] _GEN_369 = io_exe_0 != 6'h0 ? _GEN_305 : _GEN_241; // @[Rename.scala 208:30]
  wire [1:0] _GEN_370 = io_exe_0 != 6'h0 ? _GEN_306 : _GEN_242; // @[Rename.scala 208:30]
  wire [1:0] _GEN_371 = io_exe_0 != 6'h0 ? _GEN_307 : _GEN_243; // @[Rename.scala 208:30]
  wire [1:0] _GEN_372 = io_exe_0 != 6'h0 ? _GEN_308 : _GEN_244; // @[Rename.scala 208:30]
  wire [1:0] _GEN_373 = io_exe_0 != 6'h0 ? _GEN_309 : _GEN_245; // @[Rename.scala 208:30]
  wire [1:0] _GEN_374 = io_exe_0 != 6'h0 ? _GEN_310 : _GEN_246; // @[Rename.scala 208:30]
  wire [1:0] _GEN_375 = io_exe_0 != 6'h0 ? _GEN_311 : _GEN_247; // @[Rename.scala 208:30]
  wire [1:0] _GEN_376 = io_exe_0 != 6'h0 ? _GEN_312 : _GEN_248; // @[Rename.scala 208:30]
  wire [1:0] _GEN_377 = io_exe_0 != 6'h0 ? _GEN_313 : _GEN_249; // @[Rename.scala 208:30]
  wire [1:0] _GEN_378 = io_exe_0 != 6'h0 ? _GEN_314 : _GEN_250; // @[Rename.scala 208:30]
  wire [1:0] _GEN_379 = io_exe_0 != 6'h0 ? _GEN_315 : _GEN_251; // @[Rename.scala 208:30]
  wire [1:0] _GEN_380 = io_exe_0 != 6'h0 ? _GEN_316 : _GEN_252; // @[Rename.scala 208:30]
  wire [1:0] _GEN_381 = io_exe_0 != 6'h0 ? _GEN_317 : _GEN_253; // @[Rename.scala 208:30]
  wire [1:0] _GEN_382 = io_exe_0 != 6'h0 ? _GEN_318 : _GEN_254; // @[Rename.scala 208:30]
  wire [1:0] _GEN_383 = io_exe_0 != 6'h0 ? _GEN_319 : _GEN_255; // @[Rename.scala 208:30]
  wire [1:0] _GEN_385 = 6'h1 == io_exe_1 ? 2'h2 : _GEN_321; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_386 = 6'h2 == io_exe_1 ? 2'h2 : _GEN_322; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_387 = 6'h3 == io_exe_1 ? 2'h2 : _GEN_323; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_388 = 6'h4 == io_exe_1 ? 2'h2 : _GEN_324; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_389 = 6'h5 == io_exe_1 ? 2'h2 : _GEN_325; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_390 = 6'h6 == io_exe_1 ? 2'h2 : _GEN_326; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_391 = 6'h7 == io_exe_1 ? 2'h2 : _GEN_327; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_392 = 6'h8 == io_exe_1 ? 2'h2 : _GEN_328; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_393 = 6'h9 == io_exe_1 ? 2'h2 : _GEN_329; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_394 = 6'ha == io_exe_1 ? 2'h2 : _GEN_330; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_395 = 6'hb == io_exe_1 ? 2'h2 : _GEN_331; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_396 = 6'hc == io_exe_1 ? 2'h2 : _GEN_332; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_397 = 6'hd == io_exe_1 ? 2'h2 : _GEN_333; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_398 = 6'he == io_exe_1 ? 2'h2 : _GEN_334; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_399 = 6'hf == io_exe_1 ? 2'h2 : _GEN_335; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_400 = 6'h10 == io_exe_1 ? 2'h2 : _GEN_336; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_401 = 6'h11 == io_exe_1 ? 2'h2 : _GEN_337; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_402 = 6'h12 == io_exe_1 ? 2'h2 : _GEN_338; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_403 = 6'h13 == io_exe_1 ? 2'h2 : _GEN_339; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_404 = 6'h14 == io_exe_1 ? 2'h2 : _GEN_340; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_405 = 6'h15 == io_exe_1 ? 2'h2 : _GEN_341; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_406 = 6'h16 == io_exe_1 ? 2'h2 : _GEN_342; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_407 = 6'h17 == io_exe_1 ? 2'h2 : _GEN_343; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_408 = 6'h18 == io_exe_1 ? 2'h2 : _GEN_344; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_409 = 6'h19 == io_exe_1 ? 2'h2 : _GEN_345; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_410 = 6'h1a == io_exe_1 ? 2'h2 : _GEN_346; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_411 = 6'h1b == io_exe_1 ? 2'h2 : _GEN_347; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_412 = 6'h1c == io_exe_1 ? 2'h2 : _GEN_348; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_413 = 6'h1d == io_exe_1 ? 2'h2 : _GEN_349; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_414 = 6'h1e == io_exe_1 ? 2'h2 : _GEN_350; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_415 = 6'h1f == io_exe_1 ? 2'h2 : _GEN_351; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_416 = 6'h20 == io_exe_1 ? 2'h2 : _GEN_352; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_417 = 6'h21 == io_exe_1 ? 2'h2 : _GEN_353; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_418 = 6'h22 == io_exe_1 ? 2'h2 : _GEN_354; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_419 = 6'h23 == io_exe_1 ? 2'h2 : _GEN_355; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_420 = 6'h24 == io_exe_1 ? 2'h2 : _GEN_356; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_421 = 6'h25 == io_exe_1 ? 2'h2 : _GEN_357; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_422 = 6'h26 == io_exe_1 ? 2'h2 : _GEN_358; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_423 = 6'h27 == io_exe_1 ? 2'h2 : _GEN_359; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_424 = 6'h28 == io_exe_1 ? 2'h2 : _GEN_360; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_425 = 6'h29 == io_exe_1 ? 2'h2 : _GEN_361; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_426 = 6'h2a == io_exe_1 ? 2'h2 : _GEN_362; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_427 = 6'h2b == io_exe_1 ? 2'h2 : _GEN_363; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_428 = 6'h2c == io_exe_1 ? 2'h2 : _GEN_364; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_429 = 6'h2d == io_exe_1 ? 2'h2 : _GEN_365; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_430 = 6'h2e == io_exe_1 ? 2'h2 : _GEN_366; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_431 = 6'h2f == io_exe_1 ? 2'h2 : _GEN_367; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_432 = 6'h30 == io_exe_1 ? 2'h2 : _GEN_368; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_433 = 6'h31 == io_exe_1 ? 2'h2 : _GEN_369; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_434 = 6'h32 == io_exe_1 ? 2'h2 : _GEN_370; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_435 = 6'h33 == io_exe_1 ? 2'h2 : _GEN_371; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_436 = 6'h34 == io_exe_1 ? 2'h2 : _GEN_372; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_437 = 6'h35 == io_exe_1 ? 2'h2 : _GEN_373; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_438 = 6'h36 == io_exe_1 ? 2'h2 : _GEN_374; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_439 = 6'h37 == io_exe_1 ? 2'h2 : _GEN_375; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_440 = 6'h38 == io_exe_1 ? 2'h2 : _GEN_376; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_441 = 6'h39 == io_exe_1 ? 2'h2 : _GEN_377; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_442 = 6'h3a == io_exe_1 ? 2'h2 : _GEN_378; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_443 = 6'h3b == io_exe_1 ? 2'h2 : _GEN_379; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_444 = 6'h3c == io_exe_1 ? 2'h2 : _GEN_380; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_445 = 6'h3d == io_exe_1 ? 2'h2 : _GEN_381; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_446 = 6'h3e == io_exe_1 ? 2'h2 : _GEN_382; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_447 = 6'h3f == io_exe_1 ? 2'h2 : _GEN_383; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_449 = io_exe_1 != 6'h0 ? _GEN_385 : _GEN_321; // @[Rename.scala 208:30]
  wire [1:0] _GEN_450 = io_exe_1 != 6'h0 ? _GEN_386 : _GEN_322; // @[Rename.scala 208:30]
  wire [1:0] _GEN_451 = io_exe_1 != 6'h0 ? _GEN_387 : _GEN_323; // @[Rename.scala 208:30]
  wire [1:0] _GEN_452 = io_exe_1 != 6'h0 ? _GEN_388 : _GEN_324; // @[Rename.scala 208:30]
  wire [1:0] _GEN_453 = io_exe_1 != 6'h0 ? _GEN_389 : _GEN_325; // @[Rename.scala 208:30]
  wire [1:0] _GEN_454 = io_exe_1 != 6'h0 ? _GEN_390 : _GEN_326; // @[Rename.scala 208:30]
  wire [1:0] _GEN_455 = io_exe_1 != 6'h0 ? _GEN_391 : _GEN_327; // @[Rename.scala 208:30]
  wire [1:0] _GEN_456 = io_exe_1 != 6'h0 ? _GEN_392 : _GEN_328; // @[Rename.scala 208:30]
  wire [1:0] _GEN_457 = io_exe_1 != 6'h0 ? _GEN_393 : _GEN_329; // @[Rename.scala 208:30]
  wire [1:0] _GEN_458 = io_exe_1 != 6'h0 ? _GEN_394 : _GEN_330; // @[Rename.scala 208:30]
  wire [1:0] _GEN_459 = io_exe_1 != 6'h0 ? _GEN_395 : _GEN_331; // @[Rename.scala 208:30]
  wire [1:0] _GEN_460 = io_exe_1 != 6'h0 ? _GEN_396 : _GEN_332; // @[Rename.scala 208:30]
  wire [1:0] _GEN_461 = io_exe_1 != 6'h0 ? _GEN_397 : _GEN_333; // @[Rename.scala 208:30]
  wire [1:0] _GEN_462 = io_exe_1 != 6'h0 ? _GEN_398 : _GEN_334; // @[Rename.scala 208:30]
  wire [1:0] _GEN_463 = io_exe_1 != 6'h0 ? _GEN_399 : _GEN_335; // @[Rename.scala 208:30]
  wire [1:0] _GEN_464 = io_exe_1 != 6'h0 ? _GEN_400 : _GEN_336; // @[Rename.scala 208:30]
  wire [1:0] _GEN_465 = io_exe_1 != 6'h0 ? _GEN_401 : _GEN_337; // @[Rename.scala 208:30]
  wire [1:0] _GEN_466 = io_exe_1 != 6'h0 ? _GEN_402 : _GEN_338; // @[Rename.scala 208:30]
  wire [1:0] _GEN_467 = io_exe_1 != 6'h0 ? _GEN_403 : _GEN_339; // @[Rename.scala 208:30]
  wire [1:0] _GEN_468 = io_exe_1 != 6'h0 ? _GEN_404 : _GEN_340; // @[Rename.scala 208:30]
  wire [1:0] _GEN_469 = io_exe_1 != 6'h0 ? _GEN_405 : _GEN_341; // @[Rename.scala 208:30]
  wire [1:0] _GEN_470 = io_exe_1 != 6'h0 ? _GEN_406 : _GEN_342; // @[Rename.scala 208:30]
  wire [1:0] _GEN_471 = io_exe_1 != 6'h0 ? _GEN_407 : _GEN_343; // @[Rename.scala 208:30]
  wire [1:0] _GEN_472 = io_exe_1 != 6'h0 ? _GEN_408 : _GEN_344; // @[Rename.scala 208:30]
  wire [1:0] _GEN_473 = io_exe_1 != 6'h0 ? _GEN_409 : _GEN_345; // @[Rename.scala 208:30]
  wire [1:0] _GEN_474 = io_exe_1 != 6'h0 ? _GEN_410 : _GEN_346; // @[Rename.scala 208:30]
  wire [1:0] _GEN_475 = io_exe_1 != 6'h0 ? _GEN_411 : _GEN_347; // @[Rename.scala 208:30]
  wire [1:0] _GEN_476 = io_exe_1 != 6'h0 ? _GEN_412 : _GEN_348; // @[Rename.scala 208:30]
  wire [1:0] _GEN_477 = io_exe_1 != 6'h0 ? _GEN_413 : _GEN_349; // @[Rename.scala 208:30]
  wire [1:0] _GEN_478 = io_exe_1 != 6'h0 ? _GEN_414 : _GEN_350; // @[Rename.scala 208:30]
  wire [1:0] _GEN_479 = io_exe_1 != 6'h0 ? _GEN_415 : _GEN_351; // @[Rename.scala 208:30]
  wire [1:0] _GEN_480 = io_exe_1 != 6'h0 ? _GEN_416 : _GEN_352; // @[Rename.scala 208:30]
  wire [1:0] _GEN_481 = io_exe_1 != 6'h0 ? _GEN_417 : _GEN_353; // @[Rename.scala 208:30]
  wire [1:0] _GEN_482 = io_exe_1 != 6'h0 ? _GEN_418 : _GEN_354; // @[Rename.scala 208:30]
  wire [1:0] _GEN_483 = io_exe_1 != 6'h0 ? _GEN_419 : _GEN_355; // @[Rename.scala 208:30]
  wire [1:0] _GEN_484 = io_exe_1 != 6'h0 ? _GEN_420 : _GEN_356; // @[Rename.scala 208:30]
  wire [1:0] _GEN_485 = io_exe_1 != 6'h0 ? _GEN_421 : _GEN_357; // @[Rename.scala 208:30]
  wire [1:0] _GEN_486 = io_exe_1 != 6'h0 ? _GEN_422 : _GEN_358; // @[Rename.scala 208:30]
  wire [1:0] _GEN_487 = io_exe_1 != 6'h0 ? _GEN_423 : _GEN_359; // @[Rename.scala 208:30]
  wire [1:0] _GEN_488 = io_exe_1 != 6'h0 ? _GEN_424 : _GEN_360; // @[Rename.scala 208:30]
  wire [1:0] _GEN_489 = io_exe_1 != 6'h0 ? _GEN_425 : _GEN_361; // @[Rename.scala 208:30]
  wire [1:0] _GEN_490 = io_exe_1 != 6'h0 ? _GEN_426 : _GEN_362; // @[Rename.scala 208:30]
  wire [1:0] _GEN_491 = io_exe_1 != 6'h0 ? _GEN_427 : _GEN_363; // @[Rename.scala 208:30]
  wire [1:0] _GEN_492 = io_exe_1 != 6'h0 ? _GEN_428 : _GEN_364; // @[Rename.scala 208:30]
  wire [1:0] _GEN_493 = io_exe_1 != 6'h0 ? _GEN_429 : _GEN_365; // @[Rename.scala 208:30]
  wire [1:0] _GEN_494 = io_exe_1 != 6'h0 ? _GEN_430 : _GEN_366; // @[Rename.scala 208:30]
  wire [1:0] _GEN_495 = io_exe_1 != 6'h0 ? _GEN_431 : _GEN_367; // @[Rename.scala 208:30]
  wire [1:0] _GEN_496 = io_exe_1 != 6'h0 ? _GEN_432 : _GEN_368; // @[Rename.scala 208:30]
  wire [1:0] _GEN_497 = io_exe_1 != 6'h0 ? _GEN_433 : _GEN_369; // @[Rename.scala 208:30]
  wire [1:0] _GEN_498 = io_exe_1 != 6'h0 ? _GEN_434 : _GEN_370; // @[Rename.scala 208:30]
  wire [1:0] _GEN_499 = io_exe_1 != 6'h0 ? _GEN_435 : _GEN_371; // @[Rename.scala 208:30]
  wire [1:0] _GEN_500 = io_exe_1 != 6'h0 ? _GEN_436 : _GEN_372; // @[Rename.scala 208:30]
  wire [1:0] _GEN_501 = io_exe_1 != 6'h0 ? _GEN_437 : _GEN_373; // @[Rename.scala 208:30]
  wire [1:0] _GEN_502 = io_exe_1 != 6'h0 ? _GEN_438 : _GEN_374; // @[Rename.scala 208:30]
  wire [1:0] _GEN_503 = io_exe_1 != 6'h0 ? _GEN_439 : _GEN_375; // @[Rename.scala 208:30]
  wire [1:0] _GEN_504 = io_exe_1 != 6'h0 ? _GEN_440 : _GEN_376; // @[Rename.scala 208:30]
  wire [1:0] _GEN_505 = io_exe_1 != 6'h0 ? _GEN_441 : _GEN_377; // @[Rename.scala 208:30]
  wire [1:0] _GEN_506 = io_exe_1 != 6'h0 ? _GEN_442 : _GEN_378; // @[Rename.scala 208:30]
  wire [1:0] _GEN_507 = io_exe_1 != 6'h0 ? _GEN_443 : _GEN_379; // @[Rename.scala 208:30]
  wire [1:0] _GEN_508 = io_exe_1 != 6'h0 ? _GEN_444 : _GEN_380; // @[Rename.scala 208:30]
  wire [1:0] _GEN_509 = io_exe_1 != 6'h0 ? _GEN_445 : _GEN_381; // @[Rename.scala 208:30]
  wire [1:0] _GEN_510 = io_exe_1 != 6'h0 ? _GEN_446 : _GEN_382; // @[Rename.scala 208:30]
  wire [1:0] _GEN_511 = io_exe_1 != 6'h0 ? _GEN_447 : _GEN_383; // @[Rename.scala 208:30]
  wire [1:0] _GEN_513 = 6'h1 == io_exe_2 ? 2'h2 : _GEN_449; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_514 = 6'h2 == io_exe_2 ? 2'h2 : _GEN_450; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_515 = 6'h3 == io_exe_2 ? 2'h2 : _GEN_451; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_516 = 6'h4 == io_exe_2 ? 2'h2 : _GEN_452; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_517 = 6'h5 == io_exe_2 ? 2'h2 : _GEN_453; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_518 = 6'h6 == io_exe_2 ? 2'h2 : _GEN_454; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_519 = 6'h7 == io_exe_2 ? 2'h2 : _GEN_455; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_520 = 6'h8 == io_exe_2 ? 2'h2 : _GEN_456; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_521 = 6'h9 == io_exe_2 ? 2'h2 : _GEN_457; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_522 = 6'ha == io_exe_2 ? 2'h2 : _GEN_458; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_523 = 6'hb == io_exe_2 ? 2'h2 : _GEN_459; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_524 = 6'hc == io_exe_2 ? 2'h2 : _GEN_460; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_525 = 6'hd == io_exe_2 ? 2'h2 : _GEN_461; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_526 = 6'he == io_exe_2 ? 2'h2 : _GEN_462; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_527 = 6'hf == io_exe_2 ? 2'h2 : _GEN_463; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_528 = 6'h10 == io_exe_2 ? 2'h2 : _GEN_464; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_529 = 6'h11 == io_exe_2 ? 2'h2 : _GEN_465; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_530 = 6'h12 == io_exe_2 ? 2'h2 : _GEN_466; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_531 = 6'h13 == io_exe_2 ? 2'h2 : _GEN_467; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_532 = 6'h14 == io_exe_2 ? 2'h2 : _GEN_468; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_533 = 6'h15 == io_exe_2 ? 2'h2 : _GEN_469; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_534 = 6'h16 == io_exe_2 ? 2'h2 : _GEN_470; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_535 = 6'h17 == io_exe_2 ? 2'h2 : _GEN_471; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_536 = 6'h18 == io_exe_2 ? 2'h2 : _GEN_472; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_537 = 6'h19 == io_exe_2 ? 2'h2 : _GEN_473; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_538 = 6'h1a == io_exe_2 ? 2'h2 : _GEN_474; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_539 = 6'h1b == io_exe_2 ? 2'h2 : _GEN_475; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_540 = 6'h1c == io_exe_2 ? 2'h2 : _GEN_476; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_541 = 6'h1d == io_exe_2 ? 2'h2 : _GEN_477; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_542 = 6'h1e == io_exe_2 ? 2'h2 : _GEN_478; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_543 = 6'h1f == io_exe_2 ? 2'h2 : _GEN_479; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_544 = 6'h20 == io_exe_2 ? 2'h2 : _GEN_480; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_545 = 6'h21 == io_exe_2 ? 2'h2 : _GEN_481; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_546 = 6'h22 == io_exe_2 ? 2'h2 : _GEN_482; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_547 = 6'h23 == io_exe_2 ? 2'h2 : _GEN_483; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_548 = 6'h24 == io_exe_2 ? 2'h2 : _GEN_484; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_549 = 6'h25 == io_exe_2 ? 2'h2 : _GEN_485; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_550 = 6'h26 == io_exe_2 ? 2'h2 : _GEN_486; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_551 = 6'h27 == io_exe_2 ? 2'h2 : _GEN_487; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_552 = 6'h28 == io_exe_2 ? 2'h2 : _GEN_488; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_553 = 6'h29 == io_exe_2 ? 2'h2 : _GEN_489; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_554 = 6'h2a == io_exe_2 ? 2'h2 : _GEN_490; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_555 = 6'h2b == io_exe_2 ? 2'h2 : _GEN_491; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_556 = 6'h2c == io_exe_2 ? 2'h2 : _GEN_492; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_557 = 6'h2d == io_exe_2 ? 2'h2 : _GEN_493; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_558 = 6'h2e == io_exe_2 ? 2'h2 : _GEN_494; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_559 = 6'h2f == io_exe_2 ? 2'h2 : _GEN_495; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_560 = 6'h30 == io_exe_2 ? 2'h2 : _GEN_496; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_561 = 6'h31 == io_exe_2 ? 2'h2 : _GEN_497; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_562 = 6'h32 == io_exe_2 ? 2'h2 : _GEN_498; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_563 = 6'h33 == io_exe_2 ? 2'h2 : _GEN_499; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_564 = 6'h34 == io_exe_2 ? 2'h2 : _GEN_500; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_565 = 6'h35 == io_exe_2 ? 2'h2 : _GEN_501; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_566 = 6'h36 == io_exe_2 ? 2'h2 : _GEN_502; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_567 = 6'h37 == io_exe_2 ? 2'h2 : _GEN_503; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_568 = 6'h38 == io_exe_2 ? 2'h2 : _GEN_504; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_569 = 6'h39 == io_exe_2 ? 2'h2 : _GEN_505; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_570 = 6'h3a == io_exe_2 ? 2'h2 : _GEN_506; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_571 = 6'h3b == io_exe_2 ? 2'h2 : _GEN_507; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_572 = 6'h3c == io_exe_2 ? 2'h2 : _GEN_508; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_573 = 6'h3d == io_exe_2 ? 2'h2 : _GEN_509; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_574 = 6'h3e == io_exe_2 ? 2'h2 : _GEN_510; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_575 = 6'h3f == io_exe_2 ? 2'h2 : _GEN_511; // @[Rename.scala 209:{24,24}]
  wire [1:0] _GEN_577 = io_exe_2 != 6'h0 ? _GEN_513 : _GEN_449; // @[Rename.scala 208:30]
  wire [1:0] _GEN_578 = io_exe_2 != 6'h0 ? _GEN_514 : _GEN_450; // @[Rename.scala 208:30]
  wire [1:0] _GEN_579 = io_exe_2 != 6'h0 ? _GEN_515 : _GEN_451; // @[Rename.scala 208:30]
  wire [1:0] _GEN_580 = io_exe_2 != 6'h0 ? _GEN_516 : _GEN_452; // @[Rename.scala 208:30]
  wire [1:0] _GEN_581 = io_exe_2 != 6'h0 ? _GEN_517 : _GEN_453; // @[Rename.scala 208:30]
  wire [1:0] _GEN_582 = io_exe_2 != 6'h0 ? _GEN_518 : _GEN_454; // @[Rename.scala 208:30]
  wire [1:0] _GEN_583 = io_exe_2 != 6'h0 ? _GEN_519 : _GEN_455; // @[Rename.scala 208:30]
  wire [1:0] _GEN_584 = io_exe_2 != 6'h0 ? _GEN_520 : _GEN_456; // @[Rename.scala 208:30]
  wire [1:0] _GEN_585 = io_exe_2 != 6'h0 ? _GEN_521 : _GEN_457; // @[Rename.scala 208:30]
  wire [1:0] _GEN_586 = io_exe_2 != 6'h0 ? _GEN_522 : _GEN_458; // @[Rename.scala 208:30]
  wire [1:0] _GEN_587 = io_exe_2 != 6'h0 ? _GEN_523 : _GEN_459; // @[Rename.scala 208:30]
  wire [1:0] _GEN_588 = io_exe_2 != 6'h0 ? _GEN_524 : _GEN_460; // @[Rename.scala 208:30]
  wire [1:0] _GEN_589 = io_exe_2 != 6'h0 ? _GEN_525 : _GEN_461; // @[Rename.scala 208:30]
  wire [1:0] _GEN_590 = io_exe_2 != 6'h0 ? _GEN_526 : _GEN_462; // @[Rename.scala 208:30]
  wire [1:0] _GEN_591 = io_exe_2 != 6'h0 ? _GEN_527 : _GEN_463; // @[Rename.scala 208:30]
  wire [1:0] _GEN_592 = io_exe_2 != 6'h0 ? _GEN_528 : _GEN_464; // @[Rename.scala 208:30]
  wire [1:0] _GEN_593 = io_exe_2 != 6'h0 ? _GEN_529 : _GEN_465; // @[Rename.scala 208:30]
  wire [1:0] _GEN_594 = io_exe_2 != 6'h0 ? _GEN_530 : _GEN_466; // @[Rename.scala 208:30]
  wire [1:0] _GEN_595 = io_exe_2 != 6'h0 ? _GEN_531 : _GEN_467; // @[Rename.scala 208:30]
  wire [1:0] _GEN_596 = io_exe_2 != 6'h0 ? _GEN_532 : _GEN_468; // @[Rename.scala 208:30]
  wire [1:0] _GEN_597 = io_exe_2 != 6'h0 ? _GEN_533 : _GEN_469; // @[Rename.scala 208:30]
  wire [1:0] _GEN_598 = io_exe_2 != 6'h0 ? _GEN_534 : _GEN_470; // @[Rename.scala 208:30]
  wire [1:0] _GEN_599 = io_exe_2 != 6'h0 ? _GEN_535 : _GEN_471; // @[Rename.scala 208:30]
  wire [1:0] _GEN_600 = io_exe_2 != 6'h0 ? _GEN_536 : _GEN_472; // @[Rename.scala 208:30]
  wire [1:0] _GEN_601 = io_exe_2 != 6'h0 ? _GEN_537 : _GEN_473; // @[Rename.scala 208:30]
  wire [1:0] _GEN_602 = io_exe_2 != 6'h0 ? _GEN_538 : _GEN_474; // @[Rename.scala 208:30]
  wire [1:0] _GEN_603 = io_exe_2 != 6'h0 ? _GEN_539 : _GEN_475; // @[Rename.scala 208:30]
  wire [1:0] _GEN_604 = io_exe_2 != 6'h0 ? _GEN_540 : _GEN_476; // @[Rename.scala 208:30]
  wire [1:0] _GEN_605 = io_exe_2 != 6'h0 ? _GEN_541 : _GEN_477; // @[Rename.scala 208:30]
  wire [1:0] _GEN_606 = io_exe_2 != 6'h0 ? _GEN_542 : _GEN_478; // @[Rename.scala 208:30]
  wire [1:0] _GEN_607 = io_exe_2 != 6'h0 ? _GEN_543 : _GEN_479; // @[Rename.scala 208:30]
  wire [1:0] _GEN_608 = io_exe_2 != 6'h0 ? _GEN_544 : _GEN_480; // @[Rename.scala 208:30]
  wire [1:0] _GEN_609 = io_exe_2 != 6'h0 ? _GEN_545 : _GEN_481; // @[Rename.scala 208:30]
  wire [1:0] _GEN_610 = io_exe_2 != 6'h0 ? _GEN_546 : _GEN_482; // @[Rename.scala 208:30]
  wire [1:0] _GEN_611 = io_exe_2 != 6'h0 ? _GEN_547 : _GEN_483; // @[Rename.scala 208:30]
  wire [1:0] _GEN_612 = io_exe_2 != 6'h0 ? _GEN_548 : _GEN_484; // @[Rename.scala 208:30]
  wire [1:0] _GEN_613 = io_exe_2 != 6'h0 ? _GEN_549 : _GEN_485; // @[Rename.scala 208:30]
  wire [1:0] _GEN_614 = io_exe_2 != 6'h0 ? _GEN_550 : _GEN_486; // @[Rename.scala 208:30]
  wire [1:0] _GEN_615 = io_exe_2 != 6'h0 ? _GEN_551 : _GEN_487; // @[Rename.scala 208:30]
  wire [1:0] _GEN_616 = io_exe_2 != 6'h0 ? _GEN_552 : _GEN_488; // @[Rename.scala 208:30]
  wire [1:0] _GEN_617 = io_exe_2 != 6'h0 ? _GEN_553 : _GEN_489; // @[Rename.scala 208:30]
  wire [1:0] _GEN_618 = io_exe_2 != 6'h0 ? _GEN_554 : _GEN_490; // @[Rename.scala 208:30]
  wire [1:0] _GEN_619 = io_exe_2 != 6'h0 ? _GEN_555 : _GEN_491; // @[Rename.scala 208:30]
  wire [1:0] _GEN_620 = io_exe_2 != 6'h0 ? _GEN_556 : _GEN_492; // @[Rename.scala 208:30]
  wire [1:0] _GEN_621 = io_exe_2 != 6'h0 ? _GEN_557 : _GEN_493; // @[Rename.scala 208:30]
  wire [1:0] _GEN_622 = io_exe_2 != 6'h0 ? _GEN_558 : _GEN_494; // @[Rename.scala 208:30]
  wire [1:0] _GEN_623 = io_exe_2 != 6'h0 ? _GEN_559 : _GEN_495; // @[Rename.scala 208:30]
  wire [1:0] _GEN_624 = io_exe_2 != 6'h0 ? _GEN_560 : _GEN_496; // @[Rename.scala 208:30]
  wire [1:0] _GEN_625 = io_exe_2 != 6'h0 ? _GEN_561 : _GEN_497; // @[Rename.scala 208:30]
  wire [1:0] _GEN_626 = io_exe_2 != 6'h0 ? _GEN_562 : _GEN_498; // @[Rename.scala 208:30]
  wire [1:0] _GEN_627 = io_exe_2 != 6'h0 ? _GEN_563 : _GEN_499; // @[Rename.scala 208:30]
  wire [1:0] _GEN_628 = io_exe_2 != 6'h0 ? _GEN_564 : _GEN_500; // @[Rename.scala 208:30]
  wire [1:0] _GEN_629 = io_exe_2 != 6'h0 ? _GEN_565 : _GEN_501; // @[Rename.scala 208:30]
  wire [1:0] _GEN_630 = io_exe_2 != 6'h0 ? _GEN_566 : _GEN_502; // @[Rename.scala 208:30]
  wire [1:0] _GEN_631 = io_exe_2 != 6'h0 ? _GEN_567 : _GEN_503; // @[Rename.scala 208:30]
  wire [1:0] _GEN_632 = io_exe_2 != 6'h0 ? _GEN_568 : _GEN_504; // @[Rename.scala 208:30]
  wire [1:0] _GEN_633 = io_exe_2 != 6'h0 ? _GEN_569 : _GEN_505; // @[Rename.scala 208:30]
  wire [1:0] _GEN_634 = io_exe_2 != 6'h0 ? _GEN_570 : _GEN_506; // @[Rename.scala 208:30]
  wire [1:0] _GEN_635 = io_exe_2 != 6'h0 ? _GEN_571 : _GEN_507; // @[Rename.scala 208:30]
  wire [1:0] _GEN_636 = io_exe_2 != 6'h0 ? _GEN_572 : _GEN_508; // @[Rename.scala 208:30]
  wire [1:0] _GEN_637 = io_exe_2 != 6'h0 ? _GEN_573 : _GEN_509; // @[Rename.scala 208:30]
  wire [1:0] _GEN_638 = io_exe_2 != 6'h0 ? _GEN_574 : _GEN_510; // @[Rename.scala 208:30]
  wire [1:0] _GEN_639 = io_exe_2 != 6'h0 ? _GEN_575 : _GEN_511; // @[Rename.scala 208:30]
  wire [1:0] _GEN_641 = 6'h1 == io_cm_0 ? 2'h3 : _GEN_577; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_642 = 6'h2 == io_cm_0 ? 2'h3 : _GEN_578; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_643 = 6'h3 == io_cm_0 ? 2'h3 : _GEN_579; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_644 = 6'h4 == io_cm_0 ? 2'h3 : _GEN_580; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_645 = 6'h5 == io_cm_0 ? 2'h3 : _GEN_581; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_646 = 6'h6 == io_cm_0 ? 2'h3 : _GEN_582; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_647 = 6'h7 == io_cm_0 ? 2'h3 : _GEN_583; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_648 = 6'h8 == io_cm_0 ? 2'h3 : _GEN_584; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_649 = 6'h9 == io_cm_0 ? 2'h3 : _GEN_585; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_650 = 6'ha == io_cm_0 ? 2'h3 : _GEN_586; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_651 = 6'hb == io_cm_0 ? 2'h3 : _GEN_587; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_652 = 6'hc == io_cm_0 ? 2'h3 : _GEN_588; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_653 = 6'hd == io_cm_0 ? 2'h3 : _GEN_589; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_654 = 6'he == io_cm_0 ? 2'h3 : _GEN_590; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_655 = 6'hf == io_cm_0 ? 2'h3 : _GEN_591; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_656 = 6'h10 == io_cm_0 ? 2'h3 : _GEN_592; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_657 = 6'h11 == io_cm_0 ? 2'h3 : _GEN_593; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_658 = 6'h12 == io_cm_0 ? 2'h3 : _GEN_594; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_659 = 6'h13 == io_cm_0 ? 2'h3 : _GEN_595; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_660 = 6'h14 == io_cm_0 ? 2'h3 : _GEN_596; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_661 = 6'h15 == io_cm_0 ? 2'h3 : _GEN_597; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_662 = 6'h16 == io_cm_0 ? 2'h3 : _GEN_598; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_663 = 6'h17 == io_cm_0 ? 2'h3 : _GEN_599; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_664 = 6'h18 == io_cm_0 ? 2'h3 : _GEN_600; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_665 = 6'h19 == io_cm_0 ? 2'h3 : _GEN_601; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_666 = 6'h1a == io_cm_0 ? 2'h3 : _GEN_602; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_667 = 6'h1b == io_cm_0 ? 2'h3 : _GEN_603; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_668 = 6'h1c == io_cm_0 ? 2'h3 : _GEN_604; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_669 = 6'h1d == io_cm_0 ? 2'h3 : _GEN_605; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_670 = 6'h1e == io_cm_0 ? 2'h3 : _GEN_606; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_671 = 6'h1f == io_cm_0 ? 2'h3 : _GEN_607; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_672 = 6'h20 == io_cm_0 ? 2'h3 : _GEN_608; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_673 = 6'h21 == io_cm_0 ? 2'h3 : _GEN_609; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_674 = 6'h22 == io_cm_0 ? 2'h3 : _GEN_610; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_675 = 6'h23 == io_cm_0 ? 2'h3 : _GEN_611; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_676 = 6'h24 == io_cm_0 ? 2'h3 : _GEN_612; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_677 = 6'h25 == io_cm_0 ? 2'h3 : _GEN_613; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_678 = 6'h26 == io_cm_0 ? 2'h3 : _GEN_614; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_679 = 6'h27 == io_cm_0 ? 2'h3 : _GEN_615; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_680 = 6'h28 == io_cm_0 ? 2'h3 : _GEN_616; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_681 = 6'h29 == io_cm_0 ? 2'h3 : _GEN_617; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_682 = 6'h2a == io_cm_0 ? 2'h3 : _GEN_618; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_683 = 6'h2b == io_cm_0 ? 2'h3 : _GEN_619; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_684 = 6'h2c == io_cm_0 ? 2'h3 : _GEN_620; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_685 = 6'h2d == io_cm_0 ? 2'h3 : _GEN_621; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_686 = 6'h2e == io_cm_0 ? 2'h3 : _GEN_622; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_687 = 6'h2f == io_cm_0 ? 2'h3 : _GEN_623; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_688 = 6'h30 == io_cm_0 ? 2'h3 : _GEN_624; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_689 = 6'h31 == io_cm_0 ? 2'h3 : _GEN_625; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_690 = 6'h32 == io_cm_0 ? 2'h3 : _GEN_626; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_691 = 6'h33 == io_cm_0 ? 2'h3 : _GEN_627; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_692 = 6'h34 == io_cm_0 ? 2'h3 : _GEN_628; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_693 = 6'h35 == io_cm_0 ? 2'h3 : _GEN_629; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_694 = 6'h36 == io_cm_0 ? 2'h3 : _GEN_630; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_695 = 6'h37 == io_cm_0 ? 2'h3 : _GEN_631; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_696 = 6'h38 == io_cm_0 ? 2'h3 : _GEN_632; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_697 = 6'h39 == io_cm_0 ? 2'h3 : _GEN_633; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_698 = 6'h3a == io_cm_0 ? 2'h3 : _GEN_634; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_699 = 6'h3b == io_cm_0 ? 2'h3 : _GEN_635; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_700 = 6'h3c == io_cm_0 ? 2'h3 : _GEN_636; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_701 = 6'h3d == io_cm_0 ? 2'h3 : _GEN_637; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_702 = 6'h3e == io_cm_0 ? 2'h3 : _GEN_638; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_703 = 6'h3f == io_cm_0 ? 2'h3 : _GEN_639; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_705 = io_cm_0 != 6'h0 ? _GEN_641 : _GEN_577; // @[Rename.scala 214:29]
  wire [1:0] _GEN_706 = io_cm_0 != 6'h0 ? _GEN_642 : _GEN_578; // @[Rename.scala 214:29]
  wire [1:0] _GEN_707 = io_cm_0 != 6'h0 ? _GEN_643 : _GEN_579; // @[Rename.scala 214:29]
  wire [1:0] _GEN_708 = io_cm_0 != 6'h0 ? _GEN_644 : _GEN_580; // @[Rename.scala 214:29]
  wire [1:0] _GEN_709 = io_cm_0 != 6'h0 ? _GEN_645 : _GEN_581; // @[Rename.scala 214:29]
  wire [1:0] _GEN_710 = io_cm_0 != 6'h0 ? _GEN_646 : _GEN_582; // @[Rename.scala 214:29]
  wire [1:0] _GEN_711 = io_cm_0 != 6'h0 ? _GEN_647 : _GEN_583; // @[Rename.scala 214:29]
  wire [1:0] _GEN_712 = io_cm_0 != 6'h0 ? _GEN_648 : _GEN_584; // @[Rename.scala 214:29]
  wire [1:0] _GEN_713 = io_cm_0 != 6'h0 ? _GEN_649 : _GEN_585; // @[Rename.scala 214:29]
  wire [1:0] _GEN_714 = io_cm_0 != 6'h0 ? _GEN_650 : _GEN_586; // @[Rename.scala 214:29]
  wire [1:0] _GEN_715 = io_cm_0 != 6'h0 ? _GEN_651 : _GEN_587; // @[Rename.scala 214:29]
  wire [1:0] _GEN_716 = io_cm_0 != 6'h0 ? _GEN_652 : _GEN_588; // @[Rename.scala 214:29]
  wire [1:0] _GEN_717 = io_cm_0 != 6'h0 ? _GEN_653 : _GEN_589; // @[Rename.scala 214:29]
  wire [1:0] _GEN_718 = io_cm_0 != 6'h0 ? _GEN_654 : _GEN_590; // @[Rename.scala 214:29]
  wire [1:0] _GEN_719 = io_cm_0 != 6'h0 ? _GEN_655 : _GEN_591; // @[Rename.scala 214:29]
  wire [1:0] _GEN_720 = io_cm_0 != 6'h0 ? _GEN_656 : _GEN_592; // @[Rename.scala 214:29]
  wire [1:0] _GEN_721 = io_cm_0 != 6'h0 ? _GEN_657 : _GEN_593; // @[Rename.scala 214:29]
  wire [1:0] _GEN_722 = io_cm_0 != 6'h0 ? _GEN_658 : _GEN_594; // @[Rename.scala 214:29]
  wire [1:0] _GEN_723 = io_cm_0 != 6'h0 ? _GEN_659 : _GEN_595; // @[Rename.scala 214:29]
  wire [1:0] _GEN_724 = io_cm_0 != 6'h0 ? _GEN_660 : _GEN_596; // @[Rename.scala 214:29]
  wire [1:0] _GEN_725 = io_cm_0 != 6'h0 ? _GEN_661 : _GEN_597; // @[Rename.scala 214:29]
  wire [1:0] _GEN_726 = io_cm_0 != 6'h0 ? _GEN_662 : _GEN_598; // @[Rename.scala 214:29]
  wire [1:0] _GEN_727 = io_cm_0 != 6'h0 ? _GEN_663 : _GEN_599; // @[Rename.scala 214:29]
  wire [1:0] _GEN_728 = io_cm_0 != 6'h0 ? _GEN_664 : _GEN_600; // @[Rename.scala 214:29]
  wire [1:0] _GEN_729 = io_cm_0 != 6'h0 ? _GEN_665 : _GEN_601; // @[Rename.scala 214:29]
  wire [1:0] _GEN_730 = io_cm_0 != 6'h0 ? _GEN_666 : _GEN_602; // @[Rename.scala 214:29]
  wire [1:0] _GEN_731 = io_cm_0 != 6'h0 ? _GEN_667 : _GEN_603; // @[Rename.scala 214:29]
  wire [1:0] _GEN_732 = io_cm_0 != 6'h0 ? _GEN_668 : _GEN_604; // @[Rename.scala 214:29]
  wire [1:0] _GEN_733 = io_cm_0 != 6'h0 ? _GEN_669 : _GEN_605; // @[Rename.scala 214:29]
  wire [1:0] _GEN_734 = io_cm_0 != 6'h0 ? _GEN_670 : _GEN_606; // @[Rename.scala 214:29]
  wire [1:0] _GEN_735 = io_cm_0 != 6'h0 ? _GEN_671 : _GEN_607; // @[Rename.scala 214:29]
  wire [1:0] _GEN_736 = io_cm_0 != 6'h0 ? _GEN_672 : _GEN_608; // @[Rename.scala 214:29]
  wire [1:0] _GEN_737 = io_cm_0 != 6'h0 ? _GEN_673 : _GEN_609; // @[Rename.scala 214:29]
  wire [1:0] _GEN_738 = io_cm_0 != 6'h0 ? _GEN_674 : _GEN_610; // @[Rename.scala 214:29]
  wire [1:0] _GEN_739 = io_cm_0 != 6'h0 ? _GEN_675 : _GEN_611; // @[Rename.scala 214:29]
  wire [1:0] _GEN_740 = io_cm_0 != 6'h0 ? _GEN_676 : _GEN_612; // @[Rename.scala 214:29]
  wire [1:0] _GEN_741 = io_cm_0 != 6'h0 ? _GEN_677 : _GEN_613; // @[Rename.scala 214:29]
  wire [1:0] _GEN_742 = io_cm_0 != 6'h0 ? _GEN_678 : _GEN_614; // @[Rename.scala 214:29]
  wire [1:0] _GEN_743 = io_cm_0 != 6'h0 ? _GEN_679 : _GEN_615; // @[Rename.scala 214:29]
  wire [1:0] _GEN_744 = io_cm_0 != 6'h0 ? _GEN_680 : _GEN_616; // @[Rename.scala 214:29]
  wire [1:0] _GEN_745 = io_cm_0 != 6'h0 ? _GEN_681 : _GEN_617; // @[Rename.scala 214:29]
  wire [1:0] _GEN_746 = io_cm_0 != 6'h0 ? _GEN_682 : _GEN_618; // @[Rename.scala 214:29]
  wire [1:0] _GEN_747 = io_cm_0 != 6'h0 ? _GEN_683 : _GEN_619; // @[Rename.scala 214:29]
  wire [1:0] _GEN_748 = io_cm_0 != 6'h0 ? _GEN_684 : _GEN_620; // @[Rename.scala 214:29]
  wire [1:0] _GEN_749 = io_cm_0 != 6'h0 ? _GEN_685 : _GEN_621; // @[Rename.scala 214:29]
  wire [1:0] _GEN_750 = io_cm_0 != 6'h0 ? _GEN_686 : _GEN_622; // @[Rename.scala 214:29]
  wire [1:0] _GEN_751 = io_cm_0 != 6'h0 ? _GEN_687 : _GEN_623; // @[Rename.scala 214:29]
  wire [1:0] _GEN_752 = io_cm_0 != 6'h0 ? _GEN_688 : _GEN_624; // @[Rename.scala 214:29]
  wire [1:0] _GEN_753 = io_cm_0 != 6'h0 ? _GEN_689 : _GEN_625; // @[Rename.scala 214:29]
  wire [1:0] _GEN_754 = io_cm_0 != 6'h0 ? _GEN_690 : _GEN_626; // @[Rename.scala 214:29]
  wire [1:0] _GEN_755 = io_cm_0 != 6'h0 ? _GEN_691 : _GEN_627; // @[Rename.scala 214:29]
  wire [1:0] _GEN_756 = io_cm_0 != 6'h0 ? _GEN_692 : _GEN_628; // @[Rename.scala 214:29]
  wire [1:0] _GEN_757 = io_cm_0 != 6'h0 ? _GEN_693 : _GEN_629; // @[Rename.scala 214:29]
  wire [1:0] _GEN_758 = io_cm_0 != 6'h0 ? _GEN_694 : _GEN_630; // @[Rename.scala 214:29]
  wire [1:0] _GEN_759 = io_cm_0 != 6'h0 ? _GEN_695 : _GEN_631; // @[Rename.scala 214:29]
  wire [1:0] _GEN_760 = io_cm_0 != 6'h0 ? _GEN_696 : _GEN_632; // @[Rename.scala 214:29]
  wire [1:0] _GEN_761 = io_cm_0 != 6'h0 ? _GEN_697 : _GEN_633; // @[Rename.scala 214:29]
  wire [1:0] _GEN_762 = io_cm_0 != 6'h0 ? _GEN_698 : _GEN_634; // @[Rename.scala 214:29]
  wire [1:0] _GEN_763 = io_cm_0 != 6'h0 ? _GEN_699 : _GEN_635; // @[Rename.scala 214:29]
  wire [1:0] _GEN_764 = io_cm_0 != 6'h0 ? _GEN_700 : _GEN_636; // @[Rename.scala 214:29]
  wire [1:0] _GEN_765 = io_cm_0 != 6'h0 ? _GEN_701 : _GEN_637; // @[Rename.scala 214:29]
  wire [1:0] _GEN_766 = io_cm_0 != 6'h0 ? _GEN_702 : _GEN_638; // @[Rename.scala 214:29]
  wire [1:0] _GEN_767 = io_cm_0 != 6'h0 ? _GEN_703 : _GEN_639; // @[Rename.scala 214:29]
  wire [1:0] _GEN_769 = 6'h1 == io_cm_1 ? 2'h3 : _GEN_705; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_770 = 6'h2 == io_cm_1 ? 2'h3 : _GEN_706; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_771 = 6'h3 == io_cm_1 ? 2'h3 : _GEN_707; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_772 = 6'h4 == io_cm_1 ? 2'h3 : _GEN_708; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_773 = 6'h5 == io_cm_1 ? 2'h3 : _GEN_709; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_774 = 6'h6 == io_cm_1 ? 2'h3 : _GEN_710; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_775 = 6'h7 == io_cm_1 ? 2'h3 : _GEN_711; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_776 = 6'h8 == io_cm_1 ? 2'h3 : _GEN_712; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_777 = 6'h9 == io_cm_1 ? 2'h3 : _GEN_713; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_778 = 6'ha == io_cm_1 ? 2'h3 : _GEN_714; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_779 = 6'hb == io_cm_1 ? 2'h3 : _GEN_715; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_780 = 6'hc == io_cm_1 ? 2'h3 : _GEN_716; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_781 = 6'hd == io_cm_1 ? 2'h3 : _GEN_717; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_782 = 6'he == io_cm_1 ? 2'h3 : _GEN_718; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_783 = 6'hf == io_cm_1 ? 2'h3 : _GEN_719; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_784 = 6'h10 == io_cm_1 ? 2'h3 : _GEN_720; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_785 = 6'h11 == io_cm_1 ? 2'h3 : _GEN_721; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_786 = 6'h12 == io_cm_1 ? 2'h3 : _GEN_722; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_787 = 6'h13 == io_cm_1 ? 2'h3 : _GEN_723; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_788 = 6'h14 == io_cm_1 ? 2'h3 : _GEN_724; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_789 = 6'h15 == io_cm_1 ? 2'h3 : _GEN_725; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_790 = 6'h16 == io_cm_1 ? 2'h3 : _GEN_726; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_791 = 6'h17 == io_cm_1 ? 2'h3 : _GEN_727; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_792 = 6'h18 == io_cm_1 ? 2'h3 : _GEN_728; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_793 = 6'h19 == io_cm_1 ? 2'h3 : _GEN_729; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_794 = 6'h1a == io_cm_1 ? 2'h3 : _GEN_730; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_795 = 6'h1b == io_cm_1 ? 2'h3 : _GEN_731; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_796 = 6'h1c == io_cm_1 ? 2'h3 : _GEN_732; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_797 = 6'h1d == io_cm_1 ? 2'h3 : _GEN_733; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_798 = 6'h1e == io_cm_1 ? 2'h3 : _GEN_734; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_799 = 6'h1f == io_cm_1 ? 2'h3 : _GEN_735; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_800 = 6'h20 == io_cm_1 ? 2'h3 : _GEN_736; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_801 = 6'h21 == io_cm_1 ? 2'h3 : _GEN_737; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_802 = 6'h22 == io_cm_1 ? 2'h3 : _GEN_738; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_803 = 6'h23 == io_cm_1 ? 2'h3 : _GEN_739; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_804 = 6'h24 == io_cm_1 ? 2'h3 : _GEN_740; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_805 = 6'h25 == io_cm_1 ? 2'h3 : _GEN_741; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_806 = 6'h26 == io_cm_1 ? 2'h3 : _GEN_742; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_807 = 6'h27 == io_cm_1 ? 2'h3 : _GEN_743; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_808 = 6'h28 == io_cm_1 ? 2'h3 : _GEN_744; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_809 = 6'h29 == io_cm_1 ? 2'h3 : _GEN_745; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_810 = 6'h2a == io_cm_1 ? 2'h3 : _GEN_746; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_811 = 6'h2b == io_cm_1 ? 2'h3 : _GEN_747; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_812 = 6'h2c == io_cm_1 ? 2'h3 : _GEN_748; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_813 = 6'h2d == io_cm_1 ? 2'h3 : _GEN_749; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_814 = 6'h2e == io_cm_1 ? 2'h3 : _GEN_750; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_815 = 6'h2f == io_cm_1 ? 2'h3 : _GEN_751; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_816 = 6'h30 == io_cm_1 ? 2'h3 : _GEN_752; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_817 = 6'h31 == io_cm_1 ? 2'h3 : _GEN_753; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_818 = 6'h32 == io_cm_1 ? 2'h3 : _GEN_754; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_819 = 6'h33 == io_cm_1 ? 2'h3 : _GEN_755; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_820 = 6'h34 == io_cm_1 ? 2'h3 : _GEN_756; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_821 = 6'h35 == io_cm_1 ? 2'h3 : _GEN_757; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_822 = 6'h36 == io_cm_1 ? 2'h3 : _GEN_758; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_823 = 6'h37 == io_cm_1 ? 2'h3 : _GEN_759; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_824 = 6'h38 == io_cm_1 ? 2'h3 : _GEN_760; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_825 = 6'h39 == io_cm_1 ? 2'h3 : _GEN_761; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_826 = 6'h3a == io_cm_1 ? 2'h3 : _GEN_762; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_827 = 6'h3b == io_cm_1 ? 2'h3 : _GEN_763; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_828 = 6'h3c == io_cm_1 ? 2'h3 : _GEN_764; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_829 = 6'h3d == io_cm_1 ? 2'h3 : _GEN_765; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_830 = 6'h3e == io_cm_1 ? 2'h3 : _GEN_766; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_831 = 6'h3f == io_cm_1 ? 2'h3 : _GEN_767; // @[Rename.scala 215:{23,23}]
  wire [1:0] _GEN_833 = io_cm_1 != 6'h0 ? _GEN_769 : _GEN_705; // @[Rename.scala 214:29]
  wire [1:0] _GEN_834 = io_cm_1 != 6'h0 ? _GEN_770 : _GEN_706; // @[Rename.scala 214:29]
  wire [1:0] _GEN_835 = io_cm_1 != 6'h0 ? _GEN_771 : _GEN_707; // @[Rename.scala 214:29]
  wire [1:0] _GEN_836 = io_cm_1 != 6'h0 ? _GEN_772 : _GEN_708; // @[Rename.scala 214:29]
  wire [1:0] _GEN_837 = io_cm_1 != 6'h0 ? _GEN_773 : _GEN_709; // @[Rename.scala 214:29]
  wire [1:0] _GEN_838 = io_cm_1 != 6'h0 ? _GEN_774 : _GEN_710; // @[Rename.scala 214:29]
  wire [1:0] _GEN_839 = io_cm_1 != 6'h0 ? _GEN_775 : _GEN_711; // @[Rename.scala 214:29]
  wire [1:0] _GEN_840 = io_cm_1 != 6'h0 ? _GEN_776 : _GEN_712; // @[Rename.scala 214:29]
  wire [1:0] _GEN_841 = io_cm_1 != 6'h0 ? _GEN_777 : _GEN_713; // @[Rename.scala 214:29]
  wire [1:0] _GEN_842 = io_cm_1 != 6'h0 ? _GEN_778 : _GEN_714; // @[Rename.scala 214:29]
  wire [1:0] _GEN_843 = io_cm_1 != 6'h0 ? _GEN_779 : _GEN_715; // @[Rename.scala 214:29]
  wire [1:0] _GEN_844 = io_cm_1 != 6'h0 ? _GEN_780 : _GEN_716; // @[Rename.scala 214:29]
  wire [1:0] _GEN_845 = io_cm_1 != 6'h0 ? _GEN_781 : _GEN_717; // @[Rename.scala 214:29]
  wire [1:0] _GEN_846 = io_cm_1 != 6'h0 ? _GEN_782 : _GEN_718; // @[Rename.scala 214:29]
  wire [1:0] _GEN_847 = io_cm_1 != 6'h0 ? _GEN_783 : _GEN_719; // @[Rename.scala 214:29]
  wire [1:0] _GEN_848 = io_cm_1 != 6'h0 ? _GEN_784 : _GEN_720; // @[Rename.scala 214:29]
  wire [1:0] _GEN_849 = io_cm_1 != 6'h0 ? _GEN_785 : _GEN_721; // @[Rename.scala 214:29]
  wire [1:0] _GEN_850 = io_cm_1 != 6'h0 ? _GEN_786 : _GEN_722; // @[Rename.scala 214:29]
  wire [1:0] _GEN_851 = io_cm_1 != 6'h0 ? _GEN_787 : _GEN_723; // @[Rename.scala 214:29]
  wire [1:0] _GEN_852 = io_cm_1 != 6'h0 ? _GEN_788 : _GEN_724; // @[Rename.scala 214:29]
  wire [1:0] _GEN_853 = io_cm_1 != 6'h0 ? _GEN_789 : _GEN_725; // @[Rename.scala 214:29]
  wire [1:0] _GEN_854 = io_cm_1 != 6'h0 ? _GEN_790 : _GEN_726; // @[Rename.scala 214:29]
  wire [1:0] _GEN_855 = io_cm_1 != 6'h0 ? _GEN_791 : _GEN_727; // @[Rename.scala 214:29]
  wire [1:0] _GEN_856 = io_cm_1 != 6'h0 ? _GEN_792 : _GEN_728; // @[Rename.scala 214:29]
  wire [1:0] _GEN_857 = io_cm_1 != 6'h0 ? _GEN_793 : _GEN_729; // @[Rename.scala 214:29]
  wire [1:0] _GEN_858 = io_cm_1 != 6'h0 ? _GEN_794 : _GEN_730; // @[Rename.scala 214:29]
  wire [1:0] _GEN_859 = io_cm_1 != 6'h0 ? _GEN_795 : _GEN_731; // @[Rename.scala 214:29]
  wire [1:0] _GEN_860 = io_cm_1 != 6'h0 ? _GEN_796 : _GEN_732; // @[Rename.scala 214:29]
  wire [1:0] _GEN_861 = io_cm_1 != 6'h0 ? _GEN_797 : _GEN_733; // @[Rename.scala 214:29]
  wire [1:0] _GEN_862 = io_cm_1 != 6'h0 ? _GEN_798 : _GEN_734; // @[Rename.scala 214:29]
  wire [1:0] _GEN_863 = io_cm_1 != 6'h0 ? _GEN_799 : _GEN_735; // @[Rename.scala 214:29]
  wire [1:0] _GEN_864 = io_cm_1 != 6'h0 ? _GEN_800 : _GEN_736; // @[Rename.scala 214:29]
  wire [1:0] _GEN_865 = io_cm_1 != 6'h0 ? _GEN_801 : _GEN_737; // @[Rename.scala 214:29]
  wire [1:0] _GEN_866 = io_cm_1 != 6'h0 ? _GEN_802 : _GEN_738; // @[Rename.scala 214:29]
  wire [1:0] _GEN_867 = io_cm_1 != 6'h0 ? _GEN_803 : _GEN_739; // @[Rename.scala 214:29]
  wire [1:0] _GEN_868 = io_cm_1 != 6'h0 ? _GEN_804 : _GEN_740; // @[Rename.scala 214:29]
  wire [1:0] _GEN_869 = io_cm_1 != 6'h0 ? _GEN_805 : _GEN_741; // @[Rename.scala 214:29]
  wire [1:0] _GEN_870 = io_cm_1 != 6'h0 ? _GEN_806 : _GEN_742; // @[Rename.scala 214:29]
  wire [1:0] _GEN_871 = io_cm_1 != 6'h0 ? _GEN_807 : _GEN_743; // @[Rename.scala 214:29]
  wire [1:0] _GEN_872 = io_cm_1 != 6'h0 ? _GEN_808 : _GEN_744; // @[Rename.scala 214:29]
  wire [1:0] _GEN_873 = io_cm_1 != 6'h0 ? _GEN_809 : _GEN_745; // @[Rename.scala 214:29]
  wire [1:0] _GEN_874 = io_cm_1 != 6'h0 ? _GEN_810 : _GEN_746; // @[Rename.scala 214:29]
  wire [1:0] _GEN_875 = io_cm_1 != 6'h0 ? _GEN_811 : _GEN_747; // @[Rename.scala 214:29]
  wire [1:0] _GEN_876 = io_cm_1 != 6'h0 ? _GEN_812 : _GEN_748; // @[Rename.scala 214:29]
  wire [1:0] _GEN_877 = io_cm_1 != 6'h0 ? _GEN_813 : _GEN_749; // @[Rename.scala 214:29]
  wire [1:0] _GEN_878 = io_cm_1 != 6'h0 ? _GEN_814 : _GEN_750; // @[Rename.scala 214:29]
  wire [1:0] _GEN_879 = io_cm_1 != 6'h0 ? _GEN_815 : _GEN_751; // @[Rename.scala 214:29]
  wire [1:0] _GEN_880 = io_cm_1 != 6'h0 ? _GEN_816 : _GEN_752; // @[Rename.scala 214:29]
  wire [1:0] _GEN_881 = io_cm_1 != 6'h0 ? _GEN_817 : _GEN_753; // @[Rename.scala 214:29]
  wire [1:0] _GEN_882 = io_cm_1 != 6'h0 ? _GEN_818 : _GEN_754; // @[Rename.scala 214:29]
  wire [1:0] _GEN_883 = io_cm_1 != 6'h0 ? _GEN_819 : _GEN_755; // @[Rename.scala 214:29]
  wire [1:0] _GEN_884 = io_cm_1 != 6'h0 ? _GEN_820 : _GEN_756; // @[Rename.scala 214:29]
  wire [1:0] _GEN_885 = io_cm_1 != 6'h0 ? _GEN_821 : _GEN_757; // @[Rename.scala 214:29]
  wire [1:0] _GEN_886 = io_cm_1 != 6'h0 ? _GEN_822 : _GEN_758; // @[Rename.scala 214:29]
  wire [1:0] _GEN_887 = io_cm_1 != 6'h0 ? _GEN_823 : _GEN_759; // @[Rename.scala 214:29]
  wire [1:0] _GEN_888 = io_cm_1 != 6'h0 ? _GEN_824 : _GEN_760; // @[Rename.scala 214:29]
  wire [1:0] _GEN_889 = io_cm_1 != 6'h0 ? _GEN_825 : _GEN_761; // @[Rename.scala 214:29]
  wire [1:0] _GEN_890 = io_cm_1 != 6'h0 ? _GEN_826 : _GEN_762; // @[Rename.scala 214:29]
  wire [1:0] _GEN_891 = io_cm_1 != 6'h0 ? _GEN_827 : _GEN_763; // @[Rename.scala 214:29]
  wire [1:0] _GEN_892 = io_cm_1 != 6'h0 ? _GEN_828 : _GEN_764; // @[Rename.scala 214:29]
  wire [1:0] _GEN_893 = io_cm_1 != 6'h0 ? _GEN_829 : _GEN_765; // @[Rename.scala 214:29]
  wire [1:0] _GEN_894 = io_cm_1 != 6'h0 ? _GEN_830 : _GEN_766; // @[Rename.scala 214:29]
  wire [1:0] _GEN_895 = io_cm_1 != 6'h0 ? _GEN_831 : _GEN_767; // @[Rename.scala 214:29]
  wire [1:0] _GEN_897 = 6'h1 == io_free_0 ? 2'h0 : _GEN_833; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_898 = 6'h2 == io_free_0 ? 2'h0 : _GEN_834; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_899 = 6'h3 == io_free_0 ? 2'h0 : _GEN_835; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_900 = 6'h4 == io_free_0 ? 2'h0 : _GEN_836; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_901 = 6'h5 == io_free_0 ? 2'h0 : _GEN_837; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_902 = 6'h6 == io_free_0 ? 2'h0 : _GEN_838; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_903 = 6'h7 == io_free_0 ? 2'h0 : _GEN_839; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_904 = 6'h8 == io_free_0 ? 2'h0 : _GEN_840; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_905 = 6'h9 == io_free_0 ? 2'h0 : _GEN_841; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_906 = 6'ha == io_free_0 ? 2'h0 : _GEN_842; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_907 = 6'hb == io_free_0 ? 2'h0 : _GEN_843; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_908 = 6'hc == io_free_0 ? 2'h0 : _GEN_844; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_909 = 6'hd == io_free_0 ? 2'h0 : _GEN_845; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_910 = 6'he == io_free_0 ? 2'h0 : _GEN_846; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_911 = 6'hf == io_free_0 ? 2'h0 : _GEN_847; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_912 = 6'h10 == io_free_0 ? 2'h0 : _GEN_848; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_913 = 6'h11 == io_free_0 ? 2'h0 : _GEN_849; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_914 = 6'h12 == io_free_0 ? 2'h0 : _GEN_850; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_915 = 6'h13 == io_free_0 ? 2'h0 : _GEN_851; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_916 = 6'h14 == io_free_0 ? 2'h0 : _GEN_852; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_917 = 6'h15 == io_free_0 ? 2'h0 : _GEN_853; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_918 = 6'h16 == io_free_0 ? 2'h0 : _GEN_854; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_919 = 6'h17 == io_free_0 ? 2'h0 : _GEN_855; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_920 = 6'h18 == io_free_0 ? 2'h0 : _GEN_856; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_921 = 6'h19 == io_free_0 ? 2'h0 : _GEN_857; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_922 = 6'h1a == io_free_0 ? 2'h0 : _GEN_858; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_923 = 6'h1b == io_free_0 ? 2'h0 : _GEN_859; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_924 = 6'h1c == io_free_0 ? 2'h0 : _GEN_860; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_925 = 6'h1d == io_free_0 ? 2'h0 : _GEN_861; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_926 = 6'h1e == io_free_0 ? 2'h0 : _GEN_862; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_927 = 6'h1f == io_free_0 ? 2'h0 : _GEN_863; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_928 = 6'h20 == io_free_0 ? 2'h0 : _GEN_864; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_929 = 6'h21 == io_free_0 ? 2'h0 : _GEN_865; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_930 = 6'h22 == io_free_0 ? 2'h0 : _GEN_866; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_931 = 6'h23 == io_free_0 ? 2'h0 : _GEN_867; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_932 = 6'h24 == io_free_0 ? 2'h0 : _GEN_868; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_933 = 6'h25 == io_free_0 ? 2'h0 : _GEN_869; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_934 = 6'h26 == io_free_0 ? 2'h0 : _GEN_870; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_935 = 6'h27 == io_free_0 ? 2'h0 : _GEN_871; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_936 = 6'h28 == io_free_0 ? 2'h0 : _GEN_872; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_937 = 6'h29 == io_free_0 ? 2'h0 : _GEN_873; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_938 = 6'h2a == io_free_0 ? 2'h0 : _GEN_874; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_939 = 6'h2b == io_free_0 ? 2'h0 : _GEN_875; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_940 = 6'h2c == io_free_0 ? 2'h0 : _GEN_876; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_941 = 6'h2d == io_free_0 ? 2'h0 : _GEN_877; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_942 = 6'h2e == io_free_0 ? 2'h0 : _GEN_878; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_943 = 6'h2f == io_free_0 ? 2'h0 : _GEN_879; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_944 = 6'h30 == io_free_0 ? 2'h0 : _GEN_880; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_945 = 6'h31 == io_free_0 ? 2'h0 : _GEN_881; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_946 = 6'h32 == io_free_0 ? 2'h0 : _GEN_882; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_947 = 6'h33 == io_free_0 ? 2'h0 : _GEN_883; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_948 = 6'h34 == io_free_0 ? 2'h0 : _GEN_884; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_949 = 6'h35 == io_free_0 ? 2'h0 : _GEN_885; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_950 = 6'h36 == io_free_0 ? 2'h0 : _GEN_886; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_951 = 6'h37 == io_free_0 ? 2'h0 : _GEN_887; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_952 = 6'h38 == io_free_0 ? 2'h0 : _GEN_888; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_953 = 6'h39 == io_free_0 ? 2'h0 : _GEN_889; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_954 = 6'h3a == io_free_0 ? 2'h0 : _GEN_890; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_955 = 6'h3b == io_free_0 ? 2'h0 : _GEN_891; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_956 = 6'h3c == io_free_0 ? 2'h0 : _GEN_892; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_957 = 6'h3d == io_free_0 ? 2'h0 : _GEN_893; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_958 = 6'h3e == io_free_0 ? 2'h0 : _GEN_894; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_959 = 6'h3f == io_free_0 ? 2'h0 : _GEN_895; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_961 = io_free_0 != 6'h0 ? _GEN_897 : _GEN_833; // @[Rename.scala 220:31]
  wire [1:0] _GEN_962 = io_free_0 != 6'h0 ? _GEN_898 : _GEN_834; // @[Rename.scala 220:31]
  wire [1:0] _GEN_963 = io_free_0 != 6'h0 ? _GEN_899 : _GEN_835; // @[Rename.scala 220:31]
  wire [1:0] _GEN_964 = io_free_0 != 6'h0 ? _GEN_900 : _GEN_836; // @[Rename.scala 220:31]
  wire [1:0] _GEN_965 = io_free_0 != 6'h0 ? _GEN_901 : _GEN_837; // @[Rename.scala 220:31]
  wire [1:0] _GEN_966 = io_free_0 != 6'h0 ? _GEN_902 : _GEN_838; // @[Rename.scala 220:31]
  wire [1:0] _GEN_967 = io_free_0 != 6'h0 ? _GEN_903 : _GEN_839; // @[Rename.scala 220:31]
  wire [1:0] _GEN_968 = io_free_0 != 6'h0 ? _GEN_904 : _GEN_840; // @[Rename.scala 220:31]
  wire [1:0] _GEN_969 = io_free_0 != 6'h0 ? _GEN_905 : _GEN_841; // @[Rename.scala 220:31]
  wire [1:0] _GEN_970 = io_free_0 != 6'h0 ? _GEN_906 : _GEN_842; // @[Rename.scala 220:31]
  wire [1:0] _GEN_971 = io_free_0 != 6'h0 ? _GEN_907 : _GEN_843; // @[Rename.scala 220:31]
  wire [1:0] _GEN_972 = io_free_0 != 6'h0 ? _GEN_908 : _GEN_844; // @[Rename.scala 220:31]
  wire [1:0] _GEN_973 = io_free_0 != 6'h0 ? _GEN_909 : _GEN_845; // @[Rename.scala 220:31]
  wire [1:0] _GEN_974 = io_free_0 != 6'h0 ? _GEN_910 : _GEN_846; // @[Rename.scala 220:31]
  wire [1:0] _GEN_975 = io_free_0 != 6'h0 ? _GEN_911 : _GEN_847; // @[Rename.scala 220:31]
  wire [1:0] _GEN_976 = io_free_0 != 6'h0 ? _GEN_912 : _GEN_848; // @[Rename.scala 220:31]
  wire [1:0] _GEN_977 = io_free_0 != 6'h0 ? _GEN_913 : _GEN_849; // @[Rename.scala 220:31]
  wire [1:0] _GEN_978 = io_free_0 != 6'h0 ? _GEN_914 : _GEN_850; // @[Rename.scala 220:31]
  wire [1:0] _GEN_979 = io_free_0 != 6'h0 ? _GEN_915 : _GEN_851; // @[Rename.scala 220:31]
  wire [1:0] _GEN_980 = io_free_0 != 6'h0 ? _GEN_916 : _GEN_852; // @[Rename.scala 220:31]
  wire [1:0] _GEN_981 = io_free_0 != 6'h0 ? _GEN_917 : _GEN_853; // @[Rename.scala 220:31]
  wire [1:0] _GEN_982 = io_free_0 != 6'h0 ? _GEN_918 : _GEN_854; // @[Rename.scala 220:31]
  wire [1:0] _GEN_983 = io_free_0 != 6'h0 ? _GEN_919 : _GEN_855; // @[Rename.scala 220:31]
  wire [1:0] _GEN_984 = io_free_0 != 6'h0 ? _GEN_920 : _GEN_856; // @[Rename.scala 220:31]
  wire [1:0] _GEN_985 = io_free_0 != 6'h0 ? _GEN_921 : _GEN_857; // @[Rename.scala 220:31]
  wire [1:0] _GEN_986 = io_free_0 != 6'h0 ? _GEN_922 : _GEN_858; // @[Rename.scala 220:31]
  wire [1:0] _GEN_987 = io_free_0 != 6'h0 ? _GEN_923 : _GEN_859; // @[Rename.scala 220:31]
  wire [1:0] _GEN_988 = io_free_0 != 6'h0 ? _GEN_924 : _GEN_860; // @[Rename.scala 220:31]
  wire [1:0] _GEN_989 = io_free_0 != 6'h0 ? _GEN_925 : _GEN_861; // @[Rename.scala 220:31]
  wire [1:0] _GEN_990 = io_free_0 != 6'h0 ? _GEN_926 : _GEN_862; // @[Rename.scala 220:31]
  wire [1:0] _GEN_991 = io_free_0 != 6'h0 ? _GEN_927 : _GEN_863; // @[Rename.scala 220:31]
  wire [1:0] _GEN_992 = io_free_0 != 6'h0 ? _GEN_928 : _GEN_864; // @[Rename.scala 220:31]
  wire [1:0] _GEN_993 = io_free_0 != 6'h0 ? _GEN_929 : _GEN_865; // @[Rename.scala 220:31]
  wire [1:0] _GEN_994 = io_free_0 != 6'h0 ? _GEN_930 : _GEN_866; // @[Rename.scala 220:31]
  wire [1:0] _GEN_995 = io_free_0 != 6'h0 ? _GEN_931 : _GEN_867; // @[Rename.scala 220:31]
  wire [1:0] _GEN_996 = io_free_0 != 6'h0 ? _GEN_932 : _GEN_868; // @[Rename.scala 220:31]
  wire [1:0] _GEN_997 = io_free_0 != 6'h0 ? _GEN_933 : _GEN_869; // @[Rename.scala 220:31]
  wire [1:0] _GEN_998 = io_free_0 != 6'h0 ? _GEN_934 : _GEN_870; // @[Rename.scala 220:31]
  wire [1:0] _GEN_999 = io_free_0 != 6'h0 ? _GEN_935 : _GEN_871; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1000 = io_free_0 != 6'h0 ? _GEN_936 : _GEN_872; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1001 = io_free_0 != 6'h0 ? _GEN_937 : _GEN_873; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1002 = io_free_0 != 6'h0 ? _GEN_938 : _GEN_874; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1003 = io_free_0 != 6'h0 ? _GEN_939 : _GEN_875; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1004 = io_free_0 != 6'h0 ? _GEN_940 : _GEN_876; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1005 = io_free_0 != 6'h0 ? _GEN_941 : _GEN_877; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1006 = io_free_0 != 6'h0 ? _GEN_942 : _GEN_878; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1007 = io_free_0 != 6'h0 ? _GEN_943 : _GEN_879; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1008 = io_free_0 != 6'h0 ? _GEN_944 : _GEN_880; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1009 = io_free_0 != 6'h0 ? _GEN_945 : _GEN_881; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1010 = io_free_0 != 6'h0 ? _GEN_946 : _GEN_882; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1011 = io_free_0 != 6'h0 ? _GEN_947 : _GEN_883; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1012 = io_free_0 != 6'h0 ? _GEN_948 : _GEN_884; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1013 = io_free_0 != 6'h0 ? _GEN_949 : _GEN_885; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1014 = io_free_0 != 6'h0 ? _GEN_950 : _GEN_886; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1015 = io_free_0 != 6'h0 ? _GEN_951 : _GEN_887; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1016 = io_free_0 != 6'h0 ? _GEN_952 : _GEN_888; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1017 = io_free_0 != 6'h0 ? _GEN_953 : _GEN_889; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1018 = io_free_0 != 6'h0 ? _GEN_954 : _GEN_890; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1019 = io_free_0 != 6'h0 ? _GEN_955 : _GEN_891; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1020 = io_free_0 != 6'h0 ? _GEN_956 : _GEN_892; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1021 = io_free_0 != 6'h0 ? _GEN_957 : _GEN_893; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1022 = io_free_0 != 6'h0 ? _GEN_958 : _GEN_894; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1023 = io_free_0 != 6'h0 ? _GEN_959 : _GEN_895; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1025 = 6'h1 == io_free_1 ? 2'h0 : _GEN_961; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1026 = 6'h2 == io_free_1 ? 2'h0 : _GEN_962; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1027 = 6'h3 == io_free_1 ? 2'h0 : _GEN_963; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1028 = 6'h4 == io_free_1 ? 2'h0 : _GEN_964; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1029 = 6'h5 == io_free_1 ? 2'h0 : _GEN_965; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1030 = 6'h6 == io_free_1 ? 2'h0 : _GEN_966; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1031 = 6'h7 == io_free_1 ? 2'h0 : _GEN_967; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1032 = 6'h8 == io_free_1 ? 2'h0 : _GEN_968; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1033 = 6'h9 == io_free_1 ? 2'h0 : _GEN_969; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1034 = 6'ha == io_free_1 ? 2'h0 : _GEN_970; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1035 = 6'hb == io_free_1 ? 2'h0 : _GEN_971; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1036 = 6'hc == io_free_1 ? 2'h0 : _GEN_972; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1037 = 6'hd == io_free_1 ? 2'h0 : _GEN_973; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1038 = 6'he == io_free_1 ? 2'h0 : _GEN_974; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1039 = 6'hf == io_free_1 ? 2'h0 : _GEN_975; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1040 = 6'h10 == io_free_1 ? 2'h0 : _GEN_976; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1041 = 6'h11 == io_free_1 ? 2'h0 : _GEN_977; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1042 = 6'h12 == io_free_1 ? 2'h0 : _GEN_978; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1043 = 6'h13 == io_free_1 ? 2'h0 : _GEN_979; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1044 = 6'h14 == io_free_1 ? 2'h0 : _GEN_980; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1045 = 6'h15 == io_free_1 ? 2'h0 : _GEN_981; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1046 = 6'h16 == io_free_1 ? 2'h0 : _GEN_982; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1047 = 6'h17 == io_free_1 ? 2'h0 : _GEN_983; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1048 = 6'h18 == io_free_1 ? 2'h0 : _GEN_984; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1049 = 6'h19 == io_free_1 ? 2'h0 : _GEN_985; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1050 = 6'h1a == io_free_1 ? 2'h0 : _GEN_986; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1051 = 6'h1b == io_free_1 ? 2'h0 : _GEN_987; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1052 = 6'h1c == io_free_1 ? 2'h0 : _GEN_988; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1053 = 6'h1d == io_free_1 ? 2'h0 : _GEN_989; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1054 = 6'h1e == io_free_1 ? 2'h0 : _GEN_990; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1055 = 6'h1f == io_free_1 ? 2'h0 : _GEN_991; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1056 = 6'h20 == io_free_1 ? 2'h0 : _GEN_992; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1057 = 6'h21 == io_free_1 ? 2'h0 : _GEN_993; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1058 = 6'h22 == io_free_1 ? 2'h0 : _GEN_994; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1059 = 6'h23 == io_free_1 ? 2'h0 : _GEN_995; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1060 = 6'h24 == io_free_1 ? 2'h0 : _GEN_996; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1061 = 6'h25 == io_free_1 ? 2'h0 : _GEN_997; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1062 = 6'h26 == io_free_1 ? 2'h0 : _GEN_998; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1063 = 6'h27 == io_free_1 ? 2'h0 : _GEN_999; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1064 = 6'h28 == io_free_1 ? 2'h0 : _GEN_1000; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1065 = 6'h29 == io_free_1 ? 2'h0 : _GEN_1001; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1066 = 6'h2a == io_free_1 ? 2'h0 : _GEN_1002; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1067 = 6'h2b == io_free_1 ? 2'h0 : _GEN_1003; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1068 = 6'h2c == io_free_1 ? 2'h0 : _GEN_1004; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1069 = 6'h2d == io_free_1 ? 2'h0 : _GEN_1005; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1070 = 6'h2e == io_free_1 ? 2'h0 : _GEN_1006; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1071 = 6'h2f == io_free_1 ? 2'h0 : _GEN_1007; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1072 = 6'h30 == io_free_1 ? 2'h0 : _GEN_1008; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1073 = 6'h31 == io_free_1 ? 2'h0 : _GEN_1009; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1074 = 6'h32 == io_free_1 ? 2'h0 : _GEN_1010; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1075 = 6'h33 == io_free_1 ? 2'h0 : _GEN_1011; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1076 = 6'h34 == io_free_1 ? 2'h0 : _GEN_1012; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1077 = 6'h35 == io_free_1 ? 2'h0 : _GEN_1013; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1078 = 6'h36 == io_free_1 ? 2'h0 : _GEN_1014; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1079 = 6'h37 == io_free_1 ? 2'h0 : _GEN_1015; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1080 = 6'h38 == io_free_1 ? 2'h0 : _GEN_1016; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1081 = 6'h39 == io_free_1 ? 2'h0 : _GEN_1017; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1082 = 6'h3a == io_free_1 ? 2'h0 : _GEN_1018; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1083 = 6'h3b == io_free_1 ? 2'h0 : _GEN_1019; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1084 = 6'h3c == io_free_1 ? 2'h0 : _GEN_1020; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1085 = 6'h3d == io_free_1 ? 2'h0 : _GEN_1021; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1086 = 6'h3e == io_free_1 ? 2'h0 : _GEN_1022; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1087 = 6'h3f == io_free_1 ? 2'h0 : _GEN_1023; // @[Rename.scala 221:{25,25}]
  wire [1:0] _GEN_1089 = io_free_1 != 6'h0 ? _GEN_1025 : _GEN_961; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1090 = io_free_1 != 6'h0 ? _GEN_1026 : _GEN_962; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1091 = io_free_1 != 6'h0 ? _GEN_1027 : _GEN_963; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1092 = io_free_1 != 6'h0 ? _GEN_1028 : _GEN_964; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1093 = io_free_1 != 6'h0 ? _GEN_1029 : _GEN_965; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1094 = io_free_1 != 6'h0 ? _GEN_1030 : _GEN_966; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1095 = io_free_1 != 6'h0 ? _GEN_1031 : _GEN_967; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1096 = io_free_1 != 6'h0 ? _GEN_1032 : _GEN_968; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1097 = io_free_1 != 6'h0 ? _GEN_1033 : _GEN_969; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1098 = io_free_1 != 6'h0 ? _GEN_1034 : _GEN_970; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1099 = io_free_1 != 6'h0 ? _GEN_1035 : _GEN_971; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1100 = io_free_1 != 6'h0 ? _GEN_1036 : _GEN_972; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1101 = io_free_1 != 6'h0 ? _GEN_1037 : _GEN_973; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1102 = io_free_1 != 6'h0 ? _GEN_1038 : _GEN_974; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1103 = io_free_1 != 6'h0 ? _GEN_1039 : _GEN_975; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1104 = io_free_1 != 6'h0 ? _GEN_1040 : _GEN_976; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1105 = io_free_1 != 6'h0 ? _GEN_1041 : _GEN_977; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1106 = io_free_1 != 6'h0 ? _GEN_1042 : _GEN_978; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1107 = io_free_1 != 6'h0 ? _GEN_1043 : _GEN_979; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1108 = io_free_1 != 6'h0 ? _GEN_1044 : _GEN_980; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1109 = io_free_1 != 6'h0 ? _GEN_1045 : _GEN_981; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1110 = io_free_1 != 6'h0 ? _GEN_1046 : _GEN_982; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1111 = io_free_1 != 6'h0 ? _GEN_1047 : _GEN_983; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1112 = io_free_1 != 6'h0 ? _GEN_1048 : _GEN_984; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1113 = io_free_1 != 6'h0 ? _GEN_1049 : _GEN_985; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1114 = io_free_1 != 6'h0 ? _GEN_1050 : _GEN_986; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1115 = io_free_1 != 6'h0 ? _GEN_1051 : _GEN_987; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1116 = io_free_1 != 6'h0 ? _GEN_1052 : _GEN_988; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1117 = io_free_1 != 6'h0 ? _GEN_1053 : _GEN_989; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1118 = io_free_1 != 6'h0 ? _GEN_1054 : _GEN_990; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1119 = io_free_1 != 6'h0 ? _GEN_1055 : _GEN_991; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1120 = io_free_1 != 6'h0 ? _GEN_1056 : _GEN_992; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1121 = io_free_1 != 6'h0 ? _GEN_1057 : _GEN_993; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1122 = io_free_1 != 6'h0 ? _GEN_1058 : _GEN_994; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1123 = io_free_1 != 6'h0 ? _GEN_1059 : _GEN_995; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1124 = io_free_1 != 6'h0 ? _GEN_1060 : _GEN_996; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1125 = io_free_1 != 6'h0 ? _GEN_1061 : _GEN_997; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1126 = io_free_1 != 6'h0 ? _GEN_1062 : _GEN_998; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1127 = io_free_1 != 6'h0 ? _GEN_1063 : _GEN_999; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1128 = io_free_1 != 6'h0 ? _GEN_1064 : _GEN_1000; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1129 = io_free_1 != 6'h0 ? _GEN_1065 : _GEN_1001; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1130 = io_free_1 != 6'h0 ? _GEN_1066 : _GEN_1002; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1131 = io_free_1 != 6'h0 ? _GEN_1067 : _GEN_1003; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1132 = io_free_1 != 6'h0 ? _GEN_1068 : _GEN_1004; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1133 = io_free_1 != 6'h0 ? _GEN_1069 : _GEN_1005; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1134 = io_free_1 != 6'h0 ? _GEN_1070 : _GEN_1006; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1135 = io_free_1 != 6'h0 ? _GEN_1071 : _GEN_1007; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1136 = io_free_1 != 6'h0 ? _GEN_1072 : _GEN_1008; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1137 = io_free_1 != 6'h0 ? _GEN_1073 : _GEN_1009; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1138 = io_free_1 != 6'h0 ? _GEN_1074 : _GEN_1010; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1139 = io_free_1 != 6'h0 ? _GEN_1075 : _GEN_1011; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1140 = io_free_1 != 6'h0 ? _GEN_1076 : _GEN_1012; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1141 = io_free_1 != 6'h0 ? _GEN_1077 : _GEN_1013; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1142 = io_free_1 != 6'h0 ? _GEN_1078 : _GEN_1014; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1143 = io_free_1 != 6'h0 ? _GEN_1079 : _GEN_1015; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1144 = io_free_1 != 6'h0 ? _GEN_1080 : _GEN_1016; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1145 = io_free_1 != 6'h0 ? _GEN_1081 : _GEN_1017; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1146 = io_free_1 != 6'h0 ? _GEN_1082 : _GEN_1018; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1147 = io_free_1 != 6'h0 ? _GEN_1083 : _GEN_1019; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1148 = io_free_1 != 6'h0 ? _GEN_1084 : _GEN_1020; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1149 = io_free_1 != 6'h0 ? _GEN_1085 : _GEN_1021; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1150 = io_free_1 != 6'h0 ? _GEN_1086 : _GEN_1022; // @[Rename.scala 220:31]
  wire [1:0] _GEN_1151 = io_free_1 != 6'h0 ? _GEN_1087 : _GEN_1023; // @[Rename.scala 220:31]
  assign io_allocatable = free_count >= 7'h2; // @[Rename.scala 190:33]
  assign io_rd_paddr_0 = io_en & io_rd_req_0 ? _T_511 : 6'h0; // @[Rename.scala 196:24]
  assign io_rd_paddr_1 = io_en & io_rd_req_1 ? _T_643 : 6'h0; // @[Rename.scala 199:24]
  assign io_avail_list = _T_318 | _T_383; // @[Rename.scala 192:59]
  always @(posedge clock) begin
    if (reset) begin // @[Rename.scala 186:22]
      table_1 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_1 != 2'h3) begin // @[Rename.scala 227:37]
        table_1 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_1 <= _GEN_1089;
      end
    end else begin
      table_1 <= _GEN_1089;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_2 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_2 != 2'h3) begin // @[Rename.scala 227:37]
        table_2 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_2 <= _GEN_1090;
      end
    end else begin
      table_2 <= _GEN_1090;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_3 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_3 != 2'h3) begin // @[Rename.scala 227:37]
        table_3 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_3 <= _GEN_1091;
      end
    end else begin
      table_3 <= _GEN_1091;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_4 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_4 != 2'h3) begin // @[Rename.scala 227:37]
        table_4 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_4 <= _GEN_1092;
      end
    end else begin
      table_4 <= _GEN_1092;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_5 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_5 != 2'h3) begin // @[Rename.scala 227:37]
        table_5 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_5 <= _GEN_1093;
      end
    end else begin
      table_5 <= _GEN_1093;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_6 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_6 != 2'h3) begin // @[Rename.scala 227:37]
        table_6 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_6 <= _GEN_1094;
      end
    end else begin
      table_6 <= _GEN_1094;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_7 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_7 != 2'h3) begin // @[Rename.scala 227:37]
        table_7 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_7 <= _GEN_1095;
      end
    end else begin
      table_7 <= _GEN_1095;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_8 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_8 != 2'h3) begin // @[Rename.scala 227:37]
        table_8 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_8 <= _GEN_1096;
      end
    end else begin
      table_8 <= _GEN_1096;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_9 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_9 != 2'h3) begin // @[Rename.scala 227:37]
        table_9 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_9 <= _GEN_1097;
      end
    end else begin
      table_9 <= _GEN_1097;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_10 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_10 != 2'h3) begin // @[Rename.scala 227:37]
        table_10 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_10 <= _GEN_1098;
      end
    end else begin
      table_10 <= _GEN_1098;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_11 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_11 != 2'h3) begin // @[Rename.scala 227:37]
        table_11 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_11 <= _GEN_1099;
      end
    end else begin
      table_11 <= _GEN_1099;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_12 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_12 != 2'h3) begin // @[Rename.scala 227:37]
        table_12 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_12 <= _GEN_1100;
      end
    end else begin
      table_12 <= _GEN_1100;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_13 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_13 != 2'h3) begin // @[Rename.scala 227:37]
        table_13 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_13 <= _GEN_1101;
      end
    end else begin
      table_13 <= _GEN_1101;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_14 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_14 != 2'h3) begin // @[Rename.scala 227:37]
        table_14 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_14 <= _GEN_1102;
      end
    end else begin
      table_14 <= _GEN_1102;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_15 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_15 != 2'h3) begin // @[Rename.scala 227:37]
        table_15 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_15 <= _GEN_1103;
      end
    end else begin
      table_15 <= _GEN_1103;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_16 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_16 != 2'h3) begin // @[Rename.scala 227:37]
        table_16 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_16 <= _GEN_1104;
      end
    end else begin
      table_16 <= _GEN_1104;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_17 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_17 != 2'h3) begin // @[Rename.scala 227:37]
        table_17 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_17 <= _GEN_1105;
      end
    end else begin
      table_17 <= _GEN_1105;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_18 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_18 != 2'h3) begin // @[Rename.scala 227:37]
        table_18 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_18 <= _GEN_1106;
      end
    end else begin
      table_18 <= _GEN_1106;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_19 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_19 != 2'h3) begin // @[Rename.scala 227:37]
        table_19 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_19 <= _GEN_1107;
      end
    end else begin
      table_19 <= _GEN_1107;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_20 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_20 != 2'h3) begin // @[Rename.scala 227:37]
        table_20 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_20 <= _GEN_1108;
      end
    end else begin
      table_20 <= _GEN_1108;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_21 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_21 != 2'h3) begin // @[Rename.scala 227:37]
        table_21 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_21 <= _GEN_1109;
      end
    end else begin
      table_21 <= _GEN_1109;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_22 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_22 != 2'h3) begin // @[Rename.scala 227:37]
        table_22 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_22 <= _GEN_1110;
      end
    end else begin
      table_22 <= _GEN_1110;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_23 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_23 != 2'h3) begin // @[Rename.scala 227:37]
        table_23 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_23 <= _GEN_1111;
      end
    end else begin
      table_23 <= _GEN_1111;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_24 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_24 != 2'h3) begin // @[Rename.scala 227:37]
        table_24 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_24 <= _GEN_1112;
      end
    end else begin
      table_24 <= _GEN_1112;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_25 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_25 != 2'h3) begin // @[Rename.scala 227:37]
        table_25 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_25 <= _GEN_1113;
      end
    end else begin
      table_25 <= _GEN_1113;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_26 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_26 != 2'h3) begin // @[Rename.scala 227:37]
        table_26 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_26 <= _GEN_1114;
      end
    end else begin
      table_26 <= _GEN_1114;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_27 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_27 != 2'h3) begin // @[Rename.scala 227:37]
        table_27 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_27 <= _GEN_1115;
      end
    end else begin
      table_27 <= _GEN_1115;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_28 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_28 != 2'h3) begin // @[Rename.scala 227:37]
        table_28 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_28 <= _GEN_1116;
      end
    end else begin
      table_28 <= _GEN_1116;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_29 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_29 != 2'h3) begin // @[Rename.scala 227:37]
        table_29 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_29 <= _GEN_1117;
      end
    end else begin
      table_29 <= _GEN_1117;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_30 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_30 != 2'h3) begin // @[Rename.scala 227:37]
        table_30 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_30 <= _GEN_1118;
      end
    end else begin
      table_30 <= _GEN_1118;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_31 <= 2'h3; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_31 != 2'h3) begin // @[Rename.scala 227:37]
        table_31 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_31 <= _GEN_1119;
      end
    end else begin
      table_31 <= _GEN_1119;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_32 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_32 != 2'h3) begin // @[Rename.scala 227:37]
        table_32 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_32 <= _GEN_1120;
      end
    end else begin
      table_32 <= _GEN_1120;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_33 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_33 != 2'h3) begin // @[Rename.scala 227:37]
        table_33 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_33 <= _GEN_1121;
      end
    end else begin
      table_33 <= _GEN_1121;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_34 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_34 != 2'h3) begin // @[Rename.scala 227:37]
        table_34 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_34 <= _GEN_1122;
      end
    end else begin
      table_34 <= _GEN_1122;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_35 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_35 != 2'h3) begin // @[Rename.scala 227:37]
        table_35 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_35 <= _GEN_1123;
      end
    end else begin
      table_35 <= _GEN_1123;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_36 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_36 != 2'h3) begin // @[Rename.scala 227:37]
        table_36 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_36 <= _GEN_1124;
      end
    end else begin
      table_36 <= _GEN_1124;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_37 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_37 != 2'h3) begin // @[Rename.scala 227:37]
        table_37 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_37 <= _GEN_1125;
      end
    end else begin
      table_37 <= _GEN_1125;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_38 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_38 != 2'h3) begin // @[Rename.scala 227:37]
        table_38 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_38 <= _GEN_1126;
      end
    end else begin
      table_38 <= _GEN_1126;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_39 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_39 != 2'h3) begin // @[Rename.scala 227:37]
        table_39 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_39 <= _GEN_1127;
      end
    end else begin
      table_39 <= _GEN_1127;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_40 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_40 != 2'h3) begin // @[Rename.scala 227:37]
        table_40 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_40 <= _GEN_1128;
      end
    end else begin
      table_40 <= _GEN_1128;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_41 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_41 != 2'h3) begin // @[Rename.scala 227:37]
        table_41 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_41 <= _GEN_1129;
      end
    end else begin
      table_41 <= _GEN_1129;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_42 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_42 != 2'h3) begin // @[Rename.scala 227:37]
        table_42 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_42 <= _GEN_1130;
      end
    end else begin
      table_42 <= _GEN_1130;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_43 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_43 != 2'h3) begin // @[Rename.scala 227:37]
        table_43 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_43 <= _GEN_1131;
      end
    end else begin
      table_43 <= _GEN_1131;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_44 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_44 != 2'h3) begin // @[Rename.scala 227:37]
        table_44 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_44 <= _GEN_1132;
      end
    end else begin
      table_44 <= _GEN_1132;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_45 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_45 != 2'h3) begin // @[Rename.scala 227:37]
        table_45 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_45 <= _GEN_1133;
      end
    end else begin
      table_45 <= _GEN_1133;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_46 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_46 != 2'h3) begin // @[Rename.scala 227:37]
        table_46 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_46 <= _GEN_1134;
      end
    end else begin
      table_46 <= _GEN_1134;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_47 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_47 != 2'h3) begin // @[Rename.scala 227:37]
        table_47 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_47 <= _GEN_1135;
      end
    end else begin
      table_47 <= _GEN_1135;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_48 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_48 != 2'h3) begin // @[Rename.scala 227:37]
        table_48 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_48 <= _GEN_1136;
      end
    end else begin
      table_48 <= _GEN_1136;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_49 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_49 != 2'h3) begin // @[Rename.scala 227:37]
        table_49 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_49 <= _GEN_1137;
      end
    end else begin
      table_49 <= _GEN_1137;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_50 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_50 != 2'h3) begin // @[Rename.scala 227:37]
        table_50 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_50 <= _GEN_1138;
      end
    end else begin
      table_50 <= _GEN_1138;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_51 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_51 != 2'h3) begin // @[Rename.scala 227:37]
        table_51 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_51 <= _GEN_1139;
      end
    end else begin
      table_51 <= _GEN_1139;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_52 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_52 != 2'h3) begin // @[Rename.scala 227:37]
        table_52 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_52 <= _GEN_1140;
      end
    end else begin
      table_52 <= _GEN_1140;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_53 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_53 != 2'h3) begin // @[Rename.scala 227:37]
        table_53 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_53 <= _GEN_1141;
      end
    end else begin
      table_53 <= _GEN_1141;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_54 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_54 != 2'h3) begin // @[Rename.scala 227:37]
        table_54 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_54 <= _GEN_1142;
      end
    end else begin
      table_54 <= _GEN_1142;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_55 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_55 != 2'h3) begin // @[Rename.scala 227:37]
        table_55 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_55 <= _GEN_1143;
      end
    end else begin
      table_55 <= _GEN_1143;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_56 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_56 != 2'h3) begin // @[Rename.scala 227:37]
        table_56 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_56 <= _GEN_1144;
      end
    end else begin
      table_56 <= _GEN_1144;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_57 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_57 != 2'h3) begin // @[Rename.scala 227:37]
        table_57 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_57 <= _GEN_1145;
      end
    end else begin
      table_57 <= _GEN_1145;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_58 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_58 != 2'h3) begin // @[Rename.scala 227:37]
        table_58 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_58 <= _GEN_1146;
      end
    end else begin
      table_58 <= _GEN_1146;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_59 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_59 != 2'h3) begin // @[Rename.scala 227:37]
        table_59 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_59 <= _GEN_1147;
      end
    end else begin
      table_59 <= _GEN_1147;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_60 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_60 != 2'h3) begin // @[Rename.scala 227:37]
        table_60 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_60 <= _GEN_1148;
      end
    end else begin
      table_60 <= _GEN_1148;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_61 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_61 != 2'h3) begin // @[Rename.scala 227:37]
        table_61 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_61 <= _GEN_1149;
      end
    end else begin
      table_61 <= _GEN_1149;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_62 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_62 != 2'h3) begin // @[Rename.scala 227:37]
        table_62 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_62 <= _GEN_1150;
      end
    end else begin
      table_62 <= _GEN_1150;
    end
    if (reset) begin // @[Rename.scala 186:22]
      table_63 <= 2'h0; // @[Rename.scala 186:22]
    end else if (io_cm_recover) begin // @[Rename.scala 225:24]
      if (table_63 != 2'h3) begin // @[Rename.scala 227:37]
        table_63 <= 2'h0; // @[Rename.scala 228:18]
      end else begin
        table_63 <= _GEN_1151;
      end
    end else begin
      table_63 <= _GEN_1151;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  table_1 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  table_2 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  table_3 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  table_4 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  table_5 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  table_6 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  table_7 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  table_8 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  table_9 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  table_10 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  table_11 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  table_12 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  table_13 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  table_14 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  table_15 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  table_16 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  table_17 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  table_18 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  table_19 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  table_20 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  table_21 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  table_22 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  table_23 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  table_24 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  table_25 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  table_26 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  table_27 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  table_28 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  table_29 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  table_30 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  table_31 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  table_32 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  table_33 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  table_34 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  table_35 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  table_36 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  table_37 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  table_38 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  table_39 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  table_40 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  table_41 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  table_42 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  table_43 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  table_44 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  table_45 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  table_46 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  table_47 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  table_48 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  table_49 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  table_50 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  table_51 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  table_52 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  table_53 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  table_54 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  table_55 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  table_56 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  table_57 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  table_58 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  table_59 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  table_60 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  table_61 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  table_62 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  table_63 = _RAND_62[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_RenameTable(
  input        clock,
  input        reset,
  input        io_en,
  input  [4:0] io_in_0_rs1_addr,
  input  [4:0] io_in_0_rs2_addr,
  input  [4:0] io_in_1_rs1_addr,
  input  [4:0] io_in_1_rs2_addr,
  input  [4:0] io_in_1_rd_addr,
  output [5:0] io_rs1_paddr_0,
  output [5:0] io_rs1_paddr_1,
  output [5:0] io_rs2_paddr_0,
  output [5:0] io_rs2_paddr_1,
  input  [4:0] io_rd_addr_0,
  input  [4:0] io_rd_addr_1,
  output [5:0] io_rd_ppaddr_0,
  output [5:0] io_rd_ppaddr_1,
  input  [5:0] io_rd_paddr_0,
  input  [5:0] io_rd_paddr_1,
  input        io_cm_recover,
  input  [4:0] io_cm_rd_addr_0,
  input  [4:0] io_cm_rd_addr_1,
  input  [5:0] io_cm_rd_paddr_0,
  input  [5:0] io_cm_rd_paddr_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
`endif // RANDOMIZE_REG_INIT
  reg [5:0] spec_table_0; // @[Rename.scala 117:27]
  reg [5:0] spec_table_1; // @[Rename.scala 117:27]
  reg [5:0] spec_table_2; // @[Rename.scala 117:27]
  reg [5:0] spec_table_3; // @[Rename.scala 117:27]
  reg [5:0] spec_table_4; // @[Rename.scala 117:27]
  reg [5:0] spec_table_5; // @[Rename.scala 117:27]
  reg [5:0] spec_table_6; // @[Rename.scala 117:27]
  reg [5:0] spec_table_7; // @[Rename.scala 117:27]
  reg [5:0] spec_table_8; // @[Rename.scala 117:27]
  reg [5:0] spec_table_9; // @[Rename.scala 117:27]
  reg [5:0] spec_table_10; // @[Rename.scala 117:27]
  reg [5:0] spec_table_11; // @[Rename.scala 117:27]
  reg [5:0] spec_table_12; // @[Rename.scala 117:27]
  reg [5:0] spec_table_13; // @[Rename.scala 117:27]
  reg [5:0] spec_table_14; // @[Rename.scala 117:27]
  reg [5:0] spec_table_15; // @[Rename.scala 117:27]
  reg [5:0] spec_table_16; // @[Rename.scala 117:27]
  reg [5:0] spec_table_17; // @[Rename.scala 117:27]
  reg [5:0] spec_table_18; // @[Rename.scala 117:27]
  reg [5:0] spec_table_19; // @[Rename.scala 117:27]
  reg [5:0] spec_table_20; // @[Rename.scala 117:27]
  reg [5:0] spec_table_21; // @[Rename.scala 117:27]
  reg [5:0] spec_table_22; // @[Rename.scala 117:27]
  reg [5:0] spec_table_23; // @[Rename.scala 117:27]
  reg [5:0] spec_table_24; // @[Rename.scala 117:27]
  reg [5:0] spec_table_25; // @[Rename.scala 117:27]
  reg [5:0] spec_table_26; // @[Rename.scala 117:27]
  reg [5:0] spec_table_27; // @[Rename.scala 117:27]
  reg [5:0] spec_table_28; // @[Rename.scala 117:27]
  reg [5:0] spec_table_29; // @[Rename.scala 117:27]
  reg [5:0] spec_table_30; // @[Rename.scala 117:27]
  reg [5:0] spec_table_31; // @[Rename.scala 117:27]
  reg [5:0] arch_table_0; // @[Rename.scala 118:27]
  reg [5:0] arch_table_1; // @[Rename.scala 118:27]
  reg [5:0] arch_table_2; // @[Rename.scala 118:27]
  reg [5:0] arch_table_3; // @[Rename.scala 118:27]
  reg [5:0] arch_table_4; // @[Rename.scala 118:27]
  reg [5:0] arch_table_5; // @[Rename.scala 118:27]
  reg [5:0] arch_table_6; // @[Rename.scala 118:27]
  reg [5:0] arch_table_7; // @[Rename.scala 118:27]
  reg [5:0] arch_table_8; // @[Rename.scala 118:27]
  reg [5:0] arch_table_9; // @[Rename.scala 118:27]
  reg [5:0] arch_table_10; // @[Rename.scala 118:27]
  reg [5:0] arch_table_11; // @[Rename.scala 118:27]
  reg [5:0] arch_table_12; // @[Rename.scala 118:27]
  reg [5:0] arch_table_13; // @[Rename.scala 118:27]
  reg [5:0] arch_table_14; // @[Rename.scala 118:27]
  reg [5:0] arch_table_15; // @[Rename.scala 118:27]
  reg [5:0] arch_table_16; // @[Rename.scala 118:27]
  reg [5:0] arch_table_17; // @[Rename.scala 118:27]
  reg [5:0] arch_table_18; // @[Rename.scala 118:27]
  reg [5:0] arch_table_19; // @[Rename.scala 118:27]
  reg [5:0] arch_table_20; // @[Rename.scala 118:27]
  reg [5:0] arch_table_21; // @[Rename.scala 118:27]
  reg [5:0] arch_table_22; // @[Rename.scala 118:27]
  reg [5:0] arch_table_23; // @[Rename.scala 118:27]
  reg [5:0] arch_table_24; // @[Rename.scala 118:27]
  reg [5:0] arch_table_25; // @[Rename.scala 118:27]
  reg [5:0] arch_table_26; // @[Rename.scala 118:27]
  reg [5:0] arch_table_27; // @[Rename.scala 118:27]
  reg [5:0] arch_table_28; // @[Rename.scala 118:27]
  reg [5:0] arch_table_29; // @[Rename.scala 118:27]
  reg [5:0] arch_table_30; // @[Rename.scala 118:27]
  reg [5:0] arch_table_31; // @[Rename.scala 118:27]
  wire [5:0] _GEN_1 = 5'h1 == io_in_0_rs1_addr ? spec_table_1 : spec_table_0; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_2 = 5'h2 == io_in_0_rs1_addr ? spec_table_2 : _GEN_1; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_3 = 5'h3 == io_in_0_rs1_addr ? spec_table_3 : _GEN_2; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_4 = 5'h4 == io_in_0_rs1_addr ? spec_table_4 : _GEN_3; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_5 = 5'h5 == io_in_0_rs1_addr ? spec_table_5 : _GEN_4; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_6 = 5'h6 == io_in_0_rs1_addr ? spec_table_6 : _GEN_5; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_7 = 5'h7 == io_in_0_rs1_addr ? spec_table_7 : _GEN_6; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_8 = 5'h8 == io_in_0_rs1_addr ? spec_table_8 : _GEN_7; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_9 = 5'h9 == io_in_0_rs1_addr ? spec_table_9 : _GEN_8; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_10 = 5'ha == io_in_0_rs1_addr ? spec_table_10 : _GEN_9; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_11 = 5'hb == io_in_0_rs1_addr ? spec_table_11 : _GEN_10; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_12 = 5'hc == io_in_0_rs1_addr ? spec_table_12 : _GEN_11; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_13 = 5'hd == io_in_0_rs1_addr ? spec_table_13 : _GEN_12; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_14 = 5'he == io_in_0_rs1_addr ? spec_table_14 : _GEN_13; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_15 = 5'hf == io_in_0_rs1_addr ? spec_table_15 : _GEN_14; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_16 = 5'h10 == io_in_0_rs1_addr ? spec_table_16 : _GEN_15; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_17 = 5'h11 == io_in_0_rs1_addr ? spec_table_17 : _GEN_16; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_18 = 5'h12 == io_in_0_rs1_addr ? spec_table_18 : _GEN_17; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_19 = 5'h13 == io_in_0_rs1_addr ? spec_table_19 : _GEN_18; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_20 = 5'h14 == io_in_0_rs1_addr ? spec_table_20 : _GEN_19; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_21 = 5'h15 == io_in_0_rs1_addr ? spec_table_21 : _GEN_20; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_22 = 5'h16 == io_in_0_rs1_addr ? spec_table_22 : _GEN_21; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_23 = 5'h17 == io_in_0_rs1_addr ? spec_table_23 : _GEN_22; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_24 = 5'h18 == io_in_0_rs1_addr ? spec_table_24 : _GEN_23; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_25 = 5'h19 == io_in_0_rs1_addr ? spec_table_25 : _GEN_24; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_26 = 5'h1a == io_in_0_rs1_addr ? spec_table_26 : _GEN_25; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_27 = 5'h1b == io_in_0_rs1_addr ? spec_table_27 : _GEN_26; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_28 = 5'h1c == io_in_0_rs1_addr ? spec_table_28 : _GEN_27; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_29 = 5'h1d == io_in_0_rs1_addr ? spec_table_29 : _GEN_28; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_30 = 5'h1e == io_in_0_rs1_addr ? spec_table_30 : _GEN_29; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_33 = 5'h1 == io_in_0_rs2_addr ? spec_table_1 : spec_table_0; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_34 = 5'h2 == io_in_0_rs2_addr ? spec_table_2 : _GEN_33; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_35 = 5'h3 == io_in_0_rs2_addr ? spec_table_3 : _GEN_34; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_36 = 5'h4 == io_in_0_rs2_addr ? spec_table_4 : _GEN_35; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_37 = 5'h5 == io_in_0_rs2_addr ? spec_table_5 : _GEN_36; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_38 = 5'h6 == io_in_0_rs2_addr ? spec_table_6 : _GEN_37; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_39 = 5'h7 == io_in_0_rs2_addr ? spec_table_7 : _GEN_38; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_40 = 5'h8 == io_in_0_rs2_addr ? spec_table_8 : _GEN_39; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_41 = 5'h9 == io_in_0_rs2_addr ? spec_table_9 : _GEN_40; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_42 = 5'ha == io_in_0_rs2_addr ? spec_table_10 : _GEN_41; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_43 = 5'hb == io_in_0_rs2_addr ? spec_table_11 : _GEN_42; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_44 = 5'hc == io_in_0_rs2_addr ? spec_table_12 : _GEN_43; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_45 = 5'hd == io_in_0_rs2_addr ? spec_table_13 : _GEN_44; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_46 = 5'he == io_in_0_rs2_addr ? spec_table_14 : _GEN_45; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_47 = 5'hf == io_in_0_rs2_addr ? spec_table_15 : _GEN_46; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_48 = 5'h10 == io_in_0_rs2_addr ? spec_table_16 : _GEN_47; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_49 = 5'h11 == io_in_0_rs2_addr ? spec_table_17 : _GEN_48; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_50 = 5'h12 == io_in_0_rs2_addr ? spec_table_18 : _GEN_49; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_51 = 5'h13 == io_in_0_rs2_addr ? spec_table_19 : _GEN_50; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_52 = 5'h14 == io_in_0_rs2_addr ? spec_table_20 : _GEN_51; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_53 = 5'h15 == io_in_0_rs2_addr ? spec_table_21 : _GEN_52; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_54 = 5'h16 == io_in_0_rs2_addr ? spec_table_22 : _GEN_53; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_55 = 5'h17 == io_in_0_rs2_addr ? spec_table_23 : _GEN_54; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_56 = 5'h18 == io_in_0_rs2_addr ? spec_table_24 : _GEN_55; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_57 = 5'h19 == io_in_0_rs2_addr ? spec_table_25 : _GEN_56; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_58 = 5'h1a == io_in_0_rs2_addr ? spec_table_26 : _GEN_57; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_59 = 5'h1b == io_in_0_rs2_addr ? spec_table_27 : _GEN_58; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_60 = 5'h1c == io_in_0_rs2_addr ? spec_table_28 : _GEN_59; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_61 = 5'h1d == io_in_0_rs2_addr ? spec_table_29 : _GEN_60; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_62 = 5'h1e == io_in_0_rs2_addr ? spec_table_30 : _GEN_61; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_65 = 5'h1 == io_rd_addr_0 ? spec_table_1 : spec_table_0; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_66 = 5'h2 == io_rd_addr_0 ? spec_table_2 : _GEN_65; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_67 = 5'h3 == io_rd_addr_0 ? spec_table_3 : _GEN_66; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_68 = 5'h4 == io_rd_addr_0 ? spec_table_4 : _GEN_67; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_69 = 5'h5 == io_rd_addr_0 ? spec_table_5 : _GEN_68; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_70 = 5'h6 == io_rd_addr_0 ? spec_table_6 : _GEN_69; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_71 = 5'h7 == io_rd_addr_0 ? spec_table_7 : _GEN_70; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_72 = 5'h8 == io_rd_addr_0 ? spec_table_8 : _GEN_71; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_73 = 5'h9 == io_rd_addr_0 ? spec_table_9 : _GEN_72; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_74 = 5'ha == io_rd_addr_0 ? spec_table_10 : _GEN_73; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_75 = 5'hb == io_rd_addr_0 ? spec_table_11 : _GEN_74; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_76 = 5'hc == io_rd_addr_0 ? spec_table_12 : _GEN_75; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_77 = 5'hd == io_rd_addr_0 ? spec_table_13 : _GEN_76; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_78 = 5'he == io_rd_addr_0 ? spec_table_14 : _GEN_77; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_79 = 5'hf == io_rd_addr_0 ? spec_table_15 : _GEN_78; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_80 = 5'h10 == io_rd_addr_0 ? spec_table_16 : _GEN_79; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_81 = 5'h11 == io_rd_addr_0 ? spec_table_17 : _GEN_80; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_82 = 5'h12 == io_rd_addr_0 ? spec_table_18 : _GEN_81; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_83 = 5'h13 == io_rd_addr_0 ? spec_table_19 : _GEN_82; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_84 = 5'h14 == io_rd_addr_0 ? spec_table_20 : _GEN_83; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_85 = 5'h15 == io_rd_addr_0 ? spec_table_21 : _GEN_84; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_86 = 5'h16 == io_rd_addr_0 ? spec_table_22 : _GEN_85; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_87 = 5'h17 == io_rd_addr_0 ? spec_table_23 : _GEN_86; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_88 = 5'h18 == io_rd_addr_0 ? spec_table_24 : _GEN_87; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_89 = 5'h19 == io_rd_addr_0 ? spec_table_25 : _GEN_88; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_90 = 5'h1a == io_rd_addr_0 ? spec_table_26 : _GEN_89; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_91 = 5'h1b == io_rd_addr_0 ? spec_table_27 : _GEN_90; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_92 = 5'h1c == io_rd_addr_0 ? spec_table_28 : _GEN_91; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_93 = 5'h1d == io_rd_addr_0 ? spec_table_29 : _GEN_92; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_94 = 5'h1e == io_rd_addr_0 ? spec_table_30 : _GEN_93; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_97 = 5'h1 == io_in_1_rs1_addr ? spec_table_1 : spec_table_0; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_98 = 5'h2 == io_in_1_rs1_addr ? spec_table_2 : _GEN_97; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_99 = 5'h3 == io_in_1_rs1_addr ? spec_table_3 : _GEN_98; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_100 = 5'h4 == io_in_1_rs1_addr ? spec_table_4 : _GEN_99; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_101 = 5'h5 == io_in_1_rs1_addr ? spec_table_5 : _GEN_100; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_102 = 5'h6 == io_in_1_rs1_addr ? spec_table_6 : _GEN_101; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_103 = 5'h7 == io_in_1_rs1_addr ? spec_table_7 : _GEN_102; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_104 = 5'h8 == io_in_1_rs1_addr ? spec_table_8 : _GEN_103; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_105 = 5'h9 == io_in_1_rs1_addr ? spec_table_9 : _GEN_104; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_106 = 5'ha == io_in_1_rs1_addr ? spec_table_10 : _GEN_105; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_107 = 5'hb == io_in_1_rs1_addr ? spec_table_11 : _GEN_106; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_108 = 5'hc == io_in_1_rs1_addr ? spec_table_12 : _GEN_107; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_109 = 5'hd == io_in_1_rs1_addr ? spec_table_13 : _GEN_108; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_110 = 5'he == io_in_1_rs1_addr ? spec_table_14 : _GEN_109; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_111 = 5'hf == io_in_1_rs1_addr ? spec_table_15 : _GEN_110; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_112 = 5'h10 == io_in_1_rs1_addr ? spec_table_16 : _GEN_111; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_113 = 5'h11 == io_in_1_rs1_addr ? spec_table_17 : _GEN_112; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_114 = 5'h12 == io_in_1_rs1_addr ? spec_table_18 : _GEN_113; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_115 = 5'h13 == io_in_1_rs1_addr ? spec_table_19 : _GEN_114; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_116 = 5'h14 == io_in_1_rs1_addr ? spec_table_20 : _GEN_115; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_117 = 5'h15 == io_in_1_rs1_addr ? spec_table_21 : _GEN_116; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_118 = 5'h16 == io_in_1_rs1_addr ? spec_table_22 : _GEN_117; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_119 = 5'h17 == io_in_1_rs1_addr ? spec_table_23 : _GEN_118; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_120 = 5'h18 == io_in_1_rs1_addr ? spec_table_24 : _GEN_119; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_121 = 5'h19 == io_in_1_rs1_addr ? spec_table_25 : _GEN_120; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_122 = 5'h1a == io_in_1_rs1_addr ? spec_table_26 : _GEN_121; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_123 = 5'h1b == io_in_1_rs1_addr ? spec_table_27 : _GEN_122; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_124 = 5'h1c == io_in_1_rs1_addr ? spec_table_28 : _GEN_123; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_125 = 5'h1d == io_in_1_rs1_addr ? spec_table_29 : _GEN_124; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_126 = 5'h1e == io_in_1_rs1_addr ? spec_table_30 : _GEN_125; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_127 = 5'h1f == io_in_1_rs1_addr ? spec_table_31 : _GEN_126; // @[Rename.scala 121:{21,21}]
  wire [5:0] _GEN_129 = 5'h1 == io_in_1_rs2_addr ? spec_table_1 : spec_table_0; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_130 = 5'h2 == io_in_1_rs2_addr ? spec_table_2 : _GEN_129; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_131 = 5'h3 == io_in_1_rs2_addr ? spec_table_3 : _GEN_130; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_132 = 5'h4 == io_in_1_rs2_addr ? spec_table_4 : _GEN_131; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_133 = 5'h5 == io_in_1_rs2_addr ? spec_table_5 : _GEN_132; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_134 = 5'h6 == io_in_1_rs2_addr ? spec_table_6 : _GEN_133; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_135 = 5'h7 == io_in_1_rs2_addr ? spec_table_7 : _GEN_134; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_136 = 5'h8 == io_in_1_rs2_addr ? spec_table_8 : _GEN_135; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_137 = 5'h9 == io_in_1_rs2_addr ? spec_table_9 : _GEN_136; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_138 = 5'ha == io_in_1_rs2_addr ? spec_table_10 : _GEN_137; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_139 = 5'hb == io_in_1_rs2_addr ? spec_table_11 : _GEN_138; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_140 = 5'hc == io_in_1_rs2_addr ? spec_table_12 : _GEN_139; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_141 = 5'hd == io_in_1_rs2_addr ? spec_table_13 : _GEN_140; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_142 = 5'he == io_in_1_rs2_addr ? spec_table_14 : _GEN_141; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_143 = 5'hf == io_in_1_rs2_addr ? spec_table_15 : _GEN_142; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_144 = 5'h10 == io_in_1_rs2_addr ? spec_table_16 : _GEN_143; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_145 = 5'h11 == io_in_1_rs2_addr ? spec_table_17 : _GEN_144; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_146 = 5'h12 == io_in_1_rs2_addr ? spec_table_18 : _GEN_145; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_147 = 5'h13 == io_in_1_rs2_addr ? spec_table_19 : _GEN_146; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_148 = 5'h14 == io_in_1_rs2_addr ? spec_table_20 : _GEN_147; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_149 = 5'h15 == io_in_1_rs2_addr ? spec_table_21 : _GEN_148; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_150 = 5'h16 == io_in_1_rs2_addr ? spec_table_22 : _GEN_149; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_151 = 5'h17 == io_in_1_rs2_addr ? spec_table_23 : _GEN_150; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_152 = 5'h18 == io_in_1_rs2_addr ? spec_table_24 : _GEN_151; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_153 = 5'h19 == io_in_1_rs2_addr ? spec_table_25 : _GEN_152; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_154 = 5'h1a == io_in_1_rs2_addr ? spec_table_26 : _GEN_153; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_155 = 5'h1b == io_in_1_rs2_addr ? spec_table_27 : _GEN_154; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_156 = 5'h1c == io_in_1_rs2_addr ? spec_table_28 : _GEN_155; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_157 = 5'h1d == io_in_1_rs2_addr ? spec_table_29 : _GEN_156; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_158 = 5'h1e == io_in_1_rs2_addr ? spec_table_30 : _GEN_157; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_159 = 5'h1f == io_in_1_rs2_addr ? spec_table_31 : _GEN_158; // @[Rename.scala 122:{21,21}]
  wire [5:0] _GEN_161 = 5'h1 == io_rd_addr_1 ? spec_table_1 : spec_table_0; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_162 = 5'h2 == io_rd_addr_1 ? spec_table_2 : _GEN_161; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_163 = 5'h3 == io_rd_addr_1 ? spec_table_3 : _GEN_162; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_164 = 5'h4 == io_rd_addr_1 ? spec_table_4 : _GEN_163; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_165 = 5'h5 == io_rd_addr_1 ? spec_table_5 : _GEN_164; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_166 = 5'h6 == io_rd_addr_1 ? spec_table_6 : _GEN_165; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_167 = 5'h7 == io_rd_addr_1 ? spec_table_7 : _GEN_166; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_168 = 5'h8 == io_rd_addr_1 ? spec_table_8 : _GEN_167; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_169 = 5'h9 == io_rd_addr_1 ? spec_table_9 : _GEN_168; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_170 = 5'ha == io_rd_addr_1 ? spec_table_10 : _GEN_169; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_171 = 5'hb == io_rd_addr_1 ? spec_table_11 : _GEN_170; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_172 = 5'hc == io_rd_addr_1 ? spec_table_12 : _GEN_171; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_173 = 5'hd == io_rd_addr_1 ? spec_table_13 : _GEN_172; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_174 = 5'he == io_rd_addr_1 ? spec_table_14 : _GEN_173; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_175 = 5'hf == io_rd_addr_1 ? spec_table_15 : _GEN_174; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_176 = 5'h10 == io_rd_addr_1 ? spec_table_16 : _GEN_175; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_177 = 5'h11 == io_rd_addr_1 ? spec_table_17 : _GEN_176; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_178 = 5'h12 == io_rd_addr_1 ? spec_table_18 : _GEN_177; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_179 = 5'h13 == io_rd_addr_1 ? spec_table_19 : _GEN_178; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_180 = 5'h14 == io_rd_addr_1 ? spec_table_20 : _GEN_179; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_181 = 5'h15 == io_rd_addr_1 ? spec_table_21 : _GEN_180; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_182 = 5'h16 == io_rd_addr_1 ? spec_table_22 : _GEN_181; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_183 = 5'h17 == io_rd_addr_1 ? spec_table_23 : _GEN_182; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_184 = 5'h18 == io_rd_addr_1 ? spec_table_24 : _GEN_183; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_185 = 5'h19 == io_rd_addr_1 ? spec_table_25 : _GEN_184; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_186 = 5'h1a == io_rd_addr_1 ? spec_table_26 : _GEN_185; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_187 = 5'h1b == io_rd_addr_1 ? spec_table_27 : _GEN_186; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_188 = 5'h1c == io_rd_addr_1 ? spec_table_28 : _GEN_187; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_189 = 5'h1d == io_rd_addr_1 ? spec_table_29 : _GEN_188; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_190 = 5'h1e == io_rd_addr_1 ? spec_table_30 : _GEN_189; // @[Rename.scala 123:{21,21}]
  wire [5:0] _GEN_191 = 5'h1f == io_rd_addr_1 ? spec_table_31 : _GEN_190; // @[Rename.scala 123:{21,21}]
  wire  _T_1 = io_rd_addr_0 != 5'h0; // @[Rename.scala 128:65]
  wire [5:0] _GEN_195 = 5'h0 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_0; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_196 = 5'h1 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_1; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_197 = 5'h2 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_2; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_198 = 5'h3 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_3; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_199 = 5'h4 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_4; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_200 = 5'h5 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_5; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_201 = 5'h6 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_6; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_202 = 5'h7 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_7; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_203 = 5'h8 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_8; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_204 = 5'h9 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_9; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_205 = 5'ha == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_10; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_206 = 5'hb == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_11; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_207 = 5'hc == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_12; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_208 = 5'hd == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_13; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_209 = 5'he == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_14; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_210 = 5'hf == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_15; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_211 = 5'h10 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_16; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_212 = 5'h11 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_17; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_213 = 5'h12 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_18; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_214 = 5'h13 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_19; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_215 = 5'h14 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_20; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_216 = 5'h15 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_21; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_217 = 5'h16 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_22; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_218 = 5'h17 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_23; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_219 = 5'h18 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_24; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_220 = 5'h19 == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_25; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_221 = 5'h1a == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_26; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_222 = 5'h1b == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_27; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_223 = 5'h1c == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_28; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_224 = 5'h1d == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_29; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_225 = 5'h1e == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_30; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_226 = 5'h1f == io_rd_addr_0 ? io_rd_paddr_0 : spec_table_31; // @[Rename.scala 117:27 145:{35,35}]
  wire [5:0] _GEN_227 = _T_1 & io_en ? _GEN_195 : spec_table_0; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_228 = _T_1 & io_en ? _GEN_196 : spec_table_1; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_229 = _T_1 & io_en ? _GEN_197 : spec_table_2; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_230 = _T_1 & io_en ? _GEN_198 : spec_table_3; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_231 = _T_1 & io_en ? _GEN_199 : spec_table_4; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_232 = _T_1 & io_en ? _GEN_200 : spec_table_5; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_233 = _T_1 & io_en ? _GEN_201 : spec_table_6; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_234 = _T_1 & io_en ? _GEN_202 : spec_table_7; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_235 = _T_1 & io_en ? _GEN_203 : spec_table_8; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_236 = _T_1 & io_en ? _GEN_204 : spec_table_9; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_237 = _T_1 & io_en ? _GEN_205 : spec_table_10; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_238 = _T_1 & io_en ? _GEN_206 : spec_table_11; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_239 = _T_1 & io_en ? _GEN_207 : spec_table_12; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_240 = _T_1 & io_en ? _GEN_208 : spec_table_13; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_241 = _T_1 & io_en ? _GEN_209 : spec_table_14; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_242 = _T_1 & io_en ? _GEN_210 : spec_table_15; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_243 = _T_1 & io_en ? _GEN_211 : spec_table_16; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_244 = _T_1 & io_en ? _GEN_212 : spec_table_17; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_245 = _T_1 & io_en ? _GEN_213 : spec_table_18; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_246 = _T_1 & io_en ? _GEN_214 : spec_table_19; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_247 = _T_1 & io_en ? _GEN_215 : spec_table_20; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_248 = _T_1 & io_en ? _GEN_216 : spec_table_21; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_249 = _T_1 & io_en ? _GEN_217 : spec_table_22; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_250 = _T_1 & io_en ? _GEN_218 : spec_table_23; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_251 = _T_1 & io_en ? _GEN_219 : spec_table_24; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_252 = _T_1 & io_en ? _GEN_220 : spec_table_25; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_253 = _T_1 & io_en ? _GEN_221 : spec_table_26; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_254 = _T_1 & io_en ? _GEN_222 : spec_table_27; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_255 = _T_1 & io_en ? _GEN_223 : spec_table_28; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_256 = _T_1 & io_en ? _GEN_224 : spec_table_29; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_257 = _T_1 & io_en ? _GEN_225 : spec_table_30; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_258 = _T_1 & io_en ? _GEN_226 : spec_table_31; // @[Rename.scala 117:27 144:45]
  wire [5:0] _GEN_323 = 5'h0 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_0; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_324 = 5'h1 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_1; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_325 = 5'h2 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_2; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_326 = 5'h3 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_3; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_327 = 5'h4 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_4; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_328 = 5'h5 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_5; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_329 = 5'h6 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_6; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_330 = 5'h7 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_7; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_331 = 5'h8 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_8; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_332 = 5'h9 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_9; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_333 = 5'ha == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_10; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_334 = 5'hb == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_11; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_335 = 5'hc == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_12; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_336 = 5'hd == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_13; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_337 = 5'he == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_14; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_338 = 5'hf == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_15; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_339 = 5'h10 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_16; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_340 = 5'h11 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_17; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_341 = 5'h12 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_18; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_342 = 5'h13 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_19; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_343 = 5'h14 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_20; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_344 = 5'h15 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_21; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_345 = 5'h16 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_22; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_346 = 5'h17 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_23; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_347 = 5'h18 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_24; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_348 = 5'h19 == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_25; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_349 = 5'h1a == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_26; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_350 = 5'h1b == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_27; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_351 = 5'h1c == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_28; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_352 = 5'h1d == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_29; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_353 = 5'h1e == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_30; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_354 = 5'h1f == io_cm_rd_addr_0 ? io_cm_rd_paddr_0 : arch_table_31; // @[Rename.scala 118:27 150:{38,38}]
  wire [5:0] _GEN_355 = io_cm_rd_addr_0 != 5'h0 ? _GEN_323 : arch_table_0; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_356 = io_cm_rd_addr_0 != 5'h0 ? _GEN_324 : arch_table_1; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_357 = io_cm_rd_addr_0 != 5'h0 ? _GEN_325 : arch_table_2; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_358 = io_cm_rd_addr_0 != 5'h0 ? _GEN_326 : arch_table_3; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_359 = io_cm_rd_addr_0 != 5'h0 ? _GEN_327 : arch_table_4; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_360 = io_cm_rd_addr_0 != 5'h0 ? _GEN_328 : arch_table_5; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_361 = io_cm_rd_addr_0 != 5'h0 ? _GEN_329 : arch_table_6; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_362 = io_cm_rd_addr_0 != 5'h0 ? _GEN_330 : arch_table_7; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_363 = io_cm_rd_addr_0 != 5'h0 ? _GEN_331 : arch_table_8; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_364 = io_cm_rd_addr_0 != 5'h0 ? _GEN_332 : arch_table_9; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_365 = io_cm_rd_addr_0 != 5'h0 ? _GEN_333 : arch_table_10; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_366 = io_cm_rd_addr_0 != 5'h0 ? _GEN_334 : arch_table_11; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_367 = io_cm_rd_addr_0 != 5'h0 ? _GEN_335 : arch_table_12; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_368 = io_cm_rd_addr_0 != 5'h0 ? _GEN_336 : arch_table_13; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_369 = io_cm_rd_addr_0 != 5'h0 ? _GEN_337 : arch_table_14; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_370 = io_cm_rd_addr_0 != 5'h0 ? _GEN_338 : arch_table_15; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_371 = io_cm_rd_addr_0 != 5'h0 ? _GEN_339 : arch_table_16; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_372 = io_cm_rd_addr_0 != 5'h0 ? _GEN_340 : arch_table_17; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_373 = io_cm_rd_addr_0 != 5'h0 ? _GEN_341 : arch_table_18; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_374 = io_cm_rd_addr_0 != 5'h0 ? _GEN_342 : arch_table_19; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_375 = io_cm_rd_addr_0 != 5'h0 ? _GEN_343 : arch_table_20; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_376 = io_cm_rd_addr_0 != 5'h0 ? _GEN_344 : arch_table_21; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_377 = io_cm_rd_addr_0 != 5'h0 ? _GEN_345 : arch_table_22; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_378 = io_cm_rd_addr_0 != 5'h0 ? _GEN_346 : arch_table_23; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_379 = io_cm_rd_addr_0 != 5'h0 ? _GEN_347 : arch_table_24; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_380 = io_cm_rd_addr_0 != 5'h0 ? _GEN_348 : arch_table_25; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_381 = io_cm_rd_addr_0 != 5'h0 ? _GEN_349 : arch_table_26; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_382 = io_cm_rd_addr_0 != 5'h0 ? _GEN_350 : arch_table_27; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_383 = io_cm_rd_addr_0 != 5'h0 ? _GEN_351 : arch_table_28; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_384 = io_cm_rd_addr_0 != 5'h0 ? _GEN_352 : arch_table_29; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_385 = io_cm_rd_addr_0 != 5'h0 ? _GEN_353 : arch_table_30; // @[Rename.scala 118:27 149:39]
  wire [5:0] _GEN_386 = io_cm_rd_addr_0 != 5'h0 ? _GEN_354 : arch_table_31; // @[Rename.scala 118:27 149:39]
  assign io_rs1_paddr_0 = 5'h1f == io_in_0_rs1_addr ? spec_table_31 : _GEN_30; // @[Rename.scala 121:{21,21}]
  assign io_rs1_paddr_1 = io_in_1_rs1_addr == io_rd_addr_0 & io_rd_addr_0 != 5'h0 ? io_rd_paddr_0 : _GEN_127; // @[Rename.scala 121:21 128:75 129:21]
  assign io_rs2_paddr_0 = 5'h1f == io_in_0_rs2_addr ? spec_table_31 : _GEN_62; // @[Rename.scala 122:{21,21}]
  assign io_rs2_paddr_1 = io_in_1_rs2_addr == io_rd_addr_0 & _T_1 ? io_rd_paddr_0 : _GEN_159; // @[Rename.scala 122:21 131:75 132:21]
  assign io_rd_ppaddr_0 = 5'h1f == io_rd_addr_0 ? spec_table_31 : _GEN_94; // @[Rename.scala 123:{21,21}]
  assign io_rd_ppaddr_1 = io_in_1_rd_addr == io_rd_addr_0 & _T_1 ? io_rd_paddr_0 : _GEN_191; // @[Rename.scala 123:21 135:74 136:21]
  always @(posedge clock) begin
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_0 <= 6'h0; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_0 <= arch_table_0; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h0 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_0 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_0 <= _GEN_227;
      end
    end else begin
      spec_table_0 <= _GEN_227;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_1 <= 6'h1; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_1 <= arch_table_1; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h1 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_1 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_1 <= _GEN_228;
      end
    end else begin
      spec_table_1 <= _GEN_228;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_2 <= 6'h2; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_2 <= arch_table_2; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h2 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_2 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_2 <= _GEN_229;
      end
    end else begin
      spec_table_2 <= _GEN_229;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_3 <= 6'h3; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_3 <= arch_table_3; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h3 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_3 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_3 <= _GEN_230;
      end
    end else begin
      spec_table_3 <= _GEN_230;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_4 <= 6'h4; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_4 <= arch_table_4; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h4 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_4 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_4 <= _GEN_231;
      end
    end else begin
      spec_table_4 <= _GEN_231;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_5 <= 6'h5; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_5 <= arch_table_5; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h5 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_5 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_5 <= _GEN_232;
      end
    end else begin
      spec_table_5 <= _GEN_232;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_6 <= 6'h6; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_6 <= arch_table_6; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h6 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_6 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_6 <= _GEN_233;
      end
    end else begin
      spec_table_6 <= _GEN_233;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_7 <= 6'h7; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_7 <= arch_table_7; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h7 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_7 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_7 <= _GEN_234;
      end
    end else begin
      spec_table_7 <= _GEN_234;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_8 <= 6'h8; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_8 <= arch_table_8; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h8 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_8 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_8 <= _GEN_235;
      end
    end else begin
      spec_table_8 <= _GEN_235;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_9 <= 6'h9; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_9 <= arch_table_9; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h9 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_9 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_9 <= _GEN_236;
      end
    end else begin
      spec_table_9 <= _GEN_236;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_10 <= 6'ha; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_10 <= arch_table_10; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'ha == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_10 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_10 <= _GEN_237;
      end
    end else begin
      spec_table_10 <= _GEN_237;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_11 <= 6'hb; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_11 <= arch_table_11; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'hb == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_11 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_11 <= _GEN_238;
      end
    end else begin
      spec_table_11 <= _GEN_238;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_12 <= 6'hc; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_12 <= arch_table_12; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'hc == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_12 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_12 <= _GEN_239;
      end
    end else begin
      spec_table_12 <= _GEN_239;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_13 <= 6'hd; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_13 <= arch_table_13; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'hd == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_13 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_13 <= _GEN_240;
      end
    end else begin
      spec_table_13 <= _GEN_240;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_14 <= 6'he; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_14 <= arch_table_14; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'he == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_14 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_14 <= _GEN_241;
      end
    end else begin
      spec_table_14 <= _GEN_241;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_15 <= 6'hf; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_15 <= arch_table_15; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'hf == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_15 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_15 <= _GEN_242;
      end
    end else begin
      spec_table_15 <= _GEN_242;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_16 <= 6'h10; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_16 <= arch_table_16; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h10 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_16 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_16 <= _GEN_243;
      end
    end else begin
      spec_table_16 <= _GEN_243;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_17 <= 6'h11; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_17 <= arch_table_17; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h11 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_17 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_17 <= _GEN_244;
      end
    end else begin
      spec_table_17 <= _GEN_244;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_18 <= 6'h12; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_18 <= arch_table_18; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h12 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_18 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_18 <= _GEN_245;
      end
    end else begin
      spec_table_18 <= _GEN_245;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_19 <= 6'h13; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_19 <= arch_table_19; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h13 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_19 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_19 <= _GEN_246;
      end
    end else begin
      spec_table_19 <= _GEN_246;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_20 <= 6'h14; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_20 <= arch_table_20; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h14 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_20 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_20 <= _GEN_247;
      end
    end else begin
      spec_table_20 <= _GEN_247;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_21 <= 6'h15; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_21 <= arch_table_21; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h15 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_21 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_21 <= _GEN_248;
      end
    end else begin
      spec_table_21 <= _GEN_248;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_22 <= 6'h16; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_22 <= arch_table_22; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h16 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_22 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_22 <= _GEN_249;
      end
    end else begin
      spec_table_22 <= _GEN_249;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_23 <= 6'h17; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_23 <= arch_table_23; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h17 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_23 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_23 <= _GEN_250;
      end
    end else begin
      spec_table_23 <= _GEN_250;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_24 <= 6'h18; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_24 <= arch_table_24; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h18 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_24 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_24 <= _GEN_251;
      end
    end else begin
      spec_table_24 <= _GEN_251;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_25 <= 6'h19; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_25 <= arch_table_25; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h19 == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_25 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_25 <= _GEN_252;
      end
    end else begin
      spec_table_25 <= _GEN_252;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_26 <= 6'h1a; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_26 <= arch_table_26; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h1a == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_26 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_26 <= _GEN_253;
      end
    end else begin
      spec_table_26 <= _GEN_253;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_27 <= 6'h1b; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_27 <= arch_table_27; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h1b == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_27 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_27 <= _GEN_254;
      end
    end else begin
      spec_table_27 <= _GEN_254;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_28 <= 6'h1c; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_28 <= arch_table_28; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h1c == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_28 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_28 <= _GEN_255;
      end
    end else begin
      spec_table_28 <= _GEN_255;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_29 <= 6'h1d; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_29 <= arch_table_29; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h1d == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_29 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_29 <= _GEN_256;
      end
    end else begin
      spec_table_29 <= _GEN_256;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_30 <= 6'h1e; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_30 <= arch_table_30; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h1e == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_30 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_30 <= _GEN_257;
      end
    end else begin
      spec_table_30 <= _GEN_257;
    end
    if (reset) begin // @[Rename.scala 117:27]
      spec_table_31 <= 6'h1f; // @[Rename.scala 117:27]
    end else if (io_cm_recover) begin // @[Rename.scala 139:24]
      spec_table_31 <= arch_table_31; // @[Rename.scala 140:16]
    end else if (io_rd_addr_1 != 5'h0 & io_en) begin // @[Rename.scala 144:45]
      if (5'h1f == io_rd_addr_1) begin // @[Rename.scala 145:35]
        spec_table_31 <= io_rd_paddr_1; // @[Rename.scala 145:35]
      end else begin
        spec_table_31 <= _GEN_258;
      end
    end else begin
      spec_table_31 <= _GEN_258;
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_0 <= 6'h0; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h0 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_0 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_0 <= _GEN_355;
        end
      end else begin
        arch_table_0 <= _GEN_355;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_1 <= 6'h1; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h1 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_1 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_1 <= _GEN_356;
        end
      end else begin
        arch_table_1 <= _GEN_356;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_2 <= 6'h2; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h2 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_2 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_2 <= _GEN_357;
        end
      end else begin
        arch_table_2 <= _GEN_357;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_3 <= 6'h3; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h3 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_3 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_3 <= _GEN_358;
        end
      end else begin
        arch_table_3 <= _GEN_358;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_4 <= 6'h4; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h4 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_4 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_4 <= _GEN_359;
        end
      end else begin
        arch_table_4 <= _GEN_359;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_5 <= 6'h5; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h5 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_5 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_5 <= _GEN_360;
        end
      end else begin
        arch_table_5 <= _GEN_360;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_6 <= 6'h6; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h6 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_6 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_6 <= _GEN_361;
        end
      end else begin
        arch_table_6 <= _GEN_361;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_7 <= 6'h7; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h7 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_7 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_7 <= _GEN_362;
        end
      end else begin
        arch_table_7 <= _GEN_362;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_8 <= 6'h8; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h8 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_8 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_8 <= _GEN_363;
        end
      end else begin
        arch_table_8 <= _GEN_363;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_9 <= 6'h9; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h9 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_9 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_9 <= _GEN_364;
        end
      end else begin
        arch_table_9 <= _GEN_364;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_10 <= 6'ha; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'ha == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_10 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_10 <= _GEN_365;
        end
      end else begin
        arch_table_10 <= _GEN_365;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_11 <= 6'hb; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'hb == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_11 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_11 <= _GEN_366;
        end
      end else begin
        arch_table_11 <= _GEN_366;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_12 <= 6'hc; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'hc == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_12 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_12 <= _GEN_367;
        end
      end else begin
        arch_table_12 <= _GEN_367;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_13 <= 6'hd; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'hd == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_13 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_13 <= _GEN_368;
        end
      end else begin
        arch_table_13 <= _GEN_368;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_14 <= 6'he; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'he == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_14 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_14 <= _GEN_369;
        end
      end else begin
        arch_table_14 <= _GEN_369;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_15 <= 6'hf; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'hf == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_15 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_15 <= _GEN_370;
        end
      end else begin
        arch_table_15 <= _GEN_370;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_16 <= 6'h10; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h10 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_16 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_16 <= _GEN_371;
        end
      end else begin
        arch_table_16 <= _GEN_371;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_17 <= 6'h11; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h11 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_17 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_17 <= _GEN_372;
        end
      end else begin
        arch_table_17 <= _GEN_372;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_18 <= 6'h12; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h12 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_18 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_18 <= _GEN_373;
        end
      end else begin
        arch_table_18 <= _GEN_373;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_19 <= 6'h13; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h13 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_19 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_19 <= _GEN_374;
        end
      end else begin
        arch_table_19 <= _GEN_374;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_20 <= 6'h14; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h14 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_20 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_20 <= _GEN_375;
        end
      end else begin
        arch_table_20 <= _GEN_375;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_21 <= 6'h15; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h15 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_21 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_21 <= _GEN_376;
        end
      end else begin
        arch_table_21 <= _GEN_376;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_22 <= 6'h16; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h16 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_22 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_22 <= _GEN_377;
        end
      end else begin
        arch_table_22 <= _GEN_377;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_23 <= 6'h17; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h17 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_23 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_23 <= _GEN_378;
        end
      end else begin
        arch_table_23 <= _GEN_378;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_24 <= 6'h18; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h18 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_24 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_24 <= _GEN_379;
        end
      end else begin
        arch_table_24 <= _GEN_379;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_25 <= 6'h19; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h19 == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_25 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_25 <= _GEN_380;
        end
      end else begin
        arch_table_25 <= _GEN_380;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_26 <= 6'h1a; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h1a == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_26 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_26 <= _GEN_381;
        end
      end else begin
        arch_table_26 <= _GEN_381;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_27 <= 6'h1b; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h1b == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_27 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_27 <= _GEN_382;
        end
      end else begin
        arch_table_27 <= _GEN_382;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_28 <= 6'h1c; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h1c == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_28 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_28 <= _GEN_383;
        end
      end else begin
        arch_table_28 <= _GEN_383;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_29 <= 6'h1d; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h1d == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_29 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_29 <= _GEN_384;
        end
      end else begin
        arch_table_29 <= _GEN_384;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_30 <= 6'h1e; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h1e == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_30 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_30 <= _GEN_385;
        end
      end else begin
        arch_table_30 <= _GEN_385;
      end
    end
    if (reset) begin // @[Rename.scala 118:27]
      arch_table_31 <= 6'h1f; // @[Rename.scala 118:27]
    end else if (!(io_cm_recover)) begin // @[Rename.scala 139:24]
      if (io_cm_rd_addr_1 != 5'h0) begin // @[Rename.scala 149:39]
        if (5'h1f == io_cm_rd_addr_1) begin // @[Rename.scala 150:38]
          arch_table_31 <= io_cm_rd_paddr_1; // @[Rename.scala 150:38]
        end else begin
          arch_table_31 <= _GEN_386;
        end
      end else begin
        arch_table_31 <= _GEN_386;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  spec_table_0 = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  spec_table_1 = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  spec_table_2 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  spec_table_3 = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  spec_table_4 = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  spec_table_5 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  spec_table_6 = _RAND_6[5:0];
  _RAND_7 = {1{`RANDOM}};
  spec_table_7 = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  spec_table_8 = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  spec_table_9 = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  spec_table_10 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  spec_table_11 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  spec_table_12 = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  spec_table_13 = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  spec_table_14 = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  spec_table_15 = _RAND_15[5:0];
  _RAND_16 = {1{`RANDOM}};
  spec_table_16 = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  spec_table_17 = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  spec_table_18 = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  spec_table_19 = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  spec_table_20 = _RAND_20[5:0];
  _RAND_21 = {1{`RANDOM}};
  spec_table_21 = _RAND_21[5:0];
  _RAND_22 = {1{`RANDOM}};
  spec_table_22 = _RAND_22[5:0];
  _RAND_23 = {1{`RANDOM}};
  spec_table_23 = _RAND_23[5:0];
  _RAND_24 = {1{`RANDOM}};
  spec_table_24 = _RAND_24[5:0];
  _RAND_25 = {1{`RANDOM}};
  spec_table_25 = _RAND_25[5:0];
  _RAND_26 = {1{`RANDOM}};
  spec_table_26 = _RAND_26[5:0];
  _RAND_27 = {1{`RANDOM}};
  spec_table_27 = _RAND_27[5:0];
  _RAND_28 = {1{`RANDOM}};
  spec_table_28 = _RAND_28[5:0];
  _RAND_29 = {1{`RANDOM}};
  spec_table_29 = _RAND_29[5:0];
  _RAND_30 = {1{`RANDOM}};
  spec_table_30 = _RAND_30[5:0];
  _RAND_31 = {1{`RANDOM}};
  spec_table_31 = _RAND_31[5:0];
  _RAND_32 = {1{`RANDOM}};
  arch_table_0 = _RAND_32[5:0];
  _RAND_33 = {1{`RANDOM}};
  arch_table_1 = _RAND_33[5:0];
  _RAND_34 = {1{`RANDOM}};
  arch_table_2 = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  arch_table_3 = _RAND_35[5:0];
  _RAND_36 = {1{`RANDOM}};
  arch_table_4 = _RAND_36[5:0];
  _RAND_37 = {1{`RANDOM}};
  arch_table_5 = _RAND_37[5:0];
  _RAND_38 = {1{`RANDOM}};
  arch_table_6 = _RAND_38[5:0];
  _RAND_39 = {1{`RANDOM}};
  arch_table_7 = _RAND_39[5:0];
  _RAND_40 = {1{`RANDOM}};
  arch_table_8 = _RAND_40[5:0];
  _RAND_41 = {1{`RANDOM}};
  arch_table_9 = _RAND_41[5:0];
  _RAND_42 = {1{`RANDOM}};
  arch_table_10 = _RAND_42[5:0];
  _RAND_43 = {1{`RANDOM}};
  arch_table_11 = _RAND_43[5:0];
  _RAND_44 = {1{`RANDOM}};
  arch_table_12 = _RAND_44[5:0];
  _RAND_45 = {1{`RANDOM}};
  arch_table_13 = _RAND_45[5:0];
  _RAND_46 = {1{`RANDOM}};
  arch_table_14 = _RAND_46[5:0];
  _RAND_47 = {1{`RANDOM}};
  arch_table_15 = _RAND_47[5:0];
  _RAND_48 = {1{`RANDOM}};
  arch_table_16 = _RAND_48[5:0];
  _RAND_49 = {1{`RANDOM}};
  arch_table_17 = _RAND_49[5:0];
  _RAND_50 = {1{`RANDOM}};
  arch_table_18 = _RAND_50[5:0];
  _RAND_51 = {1{`RANDOM}};
  arch_table_19 = _RAND_51[5:0];
  _RAND_52 = {1{`RANDOM}};
  arch_table_20 = _RAND_52[5:0];
  _RAND_53 = {1{`RANDOM}};
  arch_table_21 = _RAND_53[5:0];
  _RAND_54 = {1{`RANDOM}};
  arch_table_22 = _RAND_54[5:0];
  _RAND_55 = {1{`RANDOM}};
  arch_table_23 = _RAND_55[5:0];
  _RAND_56 = {1{`RANDOM}};
  arch_table_24 = _RAND_56[5:0];
  _RAND_57 = {1{`RANDOM}};
  arch_table_25 = _RAND_57[5:0];
  _RAND_58 = {1{`RANDOM}};
  arch_table_26 = _RAND_58[5:0];
  _RAND_59 = {1{`RANDOM}};
  arch_table_27 = _RAND_59[5:0];
  _RAND_60 = {1{`RANDOM}};
  arch_table_28 = _RAND_60[5:0];
  _RAND_61 = {1{`RANDOM}};
  arch_table_29 = _RAND_61[5:0];
  _RAND_62 = {1{`RANDOM}};
  arch_table_30 = _RAND_62[5:0];
  _RAND_63 = {1{`RANDOM}};
  arch_table_31 = _RAND_63[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_Rename(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_vec_0_valid,
  input  [31:0] io_in_bits_vec_0_pc,
  input  [31:0] io_in_bits_vec_0_npc,
  input  [31:0] io_in_bits_vec_0_inst,
  input  [2:0]  io_in_bits_vec_0_fu_code,
  input  [3:0]  io_in_bits_vec_0_alu_code,
  input  [3:0]  io_in_bits_vec_0_jmp_code,
  input  [1:0]  io_in_bits_vec_0_mem_code,
  input  [1:0]  io_in_bits_vec_0_mem_size,
  input  [2:0]  io_in_bits_vec_0_sys_code,
  input         io_in_bits_vec_0_w_type,
  input  [1:0]  io_in_bits_vec_0_rs1_src,
  input  [1:0]  io_in_bits_vec_0_rs2_src,
  input  [4:0]  io_in_bits_vec_0_rs1_addr,
  input  [4:0]  io_in_bits_vec_0_rs2_addr,
  input  [4:0]  io_in_bits_vec_0_rd_addr,
  input         io_in_bits_vec_0_rd_en,
  input  [31:0] io_in_bits_vec_0_imm,
  input         io_in_bits_vec_0_pred_br,
  input  [31:0] io_in_bits_vec_0_pred_bpc,
  input         io_in_bits_vec_1_valid,
  input  [31:0] io_in_bits_vec_1_pc,
  input  [31:0] io_in_bits_vec_1_npc,
  input  [31:0] io_in_bits_vec_1_inst,
  input  [2:0]  io_in_bits_vec_1_fu_code,
  input  [3:0]  io_in_bits_vec_1_alu_code,
  input  [3:0]  io_in_bits_vec_1_jmp_code,
  input  [1:0]  io_in_bits_vec_1_mem_code,
  input  [1:0]  io_in_bits_vec_1_mem_size,
  input  [2:0]  io_in_bits_vec_1_sys_code,
  input         io_in_bits_vec_1_w_type,
  input  [1:0]  io_in_bits_vec_1_rs1_src,
  input  [1:0]  io_in_bits_vec_1_rs2_src,
  input  [4:0]  io_in_bits_vec_1_rs1_addr,
  input  [4:0]  io_in_bits_vec_1_rs2_addr,
  input  [4:0]  io_in_bits_vec_1_rd_addr,
  input         io_in_bits_vec_1_rd_en,
  input  [31:0] io_in_bits_vec_1_imm,
  input         io_in_bits_vec_1_pred_br,
  input  [31:0] io_in_bits_vec_1_pred_bpc,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_vec_0_valid,
  output [31:0] io_out_bits_vec_0_pc,
  output [31:0] io_out_bits_vec_0_npc,
  output [31:0] io_out_bits_vec_0_inst,
  output [2:0]  io_out_bits_vec_0_fu_code,
  output [3:0]  io_out_bits_vec_0_alu_code,
  output [3:0]  io_out_bits_vec_0_jmp_code,
  output [1:0]  io_out_bits_vec_0_mem_code,
  output [1:0]  io_out_bits_vec_0_mem_size,
  output [2:0]  io_out_bits_vec_0_sys_code,
  output        io_out_bits_vec_0_w_type,
  output [1:0]  io_out_bits_vec_0_rs1_src,
  output [1:0]  io_out_bits_vec_0_rs2_src,
  output [4:0]  io_out_bits_vec_0_rd_addr,
  output        io_out_bits_vec_0_rd_en,
  output [31:0] io_out_bits_vec_0_imm,
  output        io_out_bits_vec_0_pred_br,
  output [31:0] io_out_bits_vec_0_pred_bpc,
  output [5:0]  io_out_bits_vec_0_rs1_paddr,
  output [5:0]  io_out_bits_vec_0_rs2_paddr,
  output [5:0]  io_out_bits_vec_0_rd_paddr,
  output [5:0]  io_out_bits_vec_0_rd_ppaddr,
  output        io_out_bits_vec_1_valid,
  output [31:0] io_out_bits_vec_1_pc,
  output [31:0] io_out_bits_vec_1_npc,
  output [31:0] io_out_bits_vec_1_inst,
  output [2:0]  io_out_bits_vec_1_fu_code,
  output [3:0]  io_out_bits_vec_1_alu_code,
  output [3:0]  io_out_bits_vec_1_jmp_code,
  output [1:0]  io_out_bits_vec_1_mem_code,
  output [1:0]  io_out_bits_vec_1_mem_size,
  output [2:0]  io_out_bits_vec_1_sys_code,
  output        io_out_bits_vec_1_w_type,
  output [1:0]  io_out_bits_vec_1_rs1_src,
  output [1:0]  io_out_bits_vec_1_rs2_src,
  output [4:0]  io_out_bits_vec_1_rd_addr,
  output        io_out_bits_vec_1_rd_en,
  output [31:0] io_out_bits_vec_1_imm,
  output        io_out_bits_vec_1_pred_br,
  output [31:0] io_out_bits_vec_1_pred_bpc,
  output [5:0]  io_out_bits_vec_1_rs1_paddr,
  output [5:0]  io_out_bits_vec_1_rs2_paddr,
  output [5:0]  io_out_bits_vec_1_rd_paddr,
  output [5:0]  io_out_bits_vec_1_rd_ppaddr,
  output [63:0] io_avail_list,
  input         io_flush,
  input         io_exe_0_valid,
  input         io_exe_0_rd_en,
  input  [5:0]  io_exe_0_rd_paddr,
  input         io_exe_1_valid,
  input         io_exe_1_rd_en,
  input  [5:0]  io_exe_1_rd_paddr,
  input         io_exe_2_valid,
  input         io_exe_2_rd_en,
  input  [5:0]  io_exe_2_rd_paddr,
  input         io_cm_recover,
  input         io_cm_0_valid,
  input  [4:0]  io_cm_0_rd_addr,
  input         io_cm_0_rd_en,
  input  [5:0]  io_cm_0_rd_paddr,
  input  [5:0]  io_cm_0_rd_ppaddr,
  input         io_cm_1_valid,
  input  [4:0]  io_cm_1_rd_addr,
  input         io_cm_1_rd_en,
  input  [5:0]  io_cm_1_rd_paddr,
  input  [5:0]  io_cm_1_rd_ppaddr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
`endif // RANDOMIZE_REG_INIT
  wire  pst_clock; // @[Rename.scala 34:19]
  wire  pst_reset; // @[Rename.scala 34:19]
  wire  pst_io_en; // @[Rename.scala 34:19]
  wire  pst_io_allocatable; // @[Rename.scala 34:19]
  wire  pst_io_rd_req_0; // @[Rename.scala 34:19]
  wire  pst_io_rd_req_1; // @[Rename.scala 34:19]
  wire [5:0] pst_io_rd_paddr_0; // @[Rename.scala 34:19]
  wire [5:0] pst_io_rd_paddr_1; // @[Rename.scala 34:19]
  wire [5:0] pst_io_exe_0; // @[Rename.scala 34:19]
  wire [5:0] pst_io_exe_1; // @[Rename.scala 34:19]
  wire [5:0] pst_io_exe_2; // @[Rename.scala 34:19]
  wire [5:0] pst_io_cm_0; // @[Rename.scala 34:19]
  wire [5:0] pst_io_cm_1; // @[Rename.scala 34:19]
  wire [5:0] pst_io_free_0; // @[Rename.scala 34:19]
  wire [5:0] pst_io_free_1; // @[Rename.scala 34:19]
  wire  pst_io_cm_recover; // @[Rename.scala 34:19]
  wire [63:0] pst_io_avail_list; // @[Rename.scala 34:19]
  wire  rt_clock; // @[Rename.scala 49:18]
  wire  rt_reset; // @[Rename.scala 49:18]
  wire  rt_io_en; // @[Rename.scala 49:18]
  wire [4:0] rt_io_in_0_rs1_addr; // @[Rename.scala 49:18]
  wire [4:0] rt_io_in_0_rs2_addr; // @[Rename.scala 49:18]
  wire [4:0] rt_io_in_1_rs1_addr; // @[Rename.scala 49:18]
  wire [4:0] rt_io_in_1_rs2_addr; // @[Rename.scala 49:18]
  wire [4:0] rt_io_in_1_rd_addr; // @[Rename.scala 49:18]
  wire [5:0] rt_io_rs1_paddr_0; // @[Rename.scala 49:18]
  wire [5:0] rt_io_rs1_paddr_1; // @[Rename.scala 49:18]
  wire [5:0] rt_io_rs2_paddr_0; // @[Rename.scala 49:18]
  wire [5:0] rt_io_rs2_paddr_1; // @[Rename.scala 49:18]
  wire [4:0] rt_io_rd_addr_0; // @[Rename.scala 49:18]
  wire [4:0] rt_io_rd_addr_1; // @[Rename.scala 49:18]
  wire [5:0] rt_io_rd_ppaddr_0; // @[Rename.scala 49:18]
  wire [5:0] rt_io_rd_ppaddr_1; // @[Rename.scala 49:18]
  wire [5:0] rt_io_rd_paddr_0; // @[Rename.scala 49:18]
  wire [5:0] rt_io_rd_paddr_1; // @[Rename.scala 49:18]
  wire  rt_io_cm_recover; // @[Rename.scala 49:18]
  wire [4:0] rt_io_cm_rd_addr_0; // @[Rename.scala 49:18]
  wire [4:0] rt_io_cm_rd_addr_1; // @[Rename.scala 49:18]
  wire [5:0] rt_io_cm_rd_paddr_0; // @[Rename.scala 49:18]
  wire [5:0] rt_io_cm_rd_paddr_1; // @[Rename.scala 49:18]
  wire  _T = io_in_bits_vec_0_valid & io_in_bits_vec_0_rd_en; // @[Rename.scala 37:41]
  wire  _T_1 = io_in_bits_vec_1_valid & io_in_bits_vec_1_rd_en; // @[Rename.scala 37:41]
  wire  _T_8 = io_cm_0_valid & io_cm_0_rd_en; // @[Rename.scala 43:40]
  wire  _T_12 = io_cm_1_valid & io_cm_1_rd_en; // @[Rename.scala 43:40]
  reg  out_uop_0_valid; // @[Rename.scala 70:24]
  reg [31:0] out_uop_0_pc; // @[Rename.scala 70:24]
  reg [31:0] out_uop_0_npc; // @[Rename.scala 70:24]
  reg [31:0] out_uop_0_inst; // @[Rename.scala 70:24]
  reg [2:0] out_uop_0_fu_code; // @[Rename.scala 70:24]
  reg [3:0] out_uop_0_alu_code; // @[Rename.scala 70:24]
  reg [3:0] out_uop_0_jmp_code; // @[Rename.scala 70:24]
  reg [1:0] out_uop_0_mem_code; // @[Rename.scala 70:24]
  reg [1:0] out_uop_0_mem_size; // @[Rename.scala 70:24]
  reg [2:0] out_uop_0_sys_code; // @[Rename.scala 70:24]
  reg  out_uop_0_w_type; // @[Rename.scala 70:24]
  reg [1:0] out_uop_0_rs1_src; // @[Rename.scala 70:24]
  reg [1:0] out_uop_0_rs2_src; // @[Rename.scala 70:24]
  reg [4:0] out_uop_0_rd_addr; // @[Rename.scala 70:24]
  reg  out_uop_0_rd_en; // @[Rename.scala 70:24]
  reg [31:0] out_uop_0_imm; // @[Rename.scala 70:24]
  reg  out_uop_0_pred_br; // @[Rename.scala 70:24]
  reg [31:0] out_uop_0_pred_bpc; // @[Rename.scala 70:24]
  reg [5:0] out_uop_0_rs1_paddr; // @[Rename.scala 70:24]
  reg [5:0] out_uop_0_rs2_paddr; // @[Rename.scala 70:24]
  reg [5:0] out_uop_0_rd_paddr; // @[Rename.scala 70:24]
  reg [5:0] out_uop_0_rd_ppaddr; // @[Rename.scala 70:24]
  reg  out_uop_1_valid; // @[Rename.scala 70:24]
  reg [31:0] out_uop_1_pc; // @[Rename.scala 70:24]
  reg [31:0] out_uop_1_npc; // @[Rename.scala 70:24]
  reg [31:0] out_uop_1_inst; // @[Rename.scala 70:24]
  reg [2:0] out_uop_1_fu_code; // @[Rename.scala 70:24]
  reg [3:0] out_uop_1_alu_code; // @[Rename.scala 70:24]
  reg [3:0] out_uop_1_jmp_code; // @[Rename.scala 70:24]
  reg [1:0] out_uop_1_mem_code; // @[Rename.scala 70:24]
  reg [1:0] out_uop_1_mem_size; // @[Rename.scala 70:24]
  reg [2:0] out_uop_1_sys_code; // @[Rename.scala 70:24]
  reg  out_uop_1_w_type; // @[Rename.scala 70:24]
  reg [1:0] out_uop_1_rs1_src; // @[Rename.scala 70:24]
  reg [1:0] out_uop_1_rs2_src; // @[Rename.scala 70:24]
  reg [4:0] out_uop_1_rd_addr; // @[Rename.scala 70:24]
  reg  out_uop_1_rd_en; // @[Rename.scala 70:24]
  reg [31:0] out_uop_1_imm; // @[Rename.scala 70:24]
  reg  out_uop_1_pred_br; // @[Rename.scala 70:24]
  reg [31:0] out_uop_1_pred_bpc; // @[Rename.scala 70:24]
  reg [5:0] out_uop_1_rs1_paddr; // @[Rename.scala 70:24]
  reg [5:0] out_uop_1_rs2_paddr; // @[Rename.scala 70:24]
  reg [5:0] out_uop_1_rd_paddr; // @[Rename.scala 70:24]
  reg [5:0] out_uop_1_rd_ppaddr; // @[Rename.scala 70:24]
  reg  out_valid; // @[Rename.scala 71:26]
  wire [5:0] uop_0_rs1_paddr = rt_io_rs1_paddr_0;
  wire [5:0] uop_0_rs2_paddr = rt_io_rs2_paddr_0;
  wire [5:0] uop_0_rd_paddr = pst_io_rd_paddr_0;
  wire [5:0] uop_0_rd_ppaddr = rt_io_rd_ppaddr_0;
  wire [5:0] uop_1_rs1_paddr = rt_io_rs1_paddr_1;
  wire [5:0] uop_1_rs2_paddr = rt_io_rs2_paddr_1;
  wire [5:0] uop_1_rd_paddr = pst_io_rd_paddr_1;
  wire [5:0] uop_1_rd_ppaddr = rt_io_rd_ppaddr_1;
  ysyx_210128_PrfStateTable pst ( // @[Rename.scala 34:19]
    .clock(pst_clock),
    .reset(pst_reset),
    .io_en(pst_io_en),
    .io_allocatable(pst_io_allocatable),
    .io_rd_req_0(pst_io_rd_req_0),
    .io_rd_req_1(pst_io_rd_req_1),
    .io_rd_paddr_0(pst_io_rd_paddr_0),
    .io_rd_paddr_1(pst_io_rd_paddr_1),
    .io_exe_0(pst_io_exe_0),
    .io_exe_1(pst_io_exe_1),
    .io_exe_2(pst_io_exe_2),
    .io_cm_0(pst_io_cm_0),
    .io_cm_1(pst_io_cm_1),
    .io_free_0(pst_io_free_0),
    .io_free_1(pst_io_free_1),
    .io_cm_recover(pst_io_cm_recover),
    .io_avail_list(pst_io_avail_list)
  );
  ysyx_210128_RenameTable rt ( // @[Rename.scala 49:18]
    .clock(rt_clock),
    .reset(rt_reset),
    .io_en(rt_io_en),
    .io_in_0_rs1_addr(rt_io_in_0_rs1_addr),
    .io_in_0_rs2_addr(rt_io_in_0_rs2_addr),
    .io_in_1_rs1_addr(rt_io_in_1_rs1_addr),
    .io_in_1_rs2_addr(rt_io_in_1_rs2_addr),
    .io_in_1_rd_addr(rt_io_in_1_rd_addr),
    .io_rs1_paddr_0(rt_io_rs1_paddr_0),
    .io_rs1_paddr_1(rt_io_rs1_paddr_1),
    .io_rs2_paddr_0(rt_io_rs2_paddr_0),
    .io_rs2_paddr_1(rt_io_rs2_paddr_1),
    .io_rd_addr_0(rt_io_rd_addr_0),
    .io_rd_addr_1(rt_io_rd_addr_1),
    .io_rd_ppaddr_0(rt_io_rd_ppaddr_0),
    .io_rd_ppaddr_1(rt_io_rd_ppaddr_1),
    .io_rd_paddr_0(rt_io_rd_paddr_0),
    .io_rd_paddr_1(rt_io_rd_paddr_1),
    .io_cm_recover(rt_io_cm_recover),
    .io_cm_rd_addr_0(rt_io_cm_rd_addr_0),
    .io_cm_rd_addr_1(rt_io_cm_rd_addr_1),
    .io_cm_rd_paddr_0(rt_io_cm_rd_paddr_0),
    .io_cm_rd_paddr_1(rt_io_cm_rd_paddr_1)
  );
  assign io_in_ready = pst_io_allocatable & io_out_ready; // @[Rename.scala 66:37]
  assign io_out_valid = out_valid; // @[Rename.scala 86:16]
  assign io_out_bits_vec_0_valid = out_uop_0_valid; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_pc = out_uop_0_pc; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_npc = out_uop_0_npc; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_inst = out_uop_0_inst; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_fu_code = out_uop_0_fu_code; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_alu_code = out_uop_0_alu_code; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_jmp_code = out_uop_0_jmp_code; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_mem_code = out_uop_0_mem_code; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_mem_size = out_uop_0_mem_size; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_sys_code = out_uop_0_sys_code; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_w_type = out_uop_0_w_type; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_rs1_src = out_uop_0_rs1_src; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_rs2_src = out_uop_0_rs2_src; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_rd_addr = out_uop_0_rd_addr; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_rd_en = out_uop_0_rd_en; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_imm = out_uop_0_imm; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_pred_br = out_uop_0_pred_br; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_pred_bpc = out_uop_0_pred_bpc; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_rs1_paddr = out_uop_0_rs1_paddr; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_rs2_paddr = out_uop_0_rs2_paddr; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_rd_paddr = out_uop_0_rd_paddr; // @[Rename.scala 85:19]
  assign io_out_bits_vec_0_rd_ppaddr = out_uop_0_rd_ppaddr; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_valid = out_uop_1_valid; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_pc = out_uop_1_pc; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_npc = out_uop_1_npc; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_inst = out_uop_1_inst; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_fu_code = out_uop_1_fu_code; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_alu_code = out_uop_1_alu_code; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_jmp_code = out_uop_1_jmp_code; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_mem_code = out_uop_1_mem_code; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_mem_size = out_uop_1_mem_size; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_sys_code = out_uop_1_sys_code; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_w_type = out_uop_1_w_type; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_rs1_src = out_uop_1_rs1_src; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_rs2_src = out_uop_1_rs2_src; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_rd_addr = out_uop_1_rd_addr; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_rd_en = out_uop_1_rd_en; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_imm = out_uop_1_imm; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_pred_br = out_uop_1_pred_br; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_pred_bpc = out_uop_1_pred_bpc; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_rs1_paddr = out_uop_1_rs1_paddr; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_rs2_paddr = out_uop_1_rs2_paddr; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_rd_paddr = out_uop_1_rd_paddr; // @[Rename.scala 85:19]
  assign io_out_bits_vec_1_rd_ppaddr = out_uop_1_rd_ppaddr; // @[Rename.scala 85:19]
  assign io_avail_list = pst_io_avail_list; // @[Rename.scala 47:17]
  assign pst_clock = clock;
  assign pst_reset = reset;
  assign pst_io_en = io_out_ready & io_in_valid; // @[Rename.scala 28:25]
  assign pst_io_rd_req_0 = io_in_bits_vec_0_valid & io_in_bits_vec_0_rd_en; // @[Rename.scala 37:41]
  assign pst_io_rd_req_1 = io_in_bits_vec_1_valid & io_in_bits_vec_1_rd_en; // @[Rename.scala 37:41]
  assign pst_io_exe_0 = io_exe_0_valid & io_exe_0_rd_en ? io_exe_0_rd_paddr : 6'h0; // @[Rename.scala 40:25]
  assign pst_io_exe_1 = io_exe_1_valid & io_exe_1_rd_en ? io_exe_1_rd_paddr : 6'h0; // @[Rename.scala 40:25]
  assign pst_io_exe_2 = io_exe_2_valid & io_exe_2_rd_en ? io_exe_2_rd_paddr : 6'h0; // @[Rename.scala 40:25]
  assign pst_io_cm_0 = io_cm_0_valid & io_cm_0_rd_en ? io_cm_0_rd_paddr : 6'h0; // @[Rename.scala 43:24]
  assign pst_io_cm_1 = io_cm_1_valid & io_cm_1_rd_en ? io_cm_1_rd_paddr : 6'h0; // @[Rename.scala 43:24]
  assign pst_io_free_0 = _T_8 ? io_cm_0_rd_ppaddr : 6'h0; // @[Rename.scala 44:26]
  assign pst_io_free_1 = _T_12 ? io_cm_1_rd_ppaddr : 6'h0; // @[Rename.scala 44:26]
  assign pst_io_cm_recover = io_cm_recover; // @[Rename.scala 46:21]
  assign rt_clock = clock;
  assign rt_reset = reset;
  assign rt_io_en = io_out_ready & io_in_valid; // @[Rename.scala 28:25]
  assign rt_io_in_0_rs1_addr = io_in_bits_vec_0_rs1_addr; // @[Rename.scala 51:12]
  assign rt_io_in_0_rs2_addr = io_in_bits_vec_0_rs2_addr; // @[Rename.scala 51:12]
  assign rt_io_in_1_rs1_addr = io_in_bits_vec_1_rs1_addr; // @[Rename.scala 51:12]
  assign rt_io_in_1_rs2_addr = io_in_bits_vec_1_rs2_addr; // @[Rename.scala 51:12]
  assign rt_io_in_1_rd_addr = io_in_bits_vec_1_rd_addr; // @[Rename.scala 51:12]
  assign rt_io_rd_addr_0 = _T ? io_in_bits_vec_0_rd_addr : 5'h0; // @[Rename.scala 55:29]
  assign rt_io_rd_addr_1 = _T_1 ? io_in_bits_vec_1_rd_addr : 5'h0; // @[Rename.scala 55:29]
  assign rt_io_rd_paddr_0 = pst_io_rd_paddr_0; // @[Rename.scala 57:23]
  assign rt_io_rd_paddr_1 = pst_io_rd_paddr_1; // @[Rename.scala 57:23]
  assign rt_io_cm_recover = io_cm_recover; // @[Rename.scala 60:21]
  assign rt_io_cm_rd_addr_0 = _T_8 ? io_cm_0_rd_addr : 5'h0; // @[Rename.scala 62:32]
  assign rt_io_cm_rd_addr_1 = _T_12 ? io_cm_1_rd_addr : 5'h0; // @[Rename.scala 62:32]
  assign rt_io_cm_rd_paddr_0 = io_cm_0_rd_paddr; // @[Rename.scala 63:26]
  assign rt_io_cm_rd_paddr_1 = io_cm_1_rd_paddr; // @[Rename.scala 63:26]
  always @(posedge clock) begin
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_valid <= 1'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_valid <= 1'h0; // @[Rename.scala 75:18]
    end else begin
      out_uop_0_valid <= io_in_bits_vec_0_valid; // @[Rename.scala 80:18]
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_pc <= 32'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_pc <= 32'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_pc <= io_in_bits_vec_0_pc;
    end else begin
      out_uop_0_pc <= 32'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_npc <= 32'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_npc <= 32'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_npc <= io_in_bits_vec_0_npc;
    end else begin
      out_uop_0_npc <= 32'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_inst <= 32'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_inst <= 32'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_inst <= io_in_bits_vec_0_inst;
    end else begin
      out_uop_0_inst <= 32'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_fu_code <= 3'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_fu_code <= 3'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_fu_code <= io_in_bits_vec_0_fu_code;
    end else begin
      out_uop_0_fu_code <= 3'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_alu_code <= 4'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_alu_code <= 4'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_alu_code <= io_in_bits_vec_0_alu_code;
    end else begin
      out_uop_0_alu_code <= 4'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_jmp_code <= 4'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_jmp_code <= 4'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_jmp_code <= io_in_bits_vec_0_jmp_code;
    end else begin
      out_uop_0_jmp_code <= 4'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_mem_code <= 2'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_mem_code <= 2'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_mem_code <= io_in_bits_vec_0_mem_code;
    end else begin
      out_uop_0_mem_code <= 2'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_mem_size <= 2'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_mem_size <= 2'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_mem_size <= io_in_bits_vec_0_mem_size;
    end else begin
      out_uop_0_mem_size <= 2'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_sys_code <= 3'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_sys_code <= 3'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_sys_code <= io_in_bits_vec_0_sys_code;
    end else begin
      out_uop_0_sys_code <= 3'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_w_type <= 1'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_w_type <= 1'h0; // @[Rename.scala 75:18]
    end else begin
      out_uop_0_w_type <= io_in_bits_vec_0_valid & io_in_bits_vec_0_w_type; // @[Rename.scala 80:18]
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_rs1_src <= 2'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_rs1_src <= 2'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_rs1_src <= io_in_bits_vec_0_rs1_src;
    end else begin
      out_uop_0_rs1_src <= 2'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_rs2_src <= 2'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_rs2_src <= 2'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_rs2_src <= io_in_bits_vec_0_rs2_src;
    end else begin
      out_uop_0_rs2_src <= 2'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_rd_addr <= 5'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_rd_addr <= 5'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_rd_addr <= io_in_bits_vec_0_rd_addr;
    end else begin
      out_uop_0_rd_addr <= 5'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_rd_en <= 1'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_rd_en <= 1'h0; // @[Rename.scala 75:18]
    end else begin
      out_uop_0_rd_en <= _T; // @[Rename.scala 80:18]
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_imm <= 32'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_imm <= 32'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_imm <= io_in_bits_vec_0_imm;
    end else begin
      out_uop_0_imm <= 32'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_pred_br <= 1'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_pred_br <= 1'h0; // @[Rename.scala 75:18]
    end else begin
      out_uop_0_pred_br <= io_in_bits_vec_0_valid & io_in_bits_vec_0_pred_br; // @[Rename.scala 80:18]
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_pred_bpc <= 32'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_pred_bpc <= 32'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_pred_bpc <= io_in_bits_vec_0_pred_bpc;
    end else begin
      out_uop_0_pred_bpc <= 32'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_rs1_paddr <= 6'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_rs1_paddr <= 6'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_rs1_paddr <= uop_0_rs1_paddr;
    end else begin
      out_uop_0_rs1_paddr <= 6'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_rs2_paddr <= 6'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_rs2_paddr <= 6'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_rs2_paddr <= uop_0_rs2_paddr;
    end else begin
      out_uop_0_rs2_paddr <= 6'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_rd_paddr <= 6'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_rd_paddr <= 6'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_rd_paddr <= uop_0_rd_paddr;
    end else begin
      out_uop_0_rd_paddr <= 6'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_0_rd_ppaddr <= 6'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_0_rd_ppaddr <= 6'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_0_valid) begin // @[Rename.scala 80:24]
      out_uop_0_rd_ppaddr <= uop_0_rd_ppaddr;
    end else begin
      out_uop_0_rd_ppaddr <= 6'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_valid <= 1'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_valid <= 1'h0; // @[Rename.scala 75:18]
    end else begin
      out_uop_1_valid <= io_in_bits_vec_1_valid; // @[Rename.scala 80:18]
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_pc <= 32'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_pc <= 32'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_pc <= io_in_bits_vec_1_pc;
    end else begin
      out_uop_1_pc <= 32'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_npc <= 32'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_npc <= 32'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_npc <= io_in_bits_vec_1_npc;
    end else begin
      out_uop_1_npc <= 32'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_inst <= 32'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_inst <= 32'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_inst <= io_in_bits_vec_1_inst;
    end else begin
      out_uop_1_inst <= 32'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_fu_code <= 3'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_fu_code <= 3'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_fu_code <= io_in_bits_vec_1_fu_code;
    end else begin
      out_uop_1_fu_code <= 3'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_alu_code <= 4'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_alu_code <= 4'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_alu_code <= io_in_bits_vec_1_alu_code;
    end else begin
      out_uop_1_alu_code <= 4'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_jmp_code <= 4'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_jmp_code <= 4'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_jmp_code <= io_in_bits_vec_1_jmp_code;
    end else begin
      out_uop_1_jmp_code <= 4'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_mem_code <= 2'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_mem_code <= 2'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_mem_code <= io_in_bits_vec_1_mem_code;
    end else begin
      out_uop_1_mem_code <= 2'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_mem_size <= 2'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_mem_size <= 2'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_mem_size <= io_in_bits_vec_1_mem_size;
    end else begin
      out_uop_1_mem_size <= 2'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_sys_code <= 3'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_sys_code <= 3'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_sys_code <= io_in_bits_vec_1_sys_code;
    end else begin
      out_uop_1_sys_code <= 3'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_w_type <= 1'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_w_type <= 1'h0; // @[Rename.scala 75:18]
    end else begin
      out_uop_1_w_type <= io_in_bits_vec_1_valid & io_in_bits_vec_1_w_type; // @[Rename.scala 80:18]
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_rs1_src <= 2'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_rs1_src <= 2'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_rs1_src <= io_in_bits_vec_1_rs1_src;
    end else begin
      out_uop_1_rs1_src <= 2'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_rs2_src <= 2'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_rs2_src <= 2'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_rs2_src <= io_in_bits_vec_1_rs2_src;
    end else begin
      out_uop_1_rs2_src <= 2'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_rd_addr <= 5'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_rd_addr <= 5'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_rd_addr <= io_in_bits_vec_1_rd_addr;
    end else begin
      out_uop_1_rd_addr <= 5'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_rd_en <= 1'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_rd_en <= 1'h0; // @[Rename.scala 75:18]
    end else begin
      out_uop_1_rd_en <= _T_1; // @[Rename.scala 80:18]
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_imm <= 32'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_imm <= 32'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_imm <= io_in_bits_vec_1_imm;
    end else begin
      out_uop_1_imm <= 32'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_pred_br <= 1'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_pred_br <= 1'h0; // @[Rename.scala 75:18]
    end else begin
      out_uop_1_pred_br <= io_in_bits_vec_1_valid & io_in_bits_vec_1_pred_br; // @[Rename.scala 80:18]
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_pred_bpc <= 32'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_pred_bpc <= 32'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_pred_bpc <= io_in_bits_vec_1_pred_bpc;
    end else begin
      out_uop_1_pred_bpc <= 32'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_rs1_paddr <= 6'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_rs1_paddr <= 6'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_rs1_paddr <= uop_1_rs1_paddr;
    end else begin
      out_uop_1_rs1_paddr <= 6'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_rs2_paddr <= 6'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_rs2_paddr <= 6'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_rs2_paddr <= uop_1_rs2_paddr;
    end else begin
      out_uop_1_rs2_paddr <= 6'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_rd_paddr <= 6'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_rd_paddr <= 6'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_rd_paddr <= uop_1_rd_paddr;
    end else begin
      out_uop_1_rd_paddr <= 6'h0;
    end
    if (reset) begin // @[Rename.scala 70:24]
      out_uop_1_rd_ppaddr <= 6'h0; // @[Rename.scala 70:24]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_uop_1_rd_ppaddr <= 6'h0; // @[Rename.scala 75:18]
    end else if (io_in_bits_vec_1_valid) begin // @[Rename.scala 80:24]
      out_uop_1_rd_ppaddr <= uop_1_rd_ppaddr;
    end else begin
      out_uop_1_rd_ppaddr <= 6'h0;
    end
    if (reset) begin // @[Rename.scala 71:26]
      out_valid <= 1'h0; // @[Rename.scala 71:26]
    end else if (io_flush) begin // @[Rename.scala 73:19]
      out_valid <= 1'h0; // @[Rename.scala 77:15]
    end else begin
      out_valid <= io_in_valid; // @[Rename.scala 82:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_uop_0_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_uop_0_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  out_uop_0_npc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  out_uop_0_inst = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  out_uop_0_fu_code = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  out_uop_0_alu_code = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  out_uop_0_jmp_code = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  out_uop_0_mem_code = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  out_uop_0_mem_size = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  out_uop_0_sys_code = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  out_uop_0_w_type = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  out_uop_0_rs1_src = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  out_uop_0_rs2_src = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  out_uop_0_rd_addr = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  out_uop_0_rd_en = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  out_uop_0_imm = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  out_uop_0_pred_br = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  out_uop_0_pred_bpc = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  out_uop_0_rs1_paddr = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  out_uop_0_rs2_paddr = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  out_uop_0_rd_paddr = _RAND_20[5:0];
  _RAND_21 = {1{`RANDOM}};
  out_uop_0_rd_ppaddr = _RAND_21[5:0];
  _RAND_22 = {1{`RANDOM}};
  out_uop_1_valid = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  out_uop_1_pc = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  out_uop_1_npc = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  out_uop_1_inst = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  out_uop_1_fu_code = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  out_uop_1_alu_code = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  out_uop_1_jmp_code = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  out_uop_1_mem_code = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  out_uop_1_mem_size = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  out_uop_1_sys_code = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  out_uop_1_w_type = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  out_uop_1_rs1_src = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  out_uop_1_rs2_src = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  out_uop_1_rd_addr = _RAND_35[4:0];
  _RAND_36 = {1{`RANDOM}};
  out_uop_1_rd_en = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  out_uop_1_imm = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  out_uop_1_pred_br = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  out_uop_1_pred_bpc = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  out_uop_1_rs1_paddr = _RAND_40[5:0];
  _RAND_41 = {1{`RANDOM}};
  out_uop_1_rs2_paddr = _RAND_41[5:0];
  _RAND_42 = {1{`RANDOM}};
  out_uop_1_rd_paddr = _RAND_42[5:0];
  _RAND_43 = {1{`RANDOM}};
  out_uop_1_rd_ppaddr = _RAND_43[5:0];
  _RAND_44 = {1{`RANDOM}};
  out_valid = _RAND_44[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_StallRegister(
  input         clock,
  input         reset,
  input         io_flush,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_vec_0_valid,
  input  [31:0] io_in_bits_vec_0_pc,
  input  [31:0] io_in_bits_vec_0_npc,
  input  [31:0] io_in_bits_vec_0_inst,
  input  [2:0]  io_in_bits_vec_0_fu_code,
  input  [3:0]  io_in_bits_vec_0_alu_code,
  input  [3:0]  io_in_bits_vec_0_jmp_code,
  input  [1:0]  io_in_bits_vec_0_mem_code,
  input  [1:0]  io_in_bits_vec_0_mem_size,
  input  [2:0]  io_in_bits_vec_0_sys_code,
  input         io_in_bits_vec_0_w_type,
  input  [1:0]  io_in_bits_vec_0_rs1_src,
  input  [1:0]  io_in_bits_vec_0_rs2_src,
  input  [4:0]  io_in_bits_vec_0_rd_addr,
  input         io_in_bits_vec_0_rd_en,
  input  [31:0] io_in_bits_vec_0_imm,
  input         io_in_bits_vec_0_pred_br,
  input  [31:0] io_in_bits_vec_0_pred_bpc,
  input  [5:0]  io_in_bits_vec_0_rs1_paddr,
  input  [5:0]  io_in_bits_vec_0_rs2_paddr,
  input  [5:0]  io_in_bits_vec_0_rd_paddr,
  input  [5:0]  io_in_bits_vec_0_rd_ppaddr,
  input         io_in_bits_vec_1_valid,
  input  [31:0] io_in_bits_vec_1_pc,
  input  [31:0] io_in_bits_vec_1_npc,
  input  [31:0] io_in_bits_vec_1_inst,
  input  [2:0]  io_in_bits_vec_1_fu_code,
  input  [3:0]  io_in_bits_vec_1_alu_code,
  input  [3:0]  io_in_bits_vec_1_jmp_code,
  input  [1:0]  io_in_bits_vec_1_mem_code,
  input  [1:0]  io_in_bits_vec_1_mem_size,
  input  [2:0]  io_in_bits_vec_1_sys_code,
  input         io_in_bits_vec_1_w_type,
  input  [1:0]  io_in_bits_vec_1_rs1_src,
  input  [1:0]  io_in_bits_vec_1_rs2_src,
  input  [4:0]  io_in_bits_vec_1_rd_addr,
  input         io_in_bits_vec_1_rd_en,
  input  [31:0] io_in_bits_vec_1_imm,
  input         io_in_bits_vec_1_pred_br,
  input  [31:0] io_in_bits_vec_1_pred_bpc,
  input  [5:0]  io_in_bits_vec_1_rs1_paddr,
  input  [5:0]  io_in_bits_vec_1_rs2_paddr,
  input  [5:0]  io_in_bits_vec_1_rd_paddr,
  input  [5:0]  io_in_bits_vec_1_rd_ppaddr,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_vec_0_valid,
  output [31:0] io_out_bits_vec_0_pc,
  output [31:0] io_out_bits_vec_0_npc,
  output [31:0] io_out_bits_vec_0_inst,
  output [2:0]  io_out_bits_vec_0_fu_code,
  output [3:0]  io_out_bits_vec_0_alu_code,
  output [3:0]  io_out_bits_vec_0_jmp_code,
  output [1:0]  io_out_bits_vec_0_mem_code,
  output [1:0]  io_out_bits_vec_0_mem_size,
  output [2:0]  io_out_bits_vec_0_sys_code,
  output        io_out_bits_vec_0_w_type,
  output [1:0]  io_out_bits_vec_0_rs1_src,
  output [1:0]  io_out_bits_vec_0_rs2_src,
  output [4:0]  io_out_bits_vec_0_rd_addr,
  output        io_out_bits_vec_0_rd_en,
  output [31:0] io_out_bits_vec_0_imm,
  output        io_out_bits_vec_0_pred_br,
  output [31:0] io_out_bits_vec_0_pred_bpc,
  output [5:0]  io_out_bits_vec_0_rs1_paddr,
  output [5:0]  io_out_bits_vec_0_rs2_paddr,
  output [5:0]  io_out_bits_vec_0_rd_paddr,
  output [5:0]  io_out_bits_vec_0_rd_ppaddr,
  output        io_out_bits_vec_1_valid,
  output [31:0] io_out_bits_vec_1_pc,
  output [31:0] io_out_bits_vec_1_npc,
  output [31:0] io_out_bits_vec_1_inst,
  output [2:0]  io_out_bits_vec_1_fu_code,
  output [3:0]  io_out_bits_vec_1_alu_code,
  output [3:0]  io_out_bits_vec_1_jmp_code,
  output [1:0]  io_out_bits_vec_1_mem_code,
  output [1:0]  io_out_bits_vec_1_mem_size,
  output [2:0]  io_out_bits_vec_1_sys_code,
  output        io_out_bits_vec_1_w_type,
  output [1:0]  io_out_bits_vec_1_rs1_src,
  output [1:0]  io_out_bits_vec_1_rs2_src,
  output [4:0]  io_out_bits_vec_1_rd_addr,
  output        io_out_bits_vec_1_rd_en,
  output [31:0] io_out_bits_vec_1_imm,
  output        io_out_bits_vec_1_pred_br,
  output [31:0] io_out_bits_vec_1_pred_bpc,
  output [5:0]  io_out_bits_vec_1_rs1_paddr,
  output [5:0]  io_out_bits_vec_1_rs2_paddr,
  output [5:0]  io_out_bits_vec_1_rd_paddr,
  output [5:0]  io_out_bits_vec_1_rd_ppaddr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
`endif // RANDOMIZE_REG_INIT
  reg  reg_in_0_valid; // @[StallRegister.scala 17:23]
  reg [31:0] reg_in_0_pc; // @[StallRegister.scala 17:23]
  reg [31:0] reg_in_0_npc; // @[StallRegister.scala 17:23]
  reg [31:0] reg_in_0_inst; // @[StallRegister.scala 17:23]
  reg [2:0] reg_in_0_fu_code; // @[StallRegister.scala 17:23]
  reg [3:0] reg_in_0_alu_code; // @[StallRegister.scala 17:23]
  reg [3:0] reg_in_0_jmp_code; // @[StallRegister.scala 17:23]
  reg [1:0] reg_in_0_mem_code; // @[StallRegister.scala 17:23]
  reg [1:0] reg_in_0_mem_size; // @[StallRegister.scala 17:23]
  reg [2:0] reg_in_0_sys_code; // @[StallRegister.scala 17:23]
  reg  reg_in_0_w_type; // @[StallRegister.scala 17:23]
  reg [1:0] reg_in_0_rs1_src; // @[StallRegister.scala 17:23]
  reg [1:0] reg_in_0_rs2_src; // @[StallRegister.scala 17:23]
  reg [4:0] reg_in_0_rd_addr; // @[StallRegister.scala 17:23]
  reg  reg_in_0_rd_en; // @[StallRegister.scala 17:23]
  reg [31:0] reg_in_0_imm; // @[StallRegister.scala 17:23]
  reg  reg_in_0_pred_br; // @[StallRegister.scala 17:23]
  reg [31:0] reg_in_0_pred_bpc; // @[StallRegister.scala 17:23]
  reg [5:0] reg_in_0_rs1_paddr; // @[StallRegister.scala 17:23]
  reg [5:0] reg_in_0_rs2_paddr; // @[StallRegister.scala 17:23]
  reg [5:0] reg_in_0_rd_paddr; // @[StallRegister.scala 17:23]
  reg [5:0] reg_in_0_rd_ppaddr; // @[StallRegister.scala 17:23]
  reg  reg_in_1_valid; // @[StallRegister.scala 17:23]
  reg [31:0] reg_in_1_pc; // @[StallRegister.scala 17:23]
  reg [31:0] reg_in_1_npc; // @[StallRegister.scala 17:23]
  reg [31:0] reg_in_1_inst; // @[StallRegister.scala 17:23]
  reg [2:0] reg_in_1_fu_code; // @[StallRegister.scala 17:23]
  reg [3:0] reg_in_1_alu_code; // @[StallRegister.scala 17:23]
  reg [3:0] reg_in_1_jmp_code; // @[StallRegister.scala 17:23]
  reg [1:0] reg_in_1_mem_code; // @[StallRegister.scala 17:23]
  reg [1:0] reg_in_1_mem_size; // @[StallRegister.scala 17:23]
  reg [2:0] reg_in_1_sys_code; // @[StallRegister.scala 17:23]
  reg  reg_in_1_w_type; // @[StallRegister.scala 17:23]
  reg [1:0] reg_in_1_rs1_src; // @[StallRegister.scala 17:23]
  reg [1:0] reg_in_1_rs2_src; // @[StallRegister.scala 17:23]
  reg [4:0] reg_in_1_rd_addr; // @[StallRegister.scala 17:23]
  reg  reg_in_1_rd_en; // @[StallRegister.scala 17:23]
  reg [31:0] reg_in_1_imm; // @[StallRegister.scala 17:23]
  reg  reg_in_1_pred_br; // @[StallRegister.scala 17:23]
  reg [31:0] reg_in_1_pred_bpc; // @[StallRegister.scala 17:23]
  reg [5:0] reg_in_1_rs1_paddr; // @[StallRegister.scala 17:23]
  reg [5:0] reg_in_1_rs2_paddr; // @[StallRegister.scala 17:23]
  reg [5:0] reg_in_1_rd_paddr; // @[StallRegister.scala 17:23]
  reg [5:0] reg_in_1_rd_ppaddr; // @[StallRegister.scala 17:23]
  reg  reg_in_valid; // @[StallRegister.scala 18:29]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg  REG; // @[StallRegister.scala 22:68]
  wire  _GEN_50 = io_in_valid & ~io_flush & ~io_out_ready & REG | reg_in_valid; // @[StallRegister.scala 22:84 24:18 18:29]
  reg  REG_1; // @[StallRegister.scala 27:32]
  assign io_in_ready = io_out_ready; // @[StallRegister.scala 35:15]
  assign io_out_valid = io_out_ready & REG_1 ? reg_in_valid : io_in_valid; // @[StallRegister.scala 27:49 29:18 33:18]
  assign io_out_bits_vec_0_valid = io_out_ready & REG_1 ? reg_in_0_valid : io_in_bits_vec_0_valid; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_pc = io_out_ready & REG_1 ? reg_in_0_pc : io_in_bits_vec_0_pc; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_npc = io_out_ready & REG_1 ? reg_in_0_npc : io_in_bits_vec_0_npc; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_inst = io_out_ready & REG_1 ? reg_in_0_inst : io_in_bits_vec_0_inst; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_fu_code = io_out_ready & REG_1 ? reg_in_0_fu_code : io_in_bits_vec_0_fu_code; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_alu_code = io_out_ready & REG_1 ? reg_in_0_alu_code : io_in_bits_vec_0_alu_code; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_jmp_code = io_out_ready & REG_1 ? reg_in_0_jmp_code : io_in_bits_vec_0_jmp_code; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_mem_code = io_out_ready & REG_1 ? reg_in_0_mem_code : io_in_bits_vec_0_mem_code; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_mem_size = io_out_ready & REG_1 ? reg_in_0_mem_size : io_in_bits_vec_0_mem_size; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_sys_code = io_out_ready & REG_1 ? reg_in_0_sys_code : io_in_bits_vec_0_sys_code; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_w_type = io_out_ready & REG_1 ? reg_in_0_w_type : io_in_bits_vec_0_w_type; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_rs1_src = io_out_ready & REG_1 ? reg_in_0_rs1_src : io_in_bits_vec_0_rs1_src; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_rs2_src = io_out_ready & REG_1 ? reg_in_0_rs2_src : io_in_bits_vec_0_rs2_src; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_rd_addr = io_out_ready & REG_1 ? reg_in_0_rd_addr : io_in_bits_vec_0_rd_addr; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_rd_en = io_out_ready & REG_1 ? reg_in_0_rd_en : io_in_bits_vec_0_rd_en; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_imm = io_out_ready & REG_1 ? reg_in_0_imm : io_in_bits_vec_0_imm; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_pred_br = io_out_ready & REG_1 ? reg_in_0_pred_br : io_in_bits_vec_0_pred_br; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_pred_bpc = io_out_ready & REG_1 ? reg_in_0_pred_bpc : io_in_bits_vec_0_pred_bpc; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_rs1_paddr = io_out_ready & REG_1 ? reg_in_0_rs1_paddr : io_in_bits_vec_0_rs1_paddr; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_rs2_paddr = io_out_ready & REG_1 ? reg_in_0_rs2_paddr : io_in_bits_vec_0_rs2_paddr; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_rd_paddr = io_out_ready & REG_1 ? reg_in_0_rd_paddr : io_in_bits_vec_0_rd_paddr; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_0_rd_ppaddr = io_out_ready & REG_1 ? reg_in_0_rd_ppaddr : io_in_bits_vec_0_rd_ppaddr; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_valid = io_out_ready & REG_1 ? reg_in_1_valid : io_in_bits_vec_1_valid; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_pc = io_out_ready & REG_1 ? reg_in_1_pc : io_in_bits_vec_1_pc; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_npc = io_out_ready & REG_1 ? reg_in_1_npc : io_in_bits_vec_1_npc; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_inst = io_out_ready & REG_1 ? reg_in_1_inst : io_in_bits_vec_1_inst; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_fu_code = io_out_ready & REG_1 ? reg_in_1_fu_code : io_in_bits_vec_1_fu_code; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_alu_code = io_out_ready & REG_1 ? reg_in_1_alu_code : io_in_bits_vec_1_alu_code; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_jmp_code = io_out_ready & REG_1 ? reg_in_1_jmp_code : io_in_bits_vec_1_jmp_code; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_mem_code = io_out_ready & REG_1 ? reg_in_1_mem_code : io_in_bits_vec_1_mem_code; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_mem_size = io_out_ready & REG_1 ? reg_in_1_mem_size : io_in_bits_vec_1_mem_size; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_sys_code = io_out_ready & REG_1 ? reg_in_1_sys_code : io_in_bits_vec_1_sys_code; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_w_type = io_out_ready & REG_1 ? reg_in_1_w_type : io_in_bits_vec_1_w_type; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_rs1_src = io_out_ready & REG_1 ? reg_in_1_rs1_src : io_in_bits_vec_1_rs1_src; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_rs2_src = io_out_ready & REG_1 ? reg_in_1_rs2_src : io_in_bits_vec_1_rs2_src; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_rd_addr = io_out_ready & REG_1 ? reg_in_1_rd_addr : io_in_bits_vec_1_rd_addr; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_rd_en = io_out_ready & REG_1 ? reg_in_1_rd_en : io_in_bits_vec_1_rd_en; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_imm = io_out_ready & REG_1 ? reg_in_1_imm : io_in_bits_vec_1_imm; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_pred_br = io_out_ready & REG_1 ? reg_in_1_pred_br : io_in_bits_vec_1_pred_br; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_pred_bpc = io_out_ready & REG_1 ? reg_in_1_pred_bpc : io_in_bits_vec_1_pred_bpc; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_rs1_paddr = io_out_ready & REG_1 ? reg_in_1_rs1_paddr : io_in_bits_vec_1_rs1_paddr; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_rs2_paddr = io_out_ready & REG_1 ? reg_in_1_rs2_paddr : io_in_bits_vec_1_rs2_paddr; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_rd_paddr = io_out_ready & REG_1 ? reg_in_1_rd_paddr : io_in_bits_vec_1_rd_paddr; // @[StallRegister.scala 27:49 28:21 32:21]
  assign io_out_bits_vec_1_rd_ppaddr = io_out_ready & REG_1 ? reg_in_1_rd_ppaddr : io_in_bits_vec_1_rd_ppaddr; // @[StallRegister.scala 27:49 28:21 32:21]
  always @(posedge clock) begin
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_valid <= 1'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_valid <= io_in_bits_vec_0_valid; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_pc <= 32'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_pc <= io_in_bits_vec_0_pc; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_npc <= 32'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_npc <= io_in_bits_vec_0_npc; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_inst <= 32'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_inst <= io_in_bits_vec_0_inst; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_fu_code <= 3'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_fu_code <= io_in_bits_vec_0_fu_code; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_alu_code <= 4'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_alu_code <= io_in_bits_vec_0_alu_code; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_jmp_code <= 4'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_jmp_code <= io_in_bits_vec_0_jmp_code; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_mem_code <= 2'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_mem_code <= io_in_bits_vec_0_mem_code; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_mem_size <= 2'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_mem_size <= io_in_bits_vec_0_mem_size; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_sys_code <= 3'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_sys_code <= io_in_bits_vec_0_sys_code; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_w_type <= 1'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_w_type <= io_in_bits_vec_0_w_type; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_rs1_src <= 2'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_rs1_src <= io_in_bits_vec_0_rs1_src; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_rs2_src <= 2'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_rs2_src <= io_in_bits_vec_0_rs2_src; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_rd_addr <= 5'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_rd_addr <= io_in_bits_vec_0_rd_addr; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_rd_en <= 1'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_rd_en <= io_in_bits_vec_0_rd_en; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_imm <= 32'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_imm <= io_in_bits_vec_0_imm; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_pred_br <= 1'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_pred_br <= io_in_bits_vec_0_pred_br; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_pred_bpc <= 32'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_pred_bpc <= io_in_bits_vec_0_pred_bpc; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_rs1_paddr <= 6'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_rs1_paddr <= io_in_bits_vec_0_rs1_paddr; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_rs2_paddr <= 6'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_rs2_paddr <= io_in_bits_vec_0_rs2_paddr; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_rd_paddr <= 6'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_rd_paddr <= io_in_bits_vec_0_rd_paddr; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_0_rd_ppaddr <= 6'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_0_rd_ppaddr <= io_in_bits_vec_0_rd_ppaddr; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_valid <= 1'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_valid <= io_in_bits_vec_1_valid; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_pc <= 32'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_pc <= io_in_bits_vec_1_pc; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_npc <= 32'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_npc <= io_in_bits_vec_1_npc; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_inst <= 32'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_inst <= io_in_bits_vec_1_inst; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_fu_code <= 3'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_fu_code <= io_in_bits_vec_1_fu_code; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_alu_code <= 4'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_alu_code <= io_in_bits_vec_1_alu_code; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_jmp_code <= 4'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_jmp_code <= io_in_bits_vec_1_jmp_code; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_mem_code <= 2'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_mem_code <= io_in_bits_vec_1_mem_code; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_mem_size <= 2'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_mem_size <= io_in_bits_vec_1_mem_size; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_sys_code <= 3'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_sys_code <= io_in_bits_vec_1_sys_code; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_w_type <= 1'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_w_type <= io_in_bits_vec_1_w_type; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_rs1_src <= 2'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_rs1_src <= io_in_bits_vec_1_rs1_src; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_rs2_src <= 2'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_rs2_src <= io_in_bits_vec_1_rs2_src; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_rd_addr <= 5'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_rd_addr <= io_in_bits_vec_1_rd_addr; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_rd_en <= 1'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_rd_en <= io_in_bits_vec_1_rd_en; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_imm <= 32'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_imm <= io_in_bits_vec_1_imm; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_pred_br <= 1'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_pred_br <= io_in_bits_vec_1_pred_br; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_pred_bpc <= 32'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_pred_bpc <= io_in_bits_vec_1_pred_bpc; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_rs1_paddr <= 6'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_rs2_paddr <= 6'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_rd_paddr <= 6'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 17:23]
      reg_in_1_rd_ppaddr <= 6'h0; // @[StallRegister.scala 17:23]
    end else if (!(io_flush | _T)) begin // @[StallRegister.scala 20:36]
      if (io_in_valid & ~io_flush & ~io_out_ready & REG) begin // @[StallRegister.scala 22:84]
        reg_in_1_rd_ppaddr <= io_in_bits_vec_1_rd_ppaddr; // @[StallRegister.scala 23:12]
      end
    end
    if (reset) begin // @[StallRegister.scala 18:29]
      reg_in_valid <= 1'h0; // @[StallRegister.scala 18:29]
    end else if (io_out_ready & REG_1) begin // @[StallRegister.scala 27:49]
      reg_in_valid <= 1'h0; // @[StallRegister.scala 30:18]
    end else if (io_flush | _T) begin // @[StallRegister.scala 20:36]
      reg_in_valid <= 1'h0; // @[StallRegister.scala 21:18]
    end else begin
      reg_in_valid <= _GEN_50;
    end
    REG <= io_out_ready; // @[StallRegister.scala 22:68]
    REG_1 <= ~io_out_ready; // @[StallRegister.scala 27:33]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_in_0_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_in_0_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_in_0_npc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_in_0_inst = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_in_0_fu_code = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  reg_in_0_alu_code = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  reg_in_0_jmp_code = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  reg_in_0_mem_code = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  reg_in_0_mem_size = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  reg_in_0_sys_code = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  reg_in_0_w_type = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  reg_in_0_rs1_src = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  reg_in_0_rs2_src = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  reg_in_0_rd_addr = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  reg_in_0_rd_en = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  reg_in_0_imm = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_in_0_pred_br = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  reg_in_0_pred_bpc = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  reg_in_0_rs1_paddr = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  reg_in_0_rs2_paddr = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  reg_in_0_rd_paddr = _RAND_20[5:0];
  _RAND_21 = {1{`RANDOM}};
  reg_in_0_rd_ppaddr = _RAND_21[5:0];
  _RAND_22 = {1{`RANDOM}};
  reg_in_1_valid = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  reg_in_1_pc = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  reg_in_1_npc = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  reg_in_1_inst = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  reg_in_1_fu_code = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  reg_in_1_alu_code = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  reg_in_1_jmp_code = _RAND_28[3:0];
  _RAND_29 = {1{`RANDOM}};
  reg_in_1_mem_code = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  reg_in_1_mem_size = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  reg_in_1_sys_code = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  reg_in_1_w_type = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  reg_in_1_rs1_src = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  reg_in_1_rs2_src = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  reg_in_1_rd_addr = _RAND_35[4:0];
  _RAND_36 = {1{`RANDOM}};
  reg_in_1_rd_en = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  reg_in_1_imm = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  reg_in_1_pred_br = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  reg_in_1_pred_bpc = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  reg_in_1_rs1_paddr = _RAND_40[5:0];
  _RAND_41 = {1{`RANDOM}};
  reg_in_1_rs2_paddr = _RAND_41[5:0];
  _RAND_42 = {1{`RANDOM}};
  reg_in_1_rd_paddr = _RAND_42[5:0];
  _RAND_43 = {1{`RANDOM}};
  reg_in_1_rd_ppaddr = _RAND_43[5:0];
  _RAND_44 = {1{`RANDOM}};
  reg_in_valid = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  REG = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  REG_1 = _RAND_46[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_Rob(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_vec_0_valid,
  input  [31:0] io_in_bits_vec_0_pc,
  input  [2:0]  io_in_bits_vec_0_fu_code,
  input  [2:0]  io_in_bits_vec_0_sys_code,
  input  [4:0]  io_in_bits_vec_0_rd_addr,
  input         io_in_bits_vec_0_rd_en,
  input  [5:0]  io_in_bits_vec_0_rd_paddr,
  input  [5:0]  io_in_bits_vec_0_rd_ppaddr,
  input         io_in_bits_vec_1_valid,
  input  [31:0] io_in_bits_vec_1_pc,
  input  [2:0]  io_in_bits_vec_1_fu_code,
  input  [2:0]  io_in_bits_vec_1_sys_code,
  input  [4:0]  io_in_bits_vec_1_rd_addr,
  input         io_in_bits_vec_1_rd_en,
  input  [5:0]  io_in_bits_vec_1_rd_paddr,
  input  [5:0]  io_in_bits_vec_1_rd_ppaddr,
  output [3:0]  io_rob_addr_0,
  output [3:0]  io_rob_addr_1,
  input         io_exe_0_valid,
  input  [3:0]  io_exe_0_rob_addr,
  input         io_exe_1_valid,
  input  [3:0]  io_exe_1_rob_addr,
  input         io_exe_2_valid,
  input  [3:0]  io_exe_2_rob_addr,
  input         io_exe_ecp_0_jmp_valid,
  input         io_exe_ecp_0_jmp,
  input  [31:0] io_exe_ecp_0_jmp_pc,
  input         io_exe_ecp_0_mis,
  input         io_exe_ecp_1_jmp_valid,
  input         io_exe_ecp_1_jmp,
  input  [31:0] io_exe_ecp_1_jmp_pc,
  input         io_exe_ecp_1_mis,
  input         io_exe_ecp_2_store_valid,
  output        io_cm_0_valid,
  output [4:0]  io_cm_0_rd_addr,
  output        io_cm_0_rd_en,
  output [5:0]  io_cm_0_rd_paddr,
  output [5:0]  io_cm_0_rd_ppaddr,
  output        io_cm_1_valid,
  output [4:0]  io_cm_1_rd_addr,
  output        io_cm_1_rd_en,
  output [5:0]  io_cm_1_rd_paddr,
  output [5:0]  io_cm_1_rd_ppaddr,
  output        io_jmp_packet_valid,
  output [31:0] io_jmp_packet_inst_pc,
  output        io_jmp_packet_jmp,
  output [31:0] io_jmp_packet_jmp_pc,
  output        io_jmp_packet_mis,
  output        io_jmp_packet_sys,
  output        io_sq_deq_req,
  input         io_flush,
  output        io_sys_ready,
  input         csr_mip_mtip_intr_0,
  output [63:0] intr_mcause_0,
  output [63:0] intr_mstatus_0,
  input  [29:0] csr_mtvec_idx_0,
  input         csr_mie_mtie_0,
  output        intr_0,
  input  [63:0] csr_mstatus_0,
  output [63:0] intr_mepc_0
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] rob_pc [0:15]; // @[Rob.scala 44:24]
//   wire  rob_pc_MPORT_2_en; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_2_addr; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_2_data; // @[Rob.scala 44:24]
//   wire  rob_pc_MPORT_3_en; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_3_addr; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_3_data; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_1_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_1_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_1_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_1_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_4_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_4_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_4_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_4_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_5_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_5_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_5_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_5_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_6_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_6_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_6_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_6_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_7_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_7_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_7_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_7_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_8_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_8_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_8_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_8_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_9_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_9_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_9_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_9_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_10_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_10_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_10_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_10_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_11_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_11_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_11_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_11_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_12_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_12_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_12_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_12_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_13_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_13_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_13_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_13_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_14_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_14_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_14_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_14_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_15_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_15_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_15_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_15_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_16_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_16_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_16_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_16_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_17_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_17_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_17_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_17_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_18_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_18_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_18_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_18_en; // @[Rob.scala 44:24]
  wire [31:0] rob_pc_MPORT_19_data; // @[Rob.scala 44:24]
  wire [3:0] rob_pc_MPORT_19_addr; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_19_mask; // @[Rob.scala 44:24]
  wire  rob_pc_MPORT_19_en; // @[Rob.scala 44:24]
//   reg  rob_pc_MPORT_2_en_pipe_0;
  reg [3:0] rob_pc_MPORT_2_addr_pipe_0;
//   reg  rob_pc_MPORT_3_en_pipe_0;
  reg [3:0] rob_pc_MPORT_3_addr_pipe_0;
  reg [2:0] rob_fu_code [0:15]; // @[Rob.scala 44:24]
//   wire  rob_fu_code_MPORT_2_en; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_2_addr; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_2_data; // @[Rob.scala 44:24]
//   wire  rob_fu_code_MPORT_3_en; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_3_addr; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_3_data; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_1_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_1_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_1_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_1_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_4_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_4_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_4_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_4_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_5_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_5_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_5_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_5_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_6_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_6_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_6_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_6_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_7_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_7_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_7_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_7_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_8_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_8_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_8_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_8_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_9_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_9_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_9_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_9_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_10_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_10_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_10_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_10_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_11_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_11_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_11_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_11_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_12_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_12_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_12_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_12_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_13_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_13_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_13_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_13_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_14_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_14_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_14_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_14_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_15_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_15_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_15_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_15_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_16_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_16_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_16_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_16_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_17_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_17_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_17_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_17_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_18_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_18_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_18_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_18_en; // @[Rob.scala 44:24]
  wire [2:0] rob_fu_code_MPORT_19_data; // @[Rob.scala 44:24]
  wire [3:0] rob_fu_code_MPORT_19_addr; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_19_mask; // @[Rob.scala 44:24]
  wire  rob_fu_code_MPORT_19_en; // @[Rob.scala 44:24]
//   reg  rob_fu_code_MPORT_2_en_pipe_0;
  reg [3:0] rob_fu_code_MPORT_2_addr_pipe_0;
//   reg  rob_fu_code_MPORT_3_en_pipe_0;
  reg [3:0] rob_fu_code_MPORT_3_addr_pipe_0;
  reg [2:0] rob_sys_code [0:15]; // @[Rob.scala 44:24]
//   wire  rob_sys_code_MPORT_2_en; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_2_addr; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_2_data; // @[Rob.scala 44:24]
//   wire  rob_sys_code_MPORT_3_en; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_3_addr; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_3_data; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_1_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_1_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_1_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_1_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_4_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_4_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_4_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_4_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_5_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_5_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_5_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_5_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_6_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_6_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_6_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_6_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_7_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_7_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_7_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_7_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_8_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_8_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_8_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_8_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_9_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_9_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_9_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_9_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_10_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_10_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_10_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_10_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_11_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_11_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_11_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_11_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_12_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_12_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_12_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_12_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_13_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_13_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_13_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_13_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_14_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_14_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_14_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_14_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_15_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_15_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_15_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_15_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_16_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_16_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_16_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_16_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_17_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_17_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_17_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_17_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_18_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_18_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_18_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_18_en; // @[Rob.scala 44:24]
  wire [2:0] rob_sys_code_MPORT_19_data; // @[Rob.scala 44:24]
  wire [3:0] rob_sys_code_MPORT_19_addr; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_19_mask; // @[Rob.scala 44:24]
  wire  rob_sys_code_MPORT_19_en; // @[Rob.scala 44:24]
//   reg  rob_sys_code_MPORT_2_en_pipe_0;
  reg [3:0] rob_sys_code_MPORT_2_addr_pipe_0;
//   reg  rob_sys_code_MPORT_3_en_pipe_0;
  reg [3:0] rob_sys_code_MPORT_3_addr_pipe_0;
  reg [4:0] rob_rd_addr [0:15]; // @[Rob.scala 44:24]
//   wire  rob_rd_addr_MPORT_2_en; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_2_addr; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_2_data; // @[Rob.scala 44:24]
//   wire  rob_rd_addr_MPORT_3_en; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_3_addr; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_3_data; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_1_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_1_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_1_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_1_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_4_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_4_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_4_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_4_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_5_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_5_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_5_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_5_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_6_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_6_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_6_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_6_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_7_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_7_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_7_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_7_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_8_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_8_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_8_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_8_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_9_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_9_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_9_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_9_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_10_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_10_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_10_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_10_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_11_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_11_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_11_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_11_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_12_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_12_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_12_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_12_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_13_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_13_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_13_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_13_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_14_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_14_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_14_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_14_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_15_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_15_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_15_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_15_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_16_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_16_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_16_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_16_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_17_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_17_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_17_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_17_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_18_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_18_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_18_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_18_en; // @[Rob.scala 44:24]
  wire [4:0] rob_rd_addr_MPORT_19_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_addr_MPORT_19_addr; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_19_mask; // @[Rob.scala 44:24]
  wire  rob_rd_addr_MPORT_19_en; // @[Rob.scala 44:24]
//   reg  rob_rd_addr_MPORT_2_en_pipe_0;
  reg [3:0] rob_rd_addr_MPORT_2_addr_pipe_0;
//   reg  rob_rd_addr_MPORT_3_en_pipe_0;
  reg [3:0] rob_rd_addr_MPORT_3_addr_pipe_0;
  reg  rob_rd_en [0:15]; // @[Rob.scala 44:24]
//   wire  rob_rd_en_MPORT_2_en; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_2_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_2_data; // @[Rob.scala 44:24]
//   wire  rob_rd_en_MPORT_3_en; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_3_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_3_data; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_1_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_1_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_1_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_1_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_4_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_4_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_4_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_4_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_5_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_5_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_5_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_5_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_6_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_6_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_6_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_6_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_7_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_7_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_7_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_7_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_8_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_8_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_8_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_8_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_9_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_9_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_9_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_9_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_10_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_10_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_10_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_10_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_11_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_11_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_11_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_11_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_12_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_12_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_12_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_12_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_13_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_13_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_13_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_13_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_14_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_14_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_14_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_14_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_15_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_15_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_15_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_15_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_16_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_16_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_16_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_16_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_17_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_17_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_17_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_17_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_18_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_18_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_18_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_18_en; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_19_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_en_MPORT_19_addr; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_19_mask; // @[Rob.scala 44:24]
  wire  rob_rd_en_MPORT_19_en; // @[Rob.scala 44:24]
//   reg  rob_rd_en_MPORT_2_en_pipe_0;
  reg [3:0] rob_rd_en_MPORT_2_addr_pipe_0;
//   reg  rob_rd_en_MPORT_3_en_pipe_0;
  reg [3:0] rob_rd_en_MPORT_3_addr_pipe_0;
  reg [5:0] rob_rd_paddr [0:15]; // @[Rob.scala 44:24]
//   wire  rob_rd_paddr_MPORT_2_en; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_2_addr; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_2_data; // @[Rob.scala 44:24]
//   wire  rob_rd_paddr_MPORT_3_en; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_3_addr; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_3_data; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_1_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_1_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_1_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_1_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_4_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_4_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_4_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_4_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_5_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_5_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_5_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_5_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_6_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_6_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_6_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_6_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_7_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_7_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_7_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_7_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_8_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_8_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_8_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_8_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_9_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_9_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_9_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_9_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_10_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_10_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_10_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_10_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_11_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_11_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_11_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_11_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_12_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_12_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_12_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_12_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_13_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_13_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_13_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_13_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_14_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_14_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_14_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_14_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_15_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_15_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_15_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_15_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_16_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_16_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_16_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_16_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_17_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_17_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_17_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_17_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_18_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_18_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_18_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_18_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_paddr_MPORT_19_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_paddr_MPORT_19_addr; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_19_mask; // @[Rob.scala 44:24]
  wire  rob_rd_paddr_MPORT_19_en; // @[Rob.scala 44:24]
//   reg  rob_rd_paddr_MPORT_2_en_pipe_0;
  reg [3:0] rob_rd_paddr_MPORT_2_addr_pipe_0;
//   reg  rob_rd_paddr_MPORT_3_en_pipe_0;
  reg [3:0] rob_rd_paddr_MPORT_3_addr_pipe_0;
  reg [5:0] rob_rd_ppaddr [0:15]; // @[Rob.scala 44:24]
//   wire  rob_rd_ppaddr_MPORT_2_en; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_2_addr; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_2_data; // @[Rob.scala 44:24]
//   wire  rob_rd_ppaddr_MPORT_3_en; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_3_addr; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_3_data; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_1_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_1_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_1_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_1_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_4_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_4_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_4_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_4_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_5_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_5_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_5_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_5_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_6_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_6_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_6_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_6_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_7_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_7_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_7_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_7_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_8_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_8_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_8_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_8_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_9_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_9_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_9_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_9_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_10_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_10_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_10_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_10_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_11_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_11_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_11_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_11_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_12_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_12_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_12_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_12_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_13_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_13_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_13_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_13_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_14_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_14_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_14_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_14_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_15_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_15_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_15_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_15_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_16_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_16_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_16_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_16_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_17_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_17_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_17_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_17_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_18_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_18_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_18_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_18_en; // @[Rob.scala 44:24]
  wire [5:0] rob_rd_ppaddr_MPORT_19_data; // @[Rob.scala 44:24]
  wire [3:0] rob_rd_ppaddr_MPORT_19_addr; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_19_mask; // @[Rob.scala 44:24]
  wire  rob_rd_ppaddr_MPORT_19_en; // @[Rob.scala 44:24]
//   reg  rob_rd_ppaddr_MPORT_2_en_pipe_0;
  reg [3:0] rob_rd_ppaddr_MPORT_2_addr_pipe_0;
//   reg  rob_rd_ppaddr_MPORT_3_en_pipe_0;
  reg [3:0] rob_rd_ppaddr_MPORT_3_addr_pipe_0;
  reg [4:0] enq_vec_0; // @[Rob.scala 46:24]
  reg [4:0] enq_vec_1; // @[Rob.scala 46:24]
  reg [4:0] deq_vec_0; // @[Rob.scala 47:24]
  reg [4:0] deq_vec_1; // @[Rob.scala 47:24]
  wire [3:0] enq_ptr = enq_vec_0[3:0]; // @[Rob.scala 17:32]
  wire [3:0] deq_ptr = deq_vec_0[3:0]; // @[Rob.scala 17:32]
  wire  enq_flag = enq_vec_0[4]; // @[Rob.scala 18:33]
  wire  deq_flag = deq_vec_0[4]; // @[Rob.scala 18:33]
  wire  _T_2 = enq_flag == deq_flag; // @[Rob.scala 53:28]
  wire [3:0] _T_4 = enq_ptr - deq_ptr; // @[Rob.scala 53:50]
  wire [4:0] _GEN_2222 = {{1'd0}, enq_ptr}; // @[Rob.scala 53:71]
  wire [4:0] _T_6 = 5'h10 + _GEN_2222; // @[Rob.scala 53:71]
  wire [4:0] _GEN_2223 = {{1'd0}, deq_ptr}; // @[Rob.scala 53:81]
  wire [4:0] _T_8 = _T_6 - _GEN_2223; // @[Rob.scala 53:81]
  wire [4:0] count = enq_flag == deq_flag ? {{1'd0}, _T_4} : _T_8; // @[Rob.scala 53:18]
  wire  rob_empty = _T_2 & enq_ptr == deq_ptr; // @[Rob.scala 54:43]
  wire  _T_11 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_12 = io_in_bits_vec_0_valid + io_in_bits_vec_1_valid; // @[Bitwise.scala 47:55]
  wire [1:0] num_enq = _T_11 ? _T_12 : 2'h0; // @[Rob.scala 56:20]
  wire  shiftAmount = count[0]; // @[OneHot.scala 64:49]
  wire [1:0] _T_36 = 2'h1 << shiftAmount; // @[OneHot.scala 65:12]
  wire [1:0] _T_39 = _T_36 - 2'h1; // @[Rob.scala 121:98]
  wire [1:0] valid_vec = count >= 5'h2 ? 2'h3 : _T_39; // @[Rob.scala 121:22]
  reg  complete_15; // @[Rob.scala 70:25]
  reg  complete_14; // @[Rob.scala 70:25]
  reg  complete_13; // @[Rob.scala 70:25]
  reg  complete_12; // @[Rob.scala 70:25]
  reg  complete_11; // @[Rob.scala 70:25]
  reg  complete_10; // @[Rob.scala 70:25]
  reg  complete_9; // @[Rob.scala 70:25]
  reg  complete_8; // @[Rob.scala 70:25]
  reg  complete_7; // @[Rob.scala 70:25]
  reg  complete_6; // @[Rob.scala 70:25]
  reg  complete_5; // @[Rob.scala 70:25]
  reg  complete_4; // @[Rob.scala 70:25]
  reg  complete_3; // @[Rob.scala 70:25]
  reg  complete_2; // @[Rob.scala 70:25]
  reg  complete_1; // @[Rob.scala 70:25]
  reg  complete_0; // @[Rob.scala 70:25]
  wire  _GEN_1347 = 4'h1 == deq_ptr ? complete_1 : complete_0; // @[Rob.scala 131:{24,24}]
  wire  _GEN_1348 = 4'h2 == deq_ptr ? complete_2 : _GEN_1347; // @[Rob.scala 131:{24,24}]
  wire  _GEN_1349 = 4'h3 == deq_ptr ? complete_3 : _GEN_1348; // @[Rob.scala 131:{24,24}]
  wire  _GEN_1350 = 4'h4 == deq_ptr ? complete_4 : _GEN_1349; // @[Rob.scala 131:{24,24}]
  wire  _GEN_1351 = 4'h5 == deq_ptr ? complete_5 : _GEN_1350; // @[Rob.scala 131:{24,24}]
  wire  _GEN_1352 = 4'h6 == deq_ptr ? complete_6 : _GEN_1351; // @[Rob.scala 131:{24,24}]
  wire  _GEN_1353 = 4'h7 == deq_ptr ? complete_7 : _GEN_1352; // @[Rob.scala 131:{24,24}]
  wire  _GEN_1354 = 4'h8 == deq_ptr ? complete_8 : _GEN_1353; // @[Rob.scala 131:{24,24}]
  wire  _GEN_1355 = 4'h9 == deq_ptr ? complete_9 : _GEN_1354; // @[Rob.scala 131:{24,24}]
  wire  _GEN_1356 = 4'ha == deq_ptr ? complete_10 : _GEN_1355; // @[Rob.scala 131:{24,24}]
  wire  _GEN_1357 = 4'hb == deq_ptr ? complete_11 : _GEN_1356; // @[Rob.scala 131:{24,24}]
  wire  _GEN_1358 = 4'hc == deq_ptr ? complete_12 : _GEN_1357; // @[Rob.scala 131:{24,24}]
  wire  _GEN_1359 = 4'hd == deq_ptr ? complete_13 : _GEN_1358; // @[Rob.scala 131:{24,24}]
  wire  _GEN_1360 = 4'he == deq_ptr ? complete_14 : _GEN_1359; // @[Rob.scala 131:{24,24}]
  wire  complete_mask_0 = 4'hf == deq_ptr ? complete_15 : _GEN_1360; // @[Rob.scala 131:{24,24}]
  wire  cm_0_valid = valid_vec[0] & complete_mask_0; // @[Rob.scala 257:35]
  wire  _GEN_1363 = 4'h1 == deq_vec_1[3:0] ? complete_1 : complete_0; // @[Rob.scala 133:{48,48}]
  wire  _GEN_1364 = 4'h2 == deq_vec_1[3:0] ? complete_2 : _GEN_1363; // @[Rob.scala 133:{48,48}]
  wire  _GEN_1365 = 4'h3 == deq_vec_1[3:0] ? complete_3 : _GEN_1364; // @[Rob.scala 133:{48,48}]
  wire  _GEN_1366 = 4'h4 == deq_vec_1[3:0] ? complete_4 : _GEN_1365; // @[Rob.scala 133:{48,48}]
  wire  _GEN_1367 = 4'h5 == deq_vec_1[3:0] ? complete_5 : _GEN_1366; // @[Rob.scala 133:{48,48}]
  wire  _GEN_1368 = 4'h6 == deq_vec_1[3:0] ? complete_6 : _GEN_1367; // @[Rob.scala 133:{48,48}]
  wire  _GEN_1369 = 4'h7 == deq_vec_1[3:0] ? complete_7 : _GEN_1368; // @[Rob.scala 133:{48,48}]
  wire  _GEN_1370 = 4'h8 == deq_vec_1[3:0] ? complete_8 : _GEN_1369; // @[Rob.scala 133:{48,48}]
  wire  _GEN_1371 = 4'h9 == deq_vec_1[3:0] ? complete_9 : _GEN_1370; // @[Rob.scala 133:{48,48}]
  wire  _GEN_1372 = 4'ha == deq_vec_1[3:0] ? complete_10 : _GEN_1371; // @[Rob.scala 133:{48,48}]
  wire  _GEN_1373 = 4'hb == deq_vec_1[3:0] ? complete_11 : _GEN_1372; // @[Rob.scala 133:{48,48}]
  wire  _GEN_1374 = 4'hc == deq_vec_1[3:0] ? complete_12 : _GEN_1373; // @[Rob.scala 133:{48,48}]
  wire  _GEN_1375 = 4'hd == deq_vec_1[3:0] ? complete_13 : _GEN_1374; // @[Rob.scala 133:{48,48}]
  wire  _GEN_1376 = 4'he == deq_vec_1[3:0] ? complete_14 : _GEN_1375; // @[Rob.scala 133:{48,48}]
  wire  _GEN_1377 = 4'hf == deq_vec_1[3:0] ? complete_15 : _GEN_1376; // @[Rob.scala 133:{48,48}]
  wire  complete_mask_1 = complete_mask_0 & _GEN_1377; // @[Rob.scala 133:48]
  reg  ecp_15_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_14_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_13_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_12_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_11_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_10_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_9_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_8_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_7_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_6_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_5_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_4_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_3_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_2_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_1_jmp_valid; // @[Rob.scala 71:20]
  reg  ecp_0_jmp_valid; // @[Rob.scala 71:20]
  wire  _GEN_1472 = 4'h1 == deq_ptr ? ecp_1_jmp_valid : ecp_0_jmp_valid; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1473 = 4'h2 == deq_ptr ? ecp_2_jmp_valid : _GEN_1472; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1474 = 4'h3 == deq_ptr ? ecp_3_jmp_valid : _GEN_1473; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1475 = 4'h4 == deq_ptr ? ecp_4_jmp_valid : _GEN_1474; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1476 = 4'h5 == deq_ptr ? ecp_5_jmp_valid : _GEN_1475; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1477 = 4'h6 == deq_ptr ? ecp_6_jmp_valid : _GEN_1476; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1478 = 4'h7 == deq_ptr ? ecp_7_jmp_valid : _GEN_1477; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1479 = 4'h8 == deq_ptr ? ecp_8_jmp_valid : _GEN_1478; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1480 = 4'h9 == deq_ptr ? ecp_9_jmp_valid : _GEN_1479; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1481 = 4'ha == deq_ptr ? ecp_10_jmp_valid : _GEN_1480; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1482 = 4'hb == deq_ptr ? ecp_11_jmp_valid : _GEN_1481; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1483 = 4'hc == deq_ptr ? ecp_12_jmp_valid : _GEN_1482; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1484 = 4'hd == deq_ptr ? ecp_13_jmp_valid : _GEN_1483; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1485 = 4'he == deq_ptr ? ecp_14_jmp_valid : _GEN_1484; // @[Rob.scala 231:{16,16}]
  wire  deq_ecp_0_jmp_valid = 4'hf == deq_ptr ? ecp_15_jmp_valid : _GEN_1485; // @[Rob.scala 231:{16,16}]
  reg  ecp_15_mis; // @[Rob.scala 71:20]
  reg  ecp_14_mis; // @[Rob.scala 71:20]
  reg  ecp_13_mis; // @[Rob.scala 71:20]
  reg  ecp_12_mis; // @[Rob.scala 71:20]
  reg  ecp_11_mis; // @[Rob.scala 71:20]
  reg  ecp_10_mis; // @[Rob.scala 71:20]
  reg  ecp_9_mis; // @[Rob.scala 71:20]
  reg  ecp_8_mis; // @[Rob.scala 71:20]
  reg  ecp_7_mis; // @[Rob.scala 71:20]
  reg  ecp_6_mis; // @[Rob.scala 71:20]
  reg  ecp_5_mis; // @[Rob.scala 71:20]
  reg  ecp_4_mis; // @[Rob.scala 71:20]
  reg  ecp_3_mis; // @[Rob.scala 71:20]
  reg  ecp_2_mis; // @[Rob.scala 71:20]
  reg  ecp_1_mis; // @[Rob.scala 71:20]
  reg  ecp_0_mis; // @[Rob.scala 71:20]
  wire  _GEN_1424 = 4'h1 == deq_ptr ? ecp_1_mis : ecp_0_mis; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1425 = 4'h2 == deq_ptr ? ecp_2_mis : _GEN_1424; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1426 = 4'h3 == deq_ptr ? ecp_3_mis : _GEN_1425; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1427 = 4'h4 == deq_ptr ? ecp_4_mis : _GEN_1426; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1428 = 4'h5 == deq_ptr ? ecp_5_mis : _GEN_1427; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1429 = 4'h6 == deq_ptr ? ecp_6_mis : _GEN_1428; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1430 = 4'h7 == deq_ptr ? ecp_7_mis : _GEN_1429; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1431 = 4'h8 == deq_ptr ? ecp_8_mis : _GEN_1430; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1432 = 4'h9 == deq_ptr ? ecp_9_mis : _GEN_1431; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1433 = 4'ha == deq_ptr ? ecp_10_mis : _GEN_1432; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1434 = 4'hb == deq_ptr ? ecp_11_mis : _GEN_1433; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1435 = 4'hc == deq_ptr ? ecp_12_mis : _GEN_1434; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1436 = 4'hd == deq_ptr ? ecp_13_mis : _GEN_1435; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1437 = 4'he == deq_ptr ? ecp_14_mis : _GEN_1436; // @[Rob.scala 231:{16,16}]
  wire  deq_ecp_0_mis = 4'hf == deq_ptr ? ecp_15_mis : _GEN_1437; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1602 = 4'h1 == deq_vec_1[3:0] ? ecp_1_jmp_valid : ecp_0_jmp_valid; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1603 = 4'h2 == deq_vec_1[3:0] ? ecp_2_jmp_valid : _GEN_1602; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1604 = 4'h3 == deq_vec_1[3:0] ? ecp_3_jmp_valid : _GEN_1603; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1605 = 4'h4 == deq_vec_1[3:0] ? ecp_4_jmp_valid : _GEN_1604; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1606 = 4'h5 == deq_vec_1[3:0] ? ecp_5_jmp_valid : _GEN_1605; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1607 = 4'h6 == deq_vec_1[3:0] ? ecp_6_jmp_valid : _GEN_1606; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1608 = 4'h7 == deq_vec_1[3:0] ? ecp_7_jmp_valid : _GEN_1607; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1609 = 4'h8 == deq_vec_1[3:0] ? ecp_8_jmp_valid : _GEN_1608; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1610 = 4'h9 == deq_vec_1[3:0] ? ecp_9_jmp_valid : _GEN_1609; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1611 = 4'ha == deq_vec_1[3:0] ? ecp_10_jmp_valid : _GEN_1610; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1612 = 4'hb == deq_vec_1[3:0] ? ecp_11_jmp_valid : _GEN_1611; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1613 = 4'hc == deq_vec_1[3:0] ? ecp_12_jmp_valid : _GEN_1612; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1614 = 4'hd == deq_vec_1[3:0] ? ecp_13_jmp_valid : _GEN_1613; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1615 = 4'he == deq_vec_1[3:0] ? ecp_14_jmp_valid : _GEN_1614; // @[Rob.scala 231:{16,16}]
  wire  deq_ecp_1_jmp_valid = 4'hf == deq_vec_1[3:0] ? ecp_15_jmp_valid : _GEN_1615; // @[Rob.scala 231:{16,16}]
  wire  jmp_mask_1 = deq_ecp_0_jmp_valid ? ~deq_ecp_0_mis & ~deq_ecp_1_jmp_valid : 1'h1; // @[Rob.scala 251:25]
  reg  ecp_15_store_valid; // @[Rob.scala 71:20]
  reg  ecp_14_store_valid; // @[Rob.scala 71:20]
  reg  ecp_13_store_valid; // @[Rob.scala 71:20]
  reg  ecp_12_store_valid; // @[Rob.scala 71:20]
  reg  ecp_11_store_valid; // @[Rob.scala 71:20]
  reg  ecp_10_store_valid; // @[Rob.scala 71:20]
  reg  ecp_9_store_valid; // @[Rob.scala 71:20]
  reg  ecp_8_store_valid; // @[Rob.scala 71:20]
  reg  ecp_7_store_valid; // @[Rob.scala 71:20]
  reg  ecp_6_store_valid; // @[Rob.scala 71:20]
  reg  ecp_5_store_valid; // @[Rob.scala 71:20]
  reg  ecp_4_store_valid; // @[Rob.scala 71:20]
  reg  ecp_3_store_valid; // @[Rob.scala 71:20]
  reg  ecp_2_store_valid; // @[Rob.scala 71:20]
  reg  ecp_1_store_valid; // @[Rob.scala 71:20]
  reg  ecp_0_store_valid; // @[Rob.scala 71:20]
  wire  _GEN_1504 = 4'h1 == deq_ptr ? ecp_1_store_valid : ecp_0_store_valid; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1505 = 4'h2 == deq_ptr ? ecp_2_store_valid : _GEN_1504; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1506 = 4'h3 == deq_ptr ? ecp_3_store_valid : _GEN_1505; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1507 = 4'h4 == deq_ptr ? ecp_4_store_valid : _GEN_1506; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1508 = 4'h5 == deq_ptr ? ecp_5_store_valid : _GEN_1507; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1509 = 4'h6 == deq_ptr ? ecp_6_store_valid : _GEN_1508; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1510 = 4'h7 == deq_ptr ? ecp_7_store_valid : _GEN_1509; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1511 = 4'h8 == deq_ptr ? ecp_8_store_valid : _GEN_1510; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1512 = 4'h9 == deq_ptr ? ecp_9_store_valid : _GEN_1511; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1513 = 4'ha == deq_ptr ? ecp_10_store_valid : _GEN_1512; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1514 = 4'hb == deq_ptr ? ecp_11_store_valid : _GEN_1513; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1515 = 4'hc == deq_ptr ? ecp_12_store_valid : _GEN_1514; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1516 = 4'hd == deq_ptr ? ecp_13_store_valid : _GEN_1515; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1517 = 4'he == deq_ptr ? ecp_14_store_valid : _GEN_1516; // @[Rob.scala 231:{16,16}]
  wire  deq_ecp_0_store_valid = 4'hf == deq_ptr ? ecp_15_store_valid : _GEN_1517; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1634 = 4'h1 == deq_vec_1[3:0] ? ecp_1_store_valid : ecp_0_store_valid; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1635 = 4'h2 == deq_vec_1[3:0] ? ecp_2_store_valid : _GEN_1634; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1636 = 4'h3 == deq_vec_1[3:0] ? ecp_3_store_valid : _GEN_1635; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1637 = 4'h4 == deq_vec_1[3:0] ? ecp_4_store_valid : _GEN_1636; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1638 = 4'h5 == deq_vec_1[3:0] ? ecp_5_store_valid : _GEN_1637; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1639 = 4'h6 == deq_vec_1[3:0] ? ecp_6_store_valid : _GEN_1638; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1640 = 4'h7 == deq_vec_1[3:0] ? ecp_7_store_valid : _GEN_1639; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1641 = 4'h8 == deq_vec_1[3:0] ? ecp_8_store_valid : _GEN_1640; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1642 = 4'h9 == deq_vec_1[3:0] ? ecp_9_store_valid : _GEN_1641; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1643 = 4'ha == deq_vec_1[3:0] ? ecp_10_store_valid : _GEN_1642; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1644 = 4'hb == deq_vec_1[3:0] ? ecp_11_store_valid : _GEN_1643; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1645 = 4'hc == deq_vec_1[3:0] ? ecp_12_store_valid : _GEN_1644; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1646 = 4'hd == deq_vec_1[3:0] ? ecp_13_store_valid : _GEN_1645; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1647 = 4'he == deq_vec_1[3:0] ? ecp_14_store_valid : _GEN_1646; // @[Rob.scala 231:{16,16}]
  wire  deq_ecp_1_store_valid = 4'hf == deq_vec_1[3:0] ? ecp_15_store_valid : _GEN_1647; // @[Rob.scala 231:{16,16}]
  wire  store_mask_1 = deq_ecp_0_store_valid ? ~deq_ecp_1_store_valid : 1'h1; // @[Rob.scala 252:27]
  wire  deq_uop_0_rd_en = rob_rd_en_MPORT_2_data; // @[Rob.scala 156:21 229:16]
  wire  deq_uop_1_rd_en = rob_rd_en_MPORT_3_data; // @[Rob.scala 156:21 229:16]
  wire [4:0] deq_uop_0_rd_addr = rob_rd_addr_MPORT_2_data; // @[Rob.scala 156:21 229:16]
  wire [4:0] deq_uop_1_rd_addr = rob_rd_addr_MPORT_3_data; // @[Rob.scala 156:21 229:16]
  wire  _T_115 = cm_0_valid & deq_uop_0_rd_en & deq_uop_1_rd_en ? deq_uop_0_rd_addr != deq_uop_1_rd_addr : 1'h1; // @[Rob.scala 261:28]
  wire  cm_1_valid = valid_vec[1] & complete_mask_1 & jmp_mask_1 & store_mask_1 & _T_115; // @[Rob.scala 260:87]
  wire [1:0] num_deq = cm_0_valid + cm_1_valid; // @[Bitwise.scala 47:55]
  wire [4:0] _GEN_2224 = {{3'd0}, num_enq}; // @[Rob.scala 61:29]
  wire [5:0] next_valid_entry = count + _GEN_2224; // @[Rob.scala 61:29]
  reg  enq_ready; // @[Rob.scala 65:26]
  reg  ecp_0_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_0_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_1_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_1_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_2_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_2_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_3_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_3_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_4_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_4_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_5_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_5_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_6_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_6_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_7_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_7_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_8_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_8_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_9_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_9_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_10_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_10_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_11_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_11_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_12_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_12_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_13_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_13_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_14_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_14_jmp_pc; // @[Rob.scala 71:20]
  reg  ecp_15_jmp; // @[Rob.scala 71:20]
  reg [31:0] ecp_15_jmp_pc; // @[Rob.scala 71:20]
  wire  _T_20 = io_in_bits_vec_0_valid & _T_11; // @[Rob.scala 91:35]
  wire  _T_21 = ~io_flush; // @[Rob.scala 91:54]
  wire  _GEN_2 = 4'h0 == enq_ptr ? 1'h0 : complete_0; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_3 = 4'h1 == enq_ptr ? 1'h0 : complete_1; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_4 = 4'h2 == enq_ptr ? 1'h0 : complete_2; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_5 = 4'h3 == enq_ptr ? 1'h0 : complete_3; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_6 = 4'h4 == enq_ptr ? 1'h0 : complete_4; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_7 = 4'h5 == enq_ptr ? 1'h0 : complete_5; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_8 = 4'h6 == enq_ptr ? 1'h0 : complete_6; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_9 = 4'h7 == enq_ptr ? 1'h0 : complete_7; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_10 = 4'h8 == enq_ptr ? 1'h0 : complete_8; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_11 = 4'h9 == enq_ptr ? 1'h0 : complete_9; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_12 = 4'ha == enq_ptr ? 1'h0 : complete_10; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_13 = 4'hb == enq_ptr ? 1'h0 : complete_11; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_14 = 4'hc == enq_ptr ? 1'h0 : complete_12; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_15 = 4'hd == enq_ptr ? 1'h0 : complete_13; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_16 = 4'he == enq_ptr ? 1'h0 : complete_14; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_17 = 4'hf == enq_ptr ? 1'h0 : complete_15; // @[Rob.scala 70:25 93:{25,25}]
  wire  _GEN_34 = 4'h0 == enq_ptr ? 1'h0 : ecp_0_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_35 = 4'h1 == enq_ptr ? 1'h0 : ecp_1_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_36 = 4'h2 == enq_ptr ? 1'h0 : ecp_2_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_37 = 4'h3 == enq_ptr ? 1'h0 : ecp_3_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_38 = 4'h4 == enq_ptr ? 1'h0 : ecp_4_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_39 = 4'h5 == enq_ptr ? 1'h0 : ecp_5_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_40 = 4'h6 == enq_ptr ? 1'h0 : ecp_6_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_41 = 4'h7 == enq_ptr ? 1'h0 : ecp_7_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_42 = 4'h8 == enq_ptr ? 1'h0 : ecp_8_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_43 = 4'h9 == enq_ptr ? 1'h0 : ecp_9_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_44 = 4'ha == enq_ptr ? 1'h0 : ecp_10_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_45 = 4'hb == enq_ptr ? 1'h0 : ecp_11_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_46 = 4'hc == enq_ptr ? 1'h0 : ecp_12_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_47 = 4'hd == enq_ptr ? 1'h0 : ecp_13_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_48 = 4'he == enq_ptr ? 1'h0 : ecp_14_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_49 = 4'hf == enq_ptr ? 1'h0 : ecp_15_mis; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_50 = 4'h0 == enq_ptr ? 32'h0 : ecp_0_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_51 = 4'h1 == enq_ptr ? 32'h0 : ecp_1_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_52 = 4'h2 == enq_ptr ? 32'h0 : ecp_2_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_53 = 4'h3 == enq_ptr ? 32'h0 : ecp_3_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_54 = 4'h4 == enq_ptr ? 32'h0 : ecp_4_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_55 = 4'h5 == enq_ptr ? 32'h0 : ecp_5_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_56 = 4'h6 == enq_ptr ? 32'h0 : ecp_6_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_57 = 4'h7 == enq_ptr ? 32'h0 : ecp_7_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_58 = 4'h8 == enq_ptr ? 32'h0 : ecp_8_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_59 = 4'h9 == enq_ptr ? 32'h0 : ecp_9_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_60 = 4'ha == enq_ptr ? 32'h0 : ecp_10_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_61 = 4'hb == enq_ptr ? 32'h0 : ecp_11_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_62 = 4'hc == enq_ptr ? 32'h0 : ecp_12_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_63 = 4'hd == enq_ptr ? 32'h0 : ecp_13_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_64 = 4'he == enq_ptr ? 32'h0 : ecp_14_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire [31:0] _GEN_65 = 4'hf == enq_ptr ? 32'h0 : ecp_15_jmp_pc; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_66 = 4'h0 == enq_ptr ? 1'h0 : ecp_0_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_67 = 4'h1 == enq_ptr ? 1'h0 : ecp_1_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_68 = 4'h2 == enq_ptr ? 1'h0 : ecp_2_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_69 = 4'h3 == enq_ptr ? 1'h0 : ecp_3_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_70 = 4'h4 == enq_ptr ? 1'h0 : ecp_4_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_71 = 4'h5 == enq_ptr ? 1'h0 : ecp_5_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_72 = 4'h6 == enq_ptr ? 1'h0 : ecp_6_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_73 = 4'h7 == enq_ptr ? 1'h0 : ecp_7_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_74 = 4'h8 == enq_ptr ? 1'h0 : ecp_8_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_75 = 4'h9 == enq_ptr ? 1'h0 : ecp_9_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_76 = 4'ha == enq_ptr ? 1'h0 : ecp_10_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_77 = 4'hb == enq_ptr ? 1'h0 : ecp_11_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_78 = 4'hc == enq_ptr ? 1'h0 : ecp_12_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_79 = 4'hd == enq_ptr ? 1'h0 : ecp_13_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_80 = 4'he == enq_ptr ? 1'h0 : ecp_14_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_81 = 4'hf == enq_ptr ? 1'h0 : ecp_15_jmp; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_82 = 4'h0 == enq_ptr ? 1'h0 : ecp_0_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_83 = 4'h1 == enq_ptr ? 1'h0 : ecp_1_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_84 = 4'h2 == enq_ptr ? 1'h0 : ecp_2_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_85 = 4'h3 == enq_ptr ? 1'h0 : ecp_3_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_86 = 4'h4 == enq_ptr ? 1'h0 : ecp_4_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_87 = 4'h5 == enq_ptr ? 1'h0 : ecp_5_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_88 = 4'h6 == enq_ptr ? 1'h0 : ecp_6_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_89 = 4'h7 == enq_ptr ? 1'h0 : ecp_7_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_90 = 4'h8 == enq_ptr ? 1'h0 : ecp_8_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_91 = 4'h9 == enq_ptr ? 1'h0 : ecp_9_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_92 = 4'ha == enq_ptr ? 1'h0 : ecp_10_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_93 = 4'hb == enq_ptr ? 1'h0 : ecp_11_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_94 = 4'hc == enq_ptr ? 1'h0 : ecp_12_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_95 = 4'hd == enq_ptr ? 1'h0 : ecp_13_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_96 = 4'he == enq_ptr ? 1'h0 : ecp_14_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_97 = 4'hf == enq_ptr ? 1'h0 : ecp_15_jmp_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_114 = 4'h0 == enq_ptr ? 1'h0 : ecp_0_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_115 = 4'h1 == enq_ptr ? 1'h0 : ecp_1_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_116 = 4'h2 == enq_ptr ? 1'h0 : ecp_2_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_117 = 4'h3 == enq_ptr ? 1'h0 : ecp_3_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_118 = 4'h4 == enq_ptr ? 1'h0 : ecp_4_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_119 = 4'h5 == enq_ptr ? 1'h0 : ecp_5_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_120 = 4'h6 == enq_ptr ? 1'h0 : ecp_6_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_121 = 4'h7 == enq_ptr ? 1'h0 : ecp_7_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_122 = 4'h8 == enq_ptr ? 1'h0 : ecp_8_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_123 = 4'h9 == enq_ptr ? 1'h0 : ecp_9_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_124 = 4'ha == enq_ptr ? 1'h0 : ecp_10_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_125 = 4'hb == enq_ptr ? 1'h0 : ecp_11_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_126 = 4'hc == enq_ptr ? 1'h0 : ecp_12_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_127 = 4'hd == enq_ptr ? 1'h0 : ecp_13_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_128 = 4'he == enq_ptr ? 1'h0 : ecp_14_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_129 = 4'hf == enq_ptr ? 1'h0 : ecp_15_store_valid; // @[Rob.scala 71:20 94:{20,20}]
  wire  _GEN_159 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_2 : complete_0; // @[Rob.scala 70:25 91:65]
  wire  _GEN_160 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_3 : complete_1; // @[Rob.scala 70:25 91:65]
  wire  _GEN_161 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_4 : complete_2; // @[Rob.scala 70:25 91:65]
  wire  _GEN_162 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_5 : complete_3; // @[Rob.scala 70:25 91:65]
  wire  _GEN_163 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_6 : complete_4; // @[Rob.scala 70:25 91:65]
  wire  _GEN_164 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_7 : complete_5; // @[Rob.scala 70:25 91:65]
  wire  _GEN_165 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_8 : complete_6; // @[Rob.scala 70:25 91:65]
  wire  _GEN_166 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_9 : complete_7; // @[Rob.scala 70:25 91:65]
  wire  _GEN_167 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_10 : complete_8; // @[Rob.scala 70:25 91:65]
  wire  _GEN_168 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_11 : complete_9; // @[Rob.scala 70:25 91:65]
  wire  _GEN_169 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_12 : complete_10; // @[Rob.scala 70:25 91:65]
  wire  _GEN_170 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_13 : complete_11; // @[Rob.scala 70:25 91:65]
  wire  _GEN_171 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_14 : complete_12; // @[Rob.scala 70:25 91:65]
  wire  _GEN_172 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_15 : complete_13; // @[Rob.scala 70:25 91:65]
  wire  _GEN_173 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_16 : complete_14; // @[Rob.scala 70:25 91:65]
  wire  _GEN_174 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_17 : complete_15; // @[Rob.scala 70:25 91:65]
  wire  _GEN_191 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_34 : ecp_0_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_192 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_35 : ecp_1_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_193 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_36 : ecp_2_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_194 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_37 : ecp_3_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_195 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_38 : ecp_4_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_196 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_39 : ecp_5_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_197 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_40 : ecp_6_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_198 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_41 : ecp_7_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_199 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_42 : ecp_8_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_200 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_43 : ecp_9_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_201 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_44 : ecp_10_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_202 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_45 : ecp_11_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_203 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_46 : ecp_12_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_204 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_47 : ecp_13_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_205 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_48 : ecp_14_mis; // @[Rob.scala 71:20 91:65]
  wire  _GEN_206 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_49 : ecp_15_mis; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_207 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_50 : ecp_0_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_208 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_51 : ecp_1_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_209 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_52 : ecp_2_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_210 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_53 : ecp_3_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_211 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_54 : ecp_4_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_212 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_55 : ecp_5_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_213 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_56 : ecp_6_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_214 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_57 : ecp_7_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_215 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_58 : ecp_8_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_216 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_59 : ecp_9_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_217 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_60 : ecp_10_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_218 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_61 : ecp_11_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_219 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_62 : ecp_12_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_220 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_63 : ecp_13_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_221 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_64 : ecp_14_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire [31:0] _GEN_222 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_65 : ecp_15_jmp_pc; // @[Rob.scala 71:20 91:65]
  wire  _GEN_223 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_66 : ecp_0_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_224 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_67 : ecp_1_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_225 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_68 : ecp_2_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_226 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_69 : ecp_3_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_227 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_70 : ecp_4_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_228 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_71 : ecp_5_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_229 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_72 : ecp_6_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_230 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_73 : ecp_7_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_231 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_74 : ecp_8_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_232 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_75 : ecp_9_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_233 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_76 : ecp_10_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_234 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_77 : ecp_11_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_235 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_78 : ecp_12_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_236 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_79 : ecp_13_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_237 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_80 : ecp_14_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_238 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_81 : ecp_15_jmp; // @[Rob.scala 71:20 91:65]
  wire  _GEN_239 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_82 : ecp_0_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_240 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_83 : ecp_1_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_241 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_84 : ecp_2_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_242 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_85 : ecp_3_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_243 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_86 : ecp_4_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_244 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_87 : ecp_5_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_245 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_88 : ecp_6_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_246 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_89 : ecp_7_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_247 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_90 : ecp_8_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_248 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_91 : ecp_9_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_249 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_92 : ecp_10_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_250 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_93 : ecp_11_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_251 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_94 : ecp_12_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_252 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_95 : ecp_13_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_253 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_96 : ecp_14_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_254 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_97 : ecp_15_jmp_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_271 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_114 : ecp_0_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_272 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_115 : ecp_1_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_273 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_116 : ecp_2_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_274 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_117 : ecp_3_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_275 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_118 : ecp_4_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_276 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_119 : ecp_5_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_277 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_120 : ecp_6_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_278 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_121 : ecp_7_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_279 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_122 : ecp_8_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_280 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_123 : ecp_9_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_281 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_124 : ecp_10_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_282 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_125 : ecp_11_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_283 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_126 : ecp_12_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_284 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_127 : ecp_13_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_285 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_128 : ecp_14_store_valid; // @[Rob.scala 71:20 91:65]
  wire  _GEN_286 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? _GEN_129 : ecp_15_store_valid; // @[Rob.scala 71:20 91:65]
  wire [4:0] _GEN_289 = io_in_bits_vec_0_valid ? enq_vec_1 : enq_vec_0; // @[Rob.scala 17:{32,32}]
  wire  _T_25 = io_in_bits_vec_1_valid & _T_11; // @[Rob.scala 91:35]
  wire  _GEN_290 = 4'h0 == _GEN_289[3:0] ? 1'h0 : _GEN_159; // @[Rob.scala 93:{25,25}]
  wire  _GEN_291 = 4'h1 == _GEN_289[3:0] ? 1'h0 : _GEN_160; // @[Rob.scala 93:{25,25}]
  wire  _GEN_292 = 4'h2 == _GEN_289[3:0] ? 1'h0 : _GEN_161; // @[Rob.scala 93:{25,25}]
  wire  _GEN_293 = 4'h3 == _GEN_289[3:0] ? 1'h0 : _GEN_162; // @[Rob.scala 93:{25,25}]
  wire  _GEN_294 = 4'h4 == _GEN_289[3:0] ? 1'h0 : _GEN_163; // @[Rob.scala 93:{25,25}]
  wire  _GEN_295 = 4'h5 == _GEN_289[3:0] ? 1'h0 : _GEN_164; // @[Rob.scala 93:{25,25}]
  wire  _GEN_296 = 4'h6 == _GEN_289[3:0] ? 1'h0 : _GEN_165; // @[Rob.scala 93:{25,25}]
  wire  _GEN_297 = 4'h7 == _GEN_289[3:0] ? 1'h0 : _GEN_166; // @[Rob.scala 93:{25,25}]
  wire  _GEN_298 = 4'h8 == _GEN_289[3:0] ? 1'h0 : _GEN_167; // @[Rob.scala 93:{25,25}]
  wire  _GEN_299 = 4'h9 == _GEN_289[3:0] ? 1'h0 : _GEN_168; // @[Rob.scala 93:{25,25}]
  wire  _GEN_300 = 4'ha == _GEN_289[3:0] ? 1'h0 : _GEN_169; // @[Rob.scala 93:{25,25}]
  wire  _GEN_301 = 4'hb == _GEN_289[3:0] ? 1'h0 : _GEN_170; // @[Rob.scala 93:{25,25}]
  wire  _GEN_302 = 4'hc == _GEN_289[3:0] ? 1'h0 : _GEN_171; // @[Rob.scala 93:{25,25}]
  wire  _GEN_303 = 4'hd == _GEN_289[3:0] ? 1'h0 : _GEN_172; // @[Rob.scala 93:{25,25}]
  wire  _GEN_304 = 4'he == _GEN_289[3:0] ? 1'h0 : _GEN_173; // @[Rob.scala 93:{25,25}]
  wire  _GEN_305 = 4'hf == _GEN_289[3:0] ? 1'h0 : _GEN_174; // @[Rob.scala 93:{25,25}]
  wire  _GEN_322 = 4'h0 == _GEN_289[3:0] ? 1'h0 : _GEN_191; // @[Rob.scala 94:{20,20}]
  wire  _GEN_323 = 4'h1 == _GEN_289[3:0] ? 1'h0 : _GEN_192; // @[Rob.scala 94:{20,20}]
  wire  _GEN_324 = 4'h2 == _GEN_289[3:0] ? 1'h0 : _GEN_193; // @[Rob.scala 94:{20,20}]
  wire  _GEN_325 = 4'h3 == _GEN_289[3:0] ? 1'h0 : _GEN_194; // @[Rob.scala 94:{20,20}]
  wire  _GEN_326 = 4'h4 == _GEN_289[3:0] ? 1'h0 : _GEN_195; // @[Rob.scala 94:{20,20}]
  wire  _GEN_327 = 4'h5 == _GEN_289[3:0] ? 1'h0 : _GEN_196; // @[Rob.scala 94:{20,20}]
  wire  _GEN_328 = 4'h6 == _GEN_289[3:0] ? 1'h0 : _GEN_197; // @[Rob.scala 94:{20,20}]
  wire  _GEN_329 = 4'h7 == _GEN_289[3:0] ? 1'h0 : _GEN_198; // @[Rob.scala 94:{20,20}]
  wire  _GEN_330 = 4'h8 == _GEN_289[3:0] ? 1'h0 : _GEN_199; // @[Rob.scala 94:{20,20}]
  wire  _GEN_331 = 4'h9 == _GEN_289[3:0] ? 1'h0 : _GEN_200; // @[Rob.scala 94:{20,20}]
  wire  _GEN_332 = 4'ha == _GEN_289[3:0] ? 1'h0 : _GEN_201; // @[Rob.scala 94:{20,20}]
  wire  _GEN_333 = 4'hb == _GEN_289[3:0] ? 1'h0 : _GEN_202; // @[Rob.scala 94:{20,20}]
  wire  _GEN_334 = 4'hc == _GEN_289[3:0] ? 1'h0 : _GEN_203; // @[Rob.scala 94:{20,20}]
  wire  _GEN_335 = 4'hd == _GEN_289[3:0] ? 1'h0 : _GEN_204; // @[Rob.scala 94:{20,20}]
  wire  _GEN_336 = 4'he == _GEN_289[3:0] ? 1'h0 : _GEN_205; // @[Rob.scala 94:{20,20}]
  wire  _GEN_337 = 4'hf == _GEN_289[3:0] ? 1'h0 : _GEN_206; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_338 = 4'h0 == _GEN_289[3:0] ? 32'h0 : _GEN_207; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_339 = 4'h1 == _GEN_289[3:0] ? 32'h0 : _GEN_208; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_340 = 4'h2 == _GEN_289[3:0] ? 32'h0 : _GEN_209; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_341 = 4'h3 == _GEN_289[3:0] ? 32'h0 : _GEN_210; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_342 = 4'h4 == _GEN_289[3:0] ? 32'h0 : _GEN_211; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_343 = 4'h5 == _GEN_289[3:0] ? 32'h0 : _GEN_212; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_344 = 4'h6 == _GEN_289[3:0] ? 32'h0 : _GEN_213; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_345 = 4'h7 == _GEN_289[3:0] ? 32'h0 : _GEN_214; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_346 = 4'h8 == _GEN_289[3:0] ? 32'h0 : _GEN_215; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_347 = 4'h9 == _GEN_289[3:0] ? 32'h0 : _GEN_216; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_348 = 4'ha == _GEN_289[3:0] ? 32'h0 : _GEN_217; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_349 = 4'hb == _GEN_289[3:0] ? 32'h0 : _GEN_218; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_350 = 4'hc == _GEN_289[3:0] ? 32'h0 : _GEN_219; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_351 = 4'hd == _GEN_289[3:0] ? 32'h0 : _GEN_220; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_352 = 4'he == _GEN_289[3:0] ? 32'h0 : _GEN_221; // @[Rob.scala 94:{20,20}]
  wire [31:0] _GEN_353 = 4'hf == _GEN_289[3:0] ? 32'h0 : _GEN_222; // @[Rob.scala 94:{20,20}]
  wire  _GEN_354 = 4'h0 == _GEN_289[3:0] ? 1'h0 : _GEN_223; // @[Rob.scala 94:{20,20}]
  wire  _GEN_355 = 4'h1 == _GEN_289[3:0] ? 1'h0 : _GEN_224; // @[Rob.scala 94:{20,20}]
  wire  _GEN_356 = 4'h2 == _GEN_289[3:0] ? 1'h0 : _GEN_225; // @[Rob.scala 94:{20,20}]
  wire  _GEN_357 = 4'h3 == _GEN_289[3:0] ? 1'h0 : _GEN_226; // @[Rob.scala 94:{20,20}]
  wire  _GEN_358 = 4'h4 == _GEN_289[3:0] ? 1'h0 : _GEN_227; // @[Rob.scala 94:{20,20}]
  wire  _GEN_359 = 4'h5 == _GEN_289[3:0] ? 1'h0 : _GEN_228; // @[Rob.scala 94:{20,20}]
  wire  _GEN_360 = 4'h6 == _GEN_289[3:0] ? 1'h0 : _GEN_229; // @[Rob.scala 94:{20,20}]
  wire  _GEN_361 = 4'h7 == _GEN_289[3:0] ? 1'h0 : _GEN_230; // @[Rob.scala 94:{20,20}]
  wire  _GEN_362 = 4'h8 == _GEN_289[3:0] ? 1'h0 : _GEN_231; // @[Rob.scala 94:{20,20}]
  wire  _GEN_363 = 4'h9 == _GEN_289[3:0] ? 1'h0 : _GEN_232; // @[Rob.scala 94:{20,20}]
  wire  _GEN_364 = 4'ha == _GEN_289[3:0] ? 1'h0 : _GEN_233; // @[Rob.scala 94:{20,20}]
  wire  _GEN_365 = 4'hb == _GEN_289[3:0] ? 1'h0 : _GEN_234; // @[Rob.scala 94:{20,20}]
  wire  _GEN_366 = 4'hc == _GEN_289[3:0] ? 1'h0 : _GEN_235; // @[Rob.scala 94:{20,20}]
  wire  _GEN_367 = 4'hd == _GEN_289[3:0] ? 1'h0 : _GEN_236; // @[Rob.scala 94:{20,20}]
  wire  _GEN_368 = 4'he == _GEN_289[3:0] ? 1'h0 : _GEN_237; // @[Rob.scala 94:{20,20}]
  wire  _GEN_369 = 4'hf == _GEN_289[3:0] ? 1'h0 : _GEN_238; // @[Rob.scala 94:{20,20}]
  wire  _GEN_370 = 4'h0 == _GEN_289[3:0] ? 1'h0 : _GEN_239; // @[Rob.scala 94:{20,20}]
  wire  _GEN_371 = 4'h1 == _GEN_289[3:0] ? 1'h0 : _GEN_240; // @[Rob.scala 94:{20,20}]
  wire  _GEN_372 = 4'h2 == _GEN_289[3:0] ? 1'h0 : _GEN_241; // @[Rob.scala 94:{20,20}]
  wire  _GEN_373 = 4'h3 == _GEN_289[3:0] ? 1'h0 : _GEN_242; // @[Rob.scala 94:{20,20}]
  wire  _GEN_374 = 4'h4 == _GEN_289[3:0] ? 1'h0 : _GEN_243; // @[Rob.scala 94:{20,20}]
  wire  _GEN_375 = 4'h5 == _GEN_289[3:0] ? 1'h0 : _GEN_244; // @[Rob.scala 94:{20,20}]
  wire  _GEN_376 = 4'h6 == _GEN_289[3:0] ? 1'h0 : _GEN_245; // @[Rob.scala 94:{20,20}]
  wire  _GEN_377 = 4'h7 == _GEN_289[3:0] ? 1'h0 : _GEN_246; // @[Rob.scala 94:{20,20}]
  wire  _GEN_378 = 4'h8 == _GEN_289[3:0] ? 1'h0 : _GEN_247; // @[Rob.scala 94:{20,20}]
  wire  _GEN_379 = 4'h9 == _GEN_289[3:0] ? 1'h0 : _GEN_248; // @[Rob.scala 94:{20,20}]
  wire  _GEN_380 = 4'ha == _GEN_289[3:0] ? 1'h0 : _GEN_249; // @[Rob.scala 94:{20,20}]
  wire  _GEN_381 = 4'hb == _GEN_289[3:0] ? 1'h0 : _GEN_250; // @[Rob.scala 94:{20,20}]
  wire  _GEN_382 = 4'hc == _GEN_289[3:0] ? 1'h0 : _GEN_251; // @[Rob.scala 94:{20,20}]
  wire  _GEN_383 = 4'hd == _GEN_289[3:0] ? 1'h0 : _GEN_252; // @[Rob.scala 94:{20,20}]
  wire  _GEN_384 = 4'he == _GEN_289[3:0] ? 1'h0 : _GEN_253; // @[Rob.scala 94:{20,20}]
  wire  _GEN_385 = 4'hf == _GEN_289[3:0] ? 1'h0 : _GEN_254; // @[Rob.scala 94:{20,20}]
  wire  _GEN_402 = 4'h0 == _GEN_289[3:0] ? 1'h0 : _GEN_271; // @[Rob.scala 94:{20,20}]
  wire  _GEN_403 = 4'h1 == _GEN_289[3:0] ? 1'h0 : _GEN_272; // @[Rob.scala 94:{20,20}]
  wire  _GEN_404 = 4'h2 == _GEN_289[3:0] ? 1'h0 : _GEN_273; // @[Rob.scala 94:{20,20}]
  wire  _GEN_405 = 4'h3 == _GEN_289[3:0] ? 1'h0 : _GEN_274; // @[Rob.scala 94:{20,20}]
  wire  _GEN_406 = 4'h4 == _GEN_289[3:0] ? 1'h0 : _GEN_275; // @[Rob.scala 94:{20,20}]
  wire  _GEN_407 = 4'h5 == _GEN_289[3:0] ? 1'h0 : _GEN_276; // @[Rob.scala 94:{20,20}]
  wire  _GEN_408 = 4'h6 == _GEN_289[3:0] ? 1'h0 : _GEN_277; // @[Rob.scala 94:{20,20}]
  wire  _GEN_409 = 4'h7 == _GEN_289[3:0] ? 1'h0 : _GEN_278; // @[Rob.scala 94:{20,20}]
  wire  _GEN_410 = 4'h8 == _GEN_289[3:0] ? 1'h0 : _GEN_279; // @[Rob.scala 94:{20,20}]
  wire  _GEN_411 = 4'h9 == _GEN_289[3:0] ? 1'h0 : _GEN_280; // @[Rob.scala 94:{20,20}]
  wire  _GEN_412 = 4'ha == _GEN_289[3:0] ? 1'h0 : _GEN_281; // @[Rob.scala 94:{20,20}]
  wire  _GEN_413 = 4'hb == _GEN_289[3:0] ? 1'h0 : _GEN_282; // @[Rob.scala 94:{20,20}]
  wire  _GEN_414 = 4'hc == _GEN_289[3:0] ? 1'h0 : _GEN_283; // @[Rob.scala 94:{20,20}]
  wire  _GEN_415 = 4'hd == _GEN_289[3:0] ? 1'h0 : _GEN_284; // @[Rob.scala 94:{20,20}]
  wire  _GEN_416 = 4'he == _GEN_289[3:0] ? 1'h0 : _GEN_285; // @[Rob.scala 94:{20,20}]
  wire  _GEN_417 = 4'hf == _GEN_289[3:0] ? 1'h0 : _GEN_286; // @[Rob.scala 94:{20,20}]
  wire  _GEN_447 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_290 : _GEN_159; // @[Rob.scala 91:65]
  wire  _GEN_448 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_291 : _GEN_160; // @[Rob.scala 91:65]
  wire  _GEN_449 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_292 : _GEN_161; // @[Rob.scala 91:65]
  wire  _GEN_450 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_293 : _GEN_162; // @[Rob.scala 91:65]
  wire  _GEN_451 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_294 : _GEN_163; // @[Rob.scala 91:65]
  wire  _GEN_452 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_295 : _GEN_164; // @[Rob.scala 91:65]
  wire  _GEN_453 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_296 : _GEN_165; // @[Rob.scala 91:65]
  wire  _GEN_454 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_297 : _GEN_166; // @[Rob.scala 91:65]
  wire  _GEN_455 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_298 : _GEN_167; // @[Rob.scala 91:65]
  wire  _GEN_456 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_299 : _GEN_168; // @[Rob.scala 91:65]
  wire  _GEN_457 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_300 : _GEN_169; // @[Rob.scala 91:65]
  wire  _GEN_458 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_301 : _GEN_170; // @[Rob.scala 91:65]
  wire  _GEN_459 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_302 : _GEN_171; // @[Rob.scala 91:65]
  wire  _GEN_460 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_303 : _GEN_172; // @[Rob.scala 91:65]
  wire  _GEN_461 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_304 : _GEN_173; // @[Rob.scala 91:65]
  wire  _GEN_462 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_305 : _GEN_174; // @[Rob.scala 91:65]
  wire  _GEN_479 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_322 : _GEN_191; // @[Rob.scala 91:65]
  wire  _GEN_480 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_323 : _GEN_192; // @[Rob.scala 91:65]
  wire  _GEN_481 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_324 : _GEN_193; // @[Rob.scala 91:65]
  wire  _GEN_482 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_325 : _GEN_194; // @[Rob.scala 91:65]
  wire  _GEN_483 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_326 : _GEN_195; // @[Rob.scala 91:65]
  wire  _GEN_484 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_327 : _GEN_196; // @[Rob.scala 91:65]
  wire  _GEN_485 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_328 : _GEN_197; // @[Rob.scala 91:65]
  wire  _GEN_486 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_329 : _GEN_198; // @[Rob.scala 91:65]
  wire  _GEN_487 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_330 : _GEN_199; // @[Rob.scala 91:65]
  wire  _GEN_488 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_331 : _GEN_200; // @[Rob.scala 91:65]
  wire  _GEN_489 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_332 : _GEN_201; // @[Rob.scala 91:65]
  wire  _GEN_490 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_333 : _GEN_202; // @[Rob.scala 91:65]
  wire  _GEN_491 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_334 : _GEN_203; // @[Rob.scala 91:65]
  wire  _GEN_492 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_335 : _GEN_204; // @[Rob.scala 91:65]
  wire  _GEN_493 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_336 : _GEN_205; // @[Rob.scala 91:65]
  wire  _GEN_494 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_337 : _GEN_206; // @[Rob.scala 91:65]
  wire [31:0] _GEN_495 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_338 : _GEN_207; // @[Rob.scala 91:65]
  wire [31:0] _GEN_496 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_339 : _GEN_208; // @[Rob.scala 91:65]
  wire [31:0] _GEN_497 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_340 : _GEN_209; // @[Rob.scala 91:65]
  wire [31:0] _GEN_498 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_341 : _GEN_210; // @[Rob.scala 91:65]
  wire [31:0] _GEN_499 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_342 : _GEN_211; // @[Rob.scala 91:65]
  wire [31:0] _GEN_500 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_343 : _GEN_212; // @[Rob.scala 91:65]
  wire [31:0] _GEN_501 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_344 : _GEN_213; // @[Rob.scala 91:65]
  wire [31:0] _GEN_502 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_345 : _GEN_214; // @[Rob.scala 91:65]
  wire [31:0] _GEN_503 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_346 : _GEN_215; // @[Rob.scala 91:65]
  wire [31:0] _GEN_504 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_347 : _GEN_216; // @[Rob.scala 91:65]
  wire [31:0] _GEN_505 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_348 : _GEN_217; // @[Rob.scala 91:65]
  wire [31:0] _GEN_506 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_349 : _GEN_218; // @[Rob.scala 91:65]
  wire [31:0] _GEN_507 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_350 : _GEN_219; // @[Rob.scala 91:65]
  wire [31:0] _GEN_508 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_351 : _GEN_220; // @[Rob.scala 91:65]
  wire [31:0] _GEN_509 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_352 : _GEN_221; // @[Rob.scala 91:65]
  wire [31:0] _GEN_510 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_353 : _GEN_222; // @[Rob.scala 91:65]
  wire  _GEN_511 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_354 : _GEN_223; // @[Rob.scala 91:65]
  wire  _GEN_512 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_355 : _GEN_224; // @[Rob.scala 91:65]
  wire  _GEN_513 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_356 : _GEN_225; // @[Rob.scala 91:65]
  wire  _GEN_514 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_357 : _GEN_226; // @[Rob.scala 91:65]
  wire  _GEN_515 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_358 : _GEN_227; // @[Rob.scala 91:65]
  wire  _GEN_516 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_359 : _GEN_228; // @[Rob.scala 91:65]
  wire  _GEN_517 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_360 : _GEN_229; // @[Rob.scala 91:65]
  wire  _GEN_518 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_361 : _GEN_230; // @[Rob.scala 91:65]
  wire  _GEN_519 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_362 : _GEN_231; // @[Rob.scala 91:65]
  wire  _GEN_520 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_363 : _GEN_232; // @[Rob.scala 91:65]
  wire  _GEN_521 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_364 : _GEN_233; // @[Rob.scala 91:65]
  wire  _GEN_522 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_365 : _GEN_234; // @[Rob.scala 91:65]
  wire  _GEN_523 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_366 : _GEN_235; // @[Rob.scala 91:65]
  wire  _GEN_524 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_367 : _GEN_236; // @[Rob.scala 91:65]
  wire  _GEN_525 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_368 : _GEN_237; // @[Rob.scala 91:65]
  wire  _GEN_526 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_369 : _GEN_238; // @[Rob.scala 91:65]
  wire  _GEN_527 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_370 : _GEN_239; // @[Rob.scala 91:65]
  wire  _GEN_528 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_371 : _GEN_240; // @[Rob.scala 91:65]
  wire  _GEN_529 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_372 : _GEN_241; // @[Rob.scala 91:65]
  wire  _GEN_530 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_373 : _GEN_242; // @[Rob.scala 91:65]
  wire  _GEN_531 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_374 : _GEN_243; // @[Rob.scala 91:65]
  wire  _GEN_532 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_375 : _GEN_244; // @[Rob.scala 91:65]
  wire  _GEN_533 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_376 : _GEN_245; // @[Rob.scala 91:65]
  wire  _GEN_534 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_377 : _GEN_246; // @[Rob.scala 91:65]
  wire  _GEN_535 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_378 : _GEN_247; // @[Rob.scala 91:65]
  wire  _GEN_536 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_379 : _GEN_248; // @[Rob.scala 91:65]
  wire  _GEN_537 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_380 : _GEN_249; // @[Rob.scala 91:65]
  wire  _GEN_538 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_381 : _GEN_250; // @[Rob.scala 91:65]
  wire  _GEN_539 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_382 : _GEN_251; // @[Rob.scala 91:65]
  wire  _GEN_540 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_383 : _GEN_252; // @[Rob.scala 91:65]
  wire  _GEN_541 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_384 : _GEN_253; // @[Rob.scala 91:65]
  wire  _GEN_542 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_385 : _GEN_254; // @[Rob.scala 91:65]
  wire  _GEN_559 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_402 : _GEN_271; // @[Rob.scala 91:65]
  wire  _GEN_560 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_403 : _GEN_272; // @[Rob.scala 91:65]
  wire  _GEN_561 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_404 : _GEN_273; // @[Rob.scala 91:65]
  wire  _GEN_562 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_405 : _GEN_274; // @[Rob.scala 91:65]
  wire  _GEN_563 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_406 : _GEN_275; // @[Rob.scala 91:65]
  wire  _GEN_564 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_407 : _GEN_276; // @[Rob.scala 91:65]
  wire  _GEN_565 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_408 : _GEN_277; // @[Rob.scala 91:65]
  wire  _GEN_566 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_409 : _GEN_278; // @[Rob.scala 91:65]
  wire  _GEN_567 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_410 : _GEN_279; // @[Rob.scala 91:65]
  wire  _GEN_568 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_411 : _GEN_280; // @[Rob.scala 91:65]
  wire  _GEN_569 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_412 : _GEN_281; // @[Rob.scala 91:65]
  wire  _GEN_570 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_413 : _GEN_282; // @[Rob.scala 91:65]
  wire  _GEN_571 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_414 : _GEN_283; // @[Rob.scala 91:65]
  wire  _GEN_572 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_415 : _GEN_284; // @[Rob.scala 91:65]
  wire  _GEN_573 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_416 : _GEN_285; // @[Rob.scala 91:65]
  wire  _GEN_574 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_417 : _GEN_286; // @[Rob.scala 91:65]
  wire [4:0] next_enq_vec_0 = enq_vec_0 + _GEN_2224; // @[Rob.scala 101:44]
  wire [4:0] next_enq_vec_1 = enq_vec_1 + _GEN_2224; // @[Rob.scala 101:44]
  wire  _GEN_578 = 4'h0 == io_exe_0_rob_addr | _GEN_447; // @[Rob.scala 114:{26,26}]
  wire  _GEN_579 = 4'h1 == io_exe_0_rob_addr | _GEN_448; // @[Rob.scala 114:{26,26}]
  wire  _GEN_580 = 4'h2 == io_exe_0_rob_addr | _GEN_449; // @[Rob.scala 114:{26,26}]
  wire  _GEN_581 = 4'h3 == io_exe_0_rob_addr | _GEN_450; // @[Rob.scala 114:{26,26}]
  wire  _GEN_582 = 4'h4 == io_exe_0_rob_addr | _GEN_451; // @[Rob.scala 114:{26,26}]
  wire  _GEN_583 = 4'h5 == io_exe_0_rob_addr | _GEN_452; // @[Rob.scala 114:{26,26}]
  wire  _GEN_584 = 4'h6 == io_exe_0_rob_addr | _GEN_453; // @[Rob.scala 114:{26,26}]
  wire  _GEN_585 = 4'h7 == io_exe_0_rob_addr | _GEN_454; // @[Rob.scala 114:{26,26}]
  wire  _GEN_586 = 4'h8 == io_exe_0_rob_addr | _GEN_455; // @[Rob.scala 114:{26,26}]
  wire  _GEN_587 = 4'h9 == io_exe_0_rob_addr | _GEN_456; // @[Rob.scala 114:{26,26}]
  wire  _GEN_588 = 4'ha == io_exe_0_rob_addr | _GEN_457; // @[Rob.scala 114:{26,26}]
  wire  _GEN_589 = 4'hb == io_exe_0_rob_addr | _GEN_458; // @[Rob.scala 114:{26,26}]
  wire  _GEN_590 = 4'hc == io_exe_0_rob_addr | _GEN_459; // @[Rob.scala 114:{26,26}]
  wire  _GEN_591 = 4'hd == io_exe_0_rob_addr | _GEN_460; // @[Rob.scala 114:{26,26}]
  wire  _GEN_592 = 4'he == io_exe_0_rob_addr | _GEN_461; // @[Rob.scala 114:{26,26}]
  wire  _GEN_593 = 4'hf == io_exe_0_rob_addr | _GEN_462; // @[Rob.scala 114:{26,26}]
  wire  _GEN_610 = 4'h0 == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_479; // @[Rob.scala 115:{21,21}]
  wire  _GEN_611 = 4'h1 == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_480; // @[Rob.scala 115:{21,21}]
  wire  _GEN_612 = 4'h2 == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_481; // @[Rob.scala 115:{21,21}]
  wire  _GEN_613 = 4'h3 == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_482; // @[Rob.scala 115:{21,21}]
  wire  _GEN_614 = 4'h4 == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_483; // @[Rob.scala 115:{21,21}]
  wire  _GEN_615 = 4'h5 == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_484; // @[Rob.scala 115:{21,21}]
  wire  _GEN_616 = 4'h6 == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_485; // @[Rob.scala 115:{21,21}]
  wire  _GEN_617 = 4'h7 == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_486; // @[Rob.scala 115:{21,21}]
  wire  _GEN_618 = 4'h8 == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_487; // @[Rob.scala 115:{21,21}]
  wire  _GEN_619 = 4'h9 == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_488; // @[Rob.scala 115:{21,21}]
  wire  _GEN_620 = 4'ha == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_489; // @[Rob.scala 115:{21,21}]
  wire  _GEN_621 = 4'hb == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_490; // @[Rob.scala 115:{21,21}]
  wire  _GEN_622 = 4'hc == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_491; // @[Rob.scala 115:{21,21}]
  wire  _GEN_623 = 4'hd == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_492; // @[Rob.scala 115:{21,21}]
  wire  _GEN_624 = 4'he == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_493; // @[Rob.scala 115:{21,21}]
  wire  _GEN_625 = 4'hf == io_exe_0_rob_addr ? io_exe_ecp_0_mis : _GEN_494; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_626 = 4'h0 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_495; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_627 = 4'h1 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_496; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_628 = 4'h2 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_497; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_629 = 4'h3 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_498; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_630 = 4'h4 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_499; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_631 = 4'h5 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_500; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_632 = 4'h6 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_501; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_633 = 4'h7 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_502; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_634 = 4'h8 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_503; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_635 = 4'h9 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_504; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_636 = 4'ha == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_505; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_637 = 4'hb == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_506; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_638 = 4'hc == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_507; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_639 = 4'hd == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_508; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_640 = 4'he == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_509; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_641 = 4'hf == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_pc : _GEN_510; // @[Rob.scala 115:{21,21}]
  wire  _GEN_642 = 4'h0 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_511; // @[Rob.scala 115:{21,21}]
  wire  _GEN_643 = 4'h1 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_512; // @[Rob.scala 115:{21,21}]
  wire  _GEN_644 = 4'h2 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_513; // @[Rob.scala 115:{21,21}]
  wire  _GEN_645 = 4'h3 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_514; // @[Rob.scala 115:{21,21}]
  wire  _GEN_646 = 4'h4 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_515; // @[Rob.scala 115:{21,21}]
  wire  _GEN_647 = 4'h5 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_516; // @[Rob.scala 115:{21,21}]
  wire  _GEN_648 = 4'h6 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_517; // @[Rob.scala 115:{21,21}]
  wire  _GEN_649 = 4'h7 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_518; // @[Rob.scala 115:{21,21}]
  wire  _GEN_650 = 4'h8 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_519; // @[Rob.scala 115:{21,21}]
  wire  _GEN_651 = 4'h9 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_520; // @[Rob.scala 115:{21,21}]
  wire  _GEN_652 = 4'ha == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_521; // @[Rob.scala 115:{21,21}]
  wire  _GEN_653 = 4'hb == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_522; // @[Rob.scala 115:{21,21}]
  wire  _GEN_654 = 4'hc == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_523; // @[Rob.scala 115:{21,21}]
  wire  _GEN_655 = 4'hd == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_524; // @[Rob.scala 115:{21,21}]
  wire  _GEN_656 = 4'he == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_525; // @[Rob.scala 115:{21,21}]
  wire  _GEN_657 = 4'hf == io_exe_0_rob_addr ? io_exe_ecp_0_jmp : _GEN_526; // @[Rob.scala 115:{21,21}]
  wire  _GEN_658 = 4'h0 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_527; // @[Rob.scala 115:{21,21}]
  wire  _GEN_659 = 4'h1 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_528; // @[Rob.scala 115:{21,21}]
  wire  _GEN_660 = 4'h2 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_529; // @[Rob.scala 115:{21,21}]
  wire  _GEN_661 = 4'h3 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_530; // @[Rob.scala 115:{21,21}]
  wire  _GEN_662 = 4'h4 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_531; // @[Rob.scala 115:{21,21}]
  wire  _GEN_663 = 4'h5 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_532; // @[Rob.scala 115:{21,21}]
  wire  _GEN_664 = 4'h6 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_533; // @[Rob.scala 115:{21,21}]
  wire  _GEN_665 = 4'h7 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_534; // @[Rob.scala 115:{21,21}]
  wire  _GEN_666 = 4'h8 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_535; // @[Rob.scala 115:{21,21}]
  wire  _GEN_667 = 4'h9 == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_536; // @[Rob.scala 115:{21,21}]
  wire  _GEN_668 = 4'ha == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_537; // @[Rob.scala 115:{21,21}]
  wire  _GEN_669 = 4'hb == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_538; // @[Rob.scala 115:{21,21}]
  wire  _GEN_670 = 4'hc == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_539; // @[Rob.scala 115:{21,21}]
  wire  _GEN_671 = 4'hd == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_540; // @[Rob.scala 115:{21,21}]
  wire  _GEN_672 = 4'he == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_541; // @[Rob.scala 115:{21,21}]
  wire  _GEN_673 = 4'hf == io_exe_0_rob_addr ? io_exe_ecp_0_jmp_valid : _GEN_542; // @[Rob.scala 115:{21,21}]
  wire  _GEN_690 = 4'h0 == io_exe_0_rob_addr ? 1'h0 : _GEN_559; // @[Rob.scala 115:{21,21}]
  wire  _GEN_691 = 4'h1 == io_exe_0_rob_addr ? 1'h0 : _GEN_560; // @[Rob.scala 115:{21,21}]
  wire  _GEN_692 = 4'h2 == io_exe_0_rob_addr ? 1'h0 : _GEN_561; // @[Rob.scala 115:{21,21}]
  wire  _GEN_693 = 4'h3 == io_exe_0_rob_addr ? 1'h0 : _GEN_562; // @[Rob.scala 115:{21,21}]
  wire  _GEN_694 = 4'h4 == io_exe_0_rob_addr ? 1'h0 : _GEN_563; // @[Rob.scala 115:{21,21}]
  wire  _GEN_695 = 4'h5 == io_exe_0_rob_addr ? 1'h0 : _GEN_564; // @[Rob.scala 115:{21,21}]
  wire  _GEN_696 = 4'h6 == io_exe_0_rob_addr ? 1'h0 : _GEN_565; // @[Rob.scala 115:{21,21}]
  wire  _GEN_697 = 4'h7 == io_exe_0_rob_addr ? 1'h0 : _GEN_566; // @[Rob.scala 115:{21,21}]
  wire  _GEN_698 = 4'h8 == io_exe_0_rob_addr ? 1'h0 : _GEN_567; // @[Rob.scala 115:{21,21}]
  wire  _GEN_699 = 4'h9 == io_exe_0_rob_addr ? 1'h0 : _GEN_568; // @[Rob.scala 115:{21,21}]
  wire  _GEN_700 = 4'ha == io_exe_0_rob_addr ? 1'h0 : _GEN_569; // @[Rob.scala 115:{21,21}]
  wire  _GEN_701 = 4'hb == io_exe_0_rob_addr ? 1'h0 : _GEN_570; // @[Rob.scala 115:{21,21}]
  wire  _GEN_702 = 4'hc == io_exe_0_rob_addr ? 1'h0 : _GEN_571; // @[Rob.scala 115:{21,21}]
  wire  _GEN_703 = 4'hd == io_exe_0_rob_addr ? 1'h0 : _GEN_572; // @[Rob.scala 115:{21,21}]
  wire  _GEN_704 = 4'he == io_exe_0_rob_addr ? 1'h0 : _GEN_573; // @[Rob.scala 115:{21,21}]
  wire  _GEN_705 = 4'hf == io_exe_0_rob_addr ? 1'h0 : _GEN_574; // @[Rob.scala 115:{21,21}]
  wire  _GEN_706 = io_exe_0_valid ? _GEN_578 : _GEN_447; // @[Rob.scala 113:28]
  wire  _GEN_707 = io_exe_0_valid ? _GEN_579 : _GEN_448; // @[Rob.scala 113:28]
  wire  _GEN_708 = io_exe_0_valid ? _GEN_580 : _GEN_449; // @[Rob.scala 113:28]
  wire  _GEN_709 = io_exe_0_valid ? _GEN_581 : _GEN_450; // @[Rob.scala 113:28]
  wire  _GEN_710 = io_exe_0_valid ? _GEN_582 : _GEN_451; // @[Rob.scala 113:28]
  wire  _GEN_711 = io_exe_0_valid ? _GEN_583 : _GEN_452; // @[Rob.scala 113:28]
  wire  _GEN_712 = io_exe_0_valid ? _GEN_584 : _GEN_453; // @[Rob.scala 113:28]
  wire  _GEN_713 = io_exe_0_valid ? _GEN_585 : _GEN_454; // @[Rob.scala 113:28]
  wire  _GEN_714 = io_exe_0_valid ? _GEN_586 : _GEN_455; // @[Rob.scala 113:28]
  wire  _GEN_715 = io_exe_0_valid ? _GEN_587 : _GEN_456; // @[Rob.scala 113:28]
  wire  _GEN_716 = io_exe_0_valid ? _GEN_588 : _GEN_457; // @[Rob.scala 113:28]
  wire  _GEN_717 = io_exe_0_valid ? _GEN_589 : _GEN_458; // @[Rob.scala 113:28]
  wire  _GEN_718 = io_exe_0_valid ? _GEN_590 : _GEN_459; // @[Rob.scala 113:28]
  wire  _GEN_719 = io_exe_0_valid ? _GEN_591 : _GEN_460; // @[Rob.scala 113:28]
  wire  _GEN_720 = io_exe_0_valid ? _GEN_592 : _GEN_461; // @[Rob.scala 113:28]
  wire  _GEN_721 = io_exe_0_valid ? _GEN_593 : _GEN_462; // @[Rob.scala 113:28]
  wire  _GEN_738 = io_exe_0_valid ? _GEN_610 : _GEN_479; // @[Rob.scala 113:28]
  wire  _GEN_739 = io_exe_0_valid ? _GEN_611 : _GEN_480; // @[Rob.scala 113:28]
  wire  _GEN_740 = io_exe_0_valid ? _GEN_612 : _GEN_481; // @[Rob.scala 113:28]
  wire  _GEN_741 = io_exe_0_valid ? _GEN_613 : _GEN_482; // @[Rob.scala 113:28]
  wire  _GEN_742 = io_exe_0_valid ? _GEN_614 : _GEN_483; // @[Rob.scala 113:28]
  wire  _GEN_743 = io_exe_0_valid ? _GEN_615 : _GEN_484; // @[Rob.scala 113:28]
  wire  _GEN_744 = io_exe_0_valid ? _GEN_616 : _GEN_485; // @[Rob.scala 113:28]
  wire  _GEN_745 = io_exe_0_valid ? _GEN_617 : _GEN_486; // @[Rob.scala 113:28]
  wire  _GEN_746 = io_exe_0_valid ? _GEN_618 : _GEN_487; // @[Rob.scala 113:28]
  wire  _GEN_747 = io_exe_0_valid ? _GEN_619 : _GEN_488; // @[Rob.scala 113:28]
  wire  _GEN_748 = io_exe_0_valid ? _GEN_620 : _GEN_489; // @[Rob.scala 113:28]
  wire  _GEN_749 = io_exe_0_valid ? _GEN_621 : _GEN_490; // @[Rob.scala 113:28]
  wire  _GEN_750 = io_exe_0_valid ? _GEN_622 : _GEN_491; // @[Rob.scala 113:28]
  wire  _GEN_751 = io_exe_0_valid ? _GEN_623 : _GEN_492; // @[Rob.scala 113:28]
  wire  _GEN_752 = io_exe_0_valid ? _GEN_624 : _GEN_493; // @[Rob.scala 113:28]
  wire  _GEN_753 = io_exe_0_valid ? _GEN_625 : _GEN_494; // @[Rob.scala 113:28]
  wire [31:0] _GEN_754 = io_exe_0_valid ? _GEN_626 : _GEN_495; // @[Rob.scala 113:28]
  wire [31:0] _GEN_755 = io_exe_0_valid ? _GEN_627 : _GEN_496; // @[Rob.scala 113:28]
  wire [31:0] _GEN_756 = io_exe_0_valid ? _GEN_628 : _GEN_497; // @[Rob.scala 113:28]
  wire [31:0] _GEN_757 = io_exe_0_valid ? _GEN_629 : _GEN_498; // @[Rob.scala 113:28]
  wire [31:0] _GEN_758 = io_exe_0_valid ? _GEN_630 : _GEN_499; // @[Rob.scala 113:28]
  wire [31:0] _GEN_759 = io_exe_0_valid ? _GEN_631 : _GEN_500; // @[Rob.scala 113:28]
  wire [31:0] _GEN_760 = io_exe_0_valid ? _GEN_632 : _GEN_501; // @[Rob.scala 113:28]
  wire [31:0] _GEN_761 = io_exe_0_valid ? _GEN_633 : _GEN_502; // @[Rob.scala 113:28]
  wire [31:0] _GEN_762 = io_exe_0_valid ? _GEN_634 : _GEN_503; // @[Rob.scala 113:28]
  wire [31:0] _GEN_763 = io_exe_0_valid ? _GEN_635 : _GEN_504; // @[Rob.scala 113:28]
  wire [31:0] _GEN_764 = io_exe_0_valid ? _GEN_636 : _GEN_505; // @[Rob.scala 113:28]
  wire [31:0] _GEN_765 = io_exe_0_valid ? _GEN_637 : _GEN_506; // @[Rob.scala 113:28]
  wire [31:0] _GEN_766 = io_exe_0_valid ? _GEN_638 : _GEN_507; // @[Rob.scala 113:28]
  wire [31:0] _GEN_767 = io_exe_0_valid ? _GEN_639 : _GEN_508; // @[Rob.scala 113:28]
  wire [31:0] _GEN_768 = io_exe_0_valid ? _GEN_640 : _GEN_509; // @[Rob.scala 113:28]
  wire [31:0] _GEN_769 = io_exe_0_valid ? _GEN_641 : _GEN_510; // @[Rob.scala 113:28]
  wire  _GEN_770 = io_exe_0_valid ? _GEN_642 : _GEN_511; // @[Rob.scala 113:28]
  wire  _GEN_771 = io_exe_0_valid ? _GEN_643 : _GEN_512; // @[Rob.scala 113:28]
  wire  _GEN_772 = io_exe_0_valid ? _GEN_644 : _GEN_513; // @[Rob.scala 113:28]
  wire  _GEN_773 = io_exe_0_valid ? _GEN_645 : _GEN_514; // @[Rob.scala 113:28]
  wire  _GEN_774 = io_exe_0_valid ? _GEN_646 : _GEN_515; // @[Rob.scala 113:28]
  wire  _GEN_775 = io_exe_0_valid ? _GEN_647 : _GEN_516; // @[Rob.scala 113:28]
  wire  _GEN_776 = io_exe_0_valid ? _GEN_648 : _GEN_517; // @[Rob.scala 113:28]
  wire  _GEN_777 = io_exe_0_valid ? _GEN_649 : _GEN_518; // @[Rob.scala 113:28]
  wire  _GEN_778 = io_exe_0_valid ? _GEN_650 : _GEN_519; // @[Rob.scala 113:28]
  wire  _GEN_779 = io_exe_0_valid ? _GEN_651 : _GEN_520; // @[Rob.scala 113:28]
  wire  _GEN_780 = io_exe_0_valid ? _GEN_652 : _GEN_521; // @[Rob.scala 113:28]
  wire  _GEN_781 = io_exe_0_valid ? _GEN_653 : _GEN_522; // @[Rob.scala 113:28]
  wire  _GEN_782 = io_exe_0_valid ? _GEN_654 : _GEN_523; // @[Rob.scala 113:28]
  wire  _GEN_783 = io_exe_0_valid ? _GEN_655 : _GEN_524; // @[Rob.scala 113:28]
  wire  _GEN_784 = io_exe_0_valid ? _GEN_656 : _GEN_525; // @[Rob.scala 113:28]
  wire  _GEN_785 = io_exe_0_valid ? _GEN_657 : _GEN_526; // @[Rob.scala 113:28]
  wire  _GEN_786 = io_exe_0_valid ? _GEN_658 : _GEN_527; // @[Rob.scala 113:28]
  wire  _GEN_787 = io_exe_0_valid ? _GEN_659 : _GEN_528; // @[Rob.scala 113:28]
  wire  _GEN_788 = io_exe_0_valid ? _GEN_660 : _GEN_529; // @[Rob.scala 113:28]
  wire  _GEN_789 = io_exe_0_valid ? _GEN_661 : _GEN_530; // @[Rob.scala 113:28]
  wire  _GEN_790 = io_exe_0_valid ? _GEN_662 : _GEN_531; // @[Rob.scala 113:28]
  wire  _GEN_791 = io_exe_0_valid ? _GEN_663 : _GEN_532; // @[Rob.scala 113:28]
  wire  _GEN_792 = io_exe_0_valid ? _GEN_664 : _GEN_533; // @[Rob.scala 113:28]
  wire  _GEN_793 = io_exe_0_valid ? _GEN_665 : _GEN_534; // @[Rob.scala 113:28]
  wire  _GEN_794 = io_exe_0_valid ? _GEN_666 : _GEN_535; // @[Rob.scala 113:28]
  wire  _GEN_795 = io_exe_0_valid ? _GEN_667 : _GEN_536; // @[Rob.scala 113:28]
  wire  _GEN_796 = io_exe_0_valid ? _GEN_668 : _GEN_537; // @[Rob.scala 113:28]
  wire  _GEN_797 = io_exe_0_valid ? _GEN_669 : _GEN_538; // @[Rob.scala 113:28]
  wire  _GEN_798 = io_exe_0_valid ? _GEN_670 : _GEN_539; // @[Rob.scala 113:28]
  wire  _GEN_799 = io_exe_0_valid ? _GEN_671 : _GEN_540; // @[Rob.scala 113:28]
  wire  _GEN_800 = io_exe_0_valid ? _GEN_672 : _GEN_541; // @[Rob.scala 113:28]
  wire  _GEN_801 = io_exe_0_valid ? _GEN_673 : _GEN_542; // @[Rob.scala 113:28]
  wire  _GEN_818 = io_exe_0_valid ? _GEN_690 : _GEN_559; // @[Rob.scala 113:28]
  wire  _GEN_819 = io_exe_0_valid ? _GEN_691 : _GEN_560; // @[Rob.scala 113:28]
  wire  _GEN_820 = io_exe_0_valid ? _GEN_692 : _GEN_561; // @[Rob.scala 113:28]
  wire  _GEN_821 = io_exe_0_valid ? _GEN_693 : _GEN_562; // @[Rob.scala 113:28]
  wire  _GEN_822 = io_exe_0_valid ? _GEN_694 : _GEN_563; // @[Rob.scala 113:28]
  wire  _GEN_823 = io_exe_0_valid ? _GEN_695 : _GEN_564; // @[Rob.scala 113:28]
  wire  _GEN_824 = io_exe_0_valid ? _GEN_696 : _GEN_565; // @[Rob.scala 113:28]
  wire  _GEN_825 = io_exe_0_valid ? _GEN_697 : _GEN_566; // @[Rob.scala 113:28]
  wire  _GEN_826 = io_exe_0_valid ? _GEN_698 : _GEN_567; // @[Rob.scala 113:28]
  wire  _GEN_827 = io_exe_0_valid ? _GEN_699 : _GEN_568; // @[Rob.scala 113:28]
  wire  _GEN_828 = io_exe_0_valid ? _GEN_700 : _GEN_569; // @[Rob.scala 113:28]
  wire  _GEN_829 = io_exe_0_valid ? _GEN_701 : _GEN_570; // @[Rob.scala 113:28]
  wire  _GEN_830 = io_exe_0_valid ? _GEN_702 : _GEN_571; // @[Rob.scala 113:28]
  wire  _GEN_831 = io_exe_0_valid ? _GEN_703 : _GEN_572; // @[Rob.scala 113:28]
  wire  _GEN_832 = io_exe_0_valid ? _GEN_704 : _GEN_573; // @[Rob.scala 113:28]
  wire  _GEN_833 = io_exe_0_valid ? _GEN_705 : _GEN_574; // @[Rob.scala 113:28]
  wire  _GEN_834 = 4'h0 == io_exe_1_rob_addr | _GEN_706; // @[Rob.scala 114:{26,26}]
  wire  _GEN_835 = 4'h1 == io_exe_1_rob_addr | _GEN_707; // @[Rob.scala 114:{26,26}]
  wire  _GEN_836 = 4'h2 == io_exe_1_rob_addr | _GEN_708; // @[Rob.scala 114:{26,26}]
  wire  _GEN_837 = 4'h3 == io_exe_1_rob_addr | _GEN_709; // @[Rob.scala 114:{26,26}]
  wire  _GEN_838 = 4'h4 == io_exe_1_rob_addr | _GEN_710; // @[Rob.scala 114:{26,26}]
  wire  _GEN_839 = 4'h5 == io_exe_1_rob_addr | _GEN_711; // @[Rob.scala 114:{26,26}]
  wire  _GEN_840 = 4'h6 == io_exe_1_rob_addr | _GEN_712; // @[Rob.scala 114:{26,26}]
  wire  _GEN_841 = 4'h7 == io_exe_1_rob_addr | _GEN_713; // @[Rob.scala 114:{26,26}]
  wire  _GEN_842 = 4'h8 == io_exe_1_rob_addr | _GEN_714; // @[Rob.scala 114:{26,26}]
  wire  _GEN_843 = 4'h9 == io_exe_1_rob_addr | _GEN_715; // @[Rob.scala 114:{26,26}]
  wire  _GEN_844 = 4'ha == io_exe_1_rob_addr | _GEN_716; // @[Rob.scala 114:{26,26}]
  wire  _GEN_845 = 4'hb == io_exe_1_rob_addr | _GEN_717; // @[Rob.scala 114:{26,26}]
  wire  _GEN_846 = 4'hc == io_exe_1_rob_addr | _GEN_718; // @[Rob.scala 114:{26,26}]
  wire  _GEN_847 = 4'hd == io_exe_1_rob_addr | _GEN_719; // @[Rob.scala 114:{26,26}]
  wire  _GEN_848 = 4'he == io_exe_1_rob_addr | _GEN_720; // @[Rob.scala 114:{26,26}]
  wire  _GEN_849 = 4'hf == io_exe_1_rob_addr | _GEN_721; // @[Rob.scala 114:{26,26}]
  wire  _GEN_866 = 4'h0 == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_738; // @[Rob.scala 115:{21,21}]
  wire  _GEN_867 = 4'h1 == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_739; // @[Rob.scala 115:{21,21}]
  wire  _GEN_868 = 4'h2 == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_740; // @[Rob.scala 115:{21,21}]
  wire  _GEN_869 = 4'h3 == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_741; // @[Rob.scala 115:{21,21}]
  wire  _GEN_870 = 4'h4 == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_742; // @[Rob.scala 115:{21,21}]
  wire  _GEN_871 = 4'h5 == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_743; // @[Rob.scala 115:{21,21}]
  wire  _GEN_872 = 4'h6 == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_744; // @[Rob.scala 115:{21,21}]
  wire  _GEN_873 = 4'h7 == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_745; // @[Rob.scala 115:{21,21}]
  wire  _GEN_874 = 4'h8 == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_746; // @[Rob.scala 115:{21,21}]
  wire  _GEN_875 = 4'h9 == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_747; // @[Rob.scala 115:{21,21}]
  wire  _GEN_876 = 4'ha == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_748; // @[Rob.scala 115:{21,21}]
  wire  _GEN_877 = 4'hb == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_749; // @[Rob.scala 115:{21,21}]
  wire  _GEN_878 = 4'hc == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_750; // @[Rob.scala 115:{21,21}]
  wire  _GEN_879 = 4'hd == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_751; // @[Rob.scala 115:{21,21}]
  wire  _GEN_880 = 4'he == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_752; // @[Rob.scala 115:{21,21}]
  wire  _GEN_881 = 4'hf == io_exe_1_rob_addr ? io_exe_ecp_1_mis : _GEN_753; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_882 = 4'h0 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_754; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_883 = 4'h1 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_755; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_884 = 4'h2 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_756; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_885 = 4'h3 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_757; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_886 = 4'h4 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_758; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_887 = 4'h5 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_759; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_888 = 4'h6 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_760; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_889 = 4'h7 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_761; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_890 = 4'h8 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_762; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_891 = 4'h9 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_763; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_892 = 4'ha == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_764; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_893 = 4'hb == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_765; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_894 = 4'hc == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_766; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_895 = 4'hd == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_767; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_896 = 4'he == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_768; // @[Rob.scala 115:{21,21}]
  wire [31:0] _GEN_897 = 4'hf == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_pc : _GEN_769; // @[Rob.scala 115:{21,21}]
  wire  _GEN_898 = 4'h0 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_770; // @[Rob.scala 115:{21,21}]
  wire  _GEN_899 = 4'h1 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_771; // @[Rob.scala 115:{21,21}]
  wire  _GEN_900 = 4'h2 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_772; // @[Rob.scala 115:{21,21}]
  wire  _GEN_901 = 4'h3 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_773; // @[Rob.scala 115:{21,21}]
  wire  _GEN_902 = 4'h4 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_774; // @[Rob.scala 115:{21,21}]
  wire  _GEN_903 = 4'h5 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_775; // @[Rob.scala 115:{21,21}]
  wire  _GEN_904 = 4'h6 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_776; // @[Rob.scala 115:{21,21}]
  wire  _GEN_905 = 4'h7 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_777; // @[Rob.scala 115:{21,21}]
  wire  _GEN_906 = 4'h8 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_778; // @[Rob.scala 115:{21,21}]
  wire  _GEN_907 = 4'h9 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_779; // @[Rob.scala 115:{21,21}]
  wire  _GEN_908 = 4'ha == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_780; // @[Rob.scala 115:{21,21}]
  wire  _GEN_909 = 4'hb == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_781; // @[Rob.scala 115:{21,21}]
  wire  _GEN_910 = 4'hc == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_782; // @[Rob.scala 115:{21,21}]
  wire  _GEN_911 = 4'hd == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_783; // @[Rob.scala 115:{21,21}]
  wire  _GEN_912 = 4'he == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_784; // @[Rob.scala 115:{21,21}]
  wire  _GEN_913 = 4'hf == io_exe_1_rob_addr ? io_exe_ecp_1_jmp : _GEN_785; // @[Rob.scala 115:{21,21}]
  wire  _GEN_914 = 4'h0 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_786; // @[Rob.scala 115:{21,21}]
  wire  _GEN_915 = 4'h1 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_787; // @[Rob.scala 115:{21,21}]
  wire  _GEN_916 = 4'h2 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_788; // @[Rob.scala 115:{21,21}]
  wire  _GEN_917 = 4'h3 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_789; // @[Rob.scala 115:{21,21}]
  wire  _GEN_918 = 4'h4 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_790; // @[Rob.scala 115:{21,21}]
  wire  _GEN_919 = 4'h5 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_791; // @[Rob.scala 115:{21,21}]
  wire  _GEN_920 = 4'h6 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_792; // @[Rob.scala 115:{21,21}]
  wire  _GEN_921 = 4'h7 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_793; // @[Rob.scala 115:{21,21}]
  wire  _GEN_922 = 4'h8 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_794; // @[Rob.scala 115:{21,21}]
  wire  _GEN_923 = 4'h9 == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_795; // @[Rob.scala 115:{21,21}]
  wire  _GEN_924 = 4'ha == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_796; // @[Rob.scala 115:{21,21}]
  wire  _GEN_925 = 4'hb == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_797; // @[Rob.scala 115:{21,21}]
  wire  _GEN_926 = 4'hc == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_798; // @[Rob.scala 115:{21,21}]
  wire  _GEN_927 = 4'hd == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_799; // @[Rob.scala 115:{21,21}]
  wire  _GEN_928 = 4'he == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_800; // @[Rob.scala 115:{21,21}]
  wire  _GEN_929 = 4'hf == io_exe_1_rob_addr ? io_exe_ecp_1_jmp_valid : _GEN_801; // @[Rob.scala 115:{21,21}]
  wire  _GEN_946 = 4'h0 == io_exe_1_rob_addr ? 1'h0 : _GEN_818; // @[Rob.scala 115:{21,21}]
  wire  _GEN_947 = 4'h1 == io_exe_1_rob_addr ? 1'h0 : _GEN_819; // @[Rob.scala 115:{21,21}]
  wire  _GEN_948 = 4'h2 == io_exe_1_rob_addr ? 1'h0 : _GEN_820; // @[Rob.scala 115:{21,21}]
  wire  _GEN_949 = 4'h3 == io_exe_1_rob_addr ? 1'h0 : _GEN_821; // @[Rob.scala 115:{21,21}]
  wire  _GEN_950 = 4'h4 == io_exe_1_rob_addr ? 1'h0 : _GEN_822; // @[Rob.scala 115:{21,21}]
  wire  _GEN_951 = 4'h5 == io_exe_1_rob_addr ? 1'h0 : _GEN_823; // @[Rob.scala 115:{21,21}]
  wire  _GEN_952 = 4'h6 == io_exe_1_rob_addr ? 1'h0 : _GEN_824; // @[Rob.scala 115:{21,21}]
  wire  _GEN_953 = 4'h7 == io_exe_1_rob_addr ? 1'h0 : _GEN_825; // @[Rob.scala 115:{21,21}]
  wire  _GEN_954 = 4'h8 == io_exe_1_rob_addr ? 1'h0 : _GEN_826; // @[Rob.scala 115:{21,21}]
  wire  _GEN_955 = 4'h9 == io_exe_1_rob_addr ? 1'h0 : _GEN_827; // @[Rob.scala 115:{21,21}]
  wire  _GEN_956 = 4'ha == io_exe_1_rob_addr ? 1'h0 : _GEN_828; // @[Rob.scala 115:{21,21}]
  wire  _GEN_957 = 4'hb == io_exe_1_rob_addr ? 1'h0 : _GEN_829; // @[Rob.scala 115:{21,21}]
  wire  _GEN_958 = 4'hc == io_exe_1_rob_addr ? 1'h0 : _GEN_830; // @[Rob.scala 115:{21,21}]
  wire  _GEN_959 = 4'hd == io_exe_1_rob_addr ? 1'h0 : _GEN_831; // @[Rob.scala 115:{21,21}]
  wire  _GEN_960 = 4'he == io_exe_1_rob_addr ? 1'h0 : _GEN_832; // @[Rob.scala 115:{21,21}]
  wire  _GEN_961 = 4'hf == io_exe_1_rob_addr ? 1'h0 : _GEN_833; // @[Rob.scala 115:{21,21}]
  wire  _GEN_962 = io_exe_1_valid ? _GEN_834 : _GEN_706; // @[Rob.scala 113:28]
  wire  _GEN_963 = io_exe_1_valid ? _GEN_835 : _GEN_707; // @[Rob.scala 113:28]
  wire  _GEN_964 = io_exe_1_valid ? _GEN_836 : _GEN_708; // @[Rob.scala 113:28]
  wire  _GEN_965 = io_exe_1_valid ? _GEN_837 : _GEN_709; // @[Rob.scala 113:28]
  wire  _GEN_966 = io_exe_1_valid ? _GEN_838 : _GEN_710; // @[Rob.scala 113:28]
  wire  _GEN_967 = io_exe_1_valid ? _GEN_839 : _GEN_711; // @[Rob.scala 113:28]
  wire  _GEN_968 = io_exe_1_valid ? _GEN_840 : _GEN_712; // @[Rob.scala 113:28]
  wire  _GEN_969 = io_exe_1_valid ? _GEN_841 : _GEN_713; // @[Rob.scala 113:28]
  wire  _GEN_970 = io_exe_1_valid ? _GEN_842 : _GEN_714; // @[Rob.scala 113:28]
  wire  _GEN_971 = io_exe_1_valid ? _GEN_843 : _GEN_715; // @[Rob.scala 113:28]
  wire  _GEN_972 = io_exe_1_valid ? _GEN_844 : _GEN_716; // @[Rob.scala 113:28]
  wire  _GEN_973 = io_exe_1_valid ? _GEN_845 : _GEN_717; // @[Rob.scala 113:28]
  wire  _GEN_974 = io_exe_1_valid ? _GEN_846 : _GEN_718; // @[Rob.scala 113:28]
  wire  _GEN_975 = io_exe_1_valid ? _GEN_847 : _GEN_719; // @[Rob.scala 113:28]
  wire  _GEN_976 = io_exe_1_valid ? _GEN_848 : _GEN_720; // @[Rob.scala 113:28]
  wire  _GEN_977 = io_exe_1_valid ? _GEN_849 : _GEN_721; // @[Rob.scala 113:28]
  wire  _GEN_994 = io_exe_1_valid ? _GEN_866 : _GEN_738; // @[Rob.scala 113:28]
  wire  _GEN_995 = io_exe_1_valid ? _GEN_867 : _GEN_739; // @[Rob.scala 113:28]
  wire  _GEN_996 = io_exe_1_valid ? _GEN_868 : _GEN_740; // @[Rob.scala 113:28]
  wire  _GEN_997 = io_exe_1_valid ? _GEN_869 : _GEN_741; // @[Rob.scala 113:28]
  wire  _GEN_998 = io_exe_1_valid ? _GEN_870 : _GEN_742; // @[Rob.scala 113:28]
  wire  _GEN_999 = io_exe_1_valid ? _GEN_871 : _GEN_743; // @[Rob.scala 113:28]
  wire  _GEN_1000 = io_exe_1_valid ? _GEN_872 : _GEN_744; // @[Rob.scala 113:28]
  wire  _GEN_1001 = io_exe_1_valid ? _GEN_873 : _GEN_745; // @[Rob.scala 113:28]
  wire  _GEN_1002 = io_exe_1_valid ? _GEN_874 : _GEN_746; // @[Rob.scala 113:28]
  wire  _GEN_1003 = io_exe_1_valid ? _GEN_875 : _GEN_747; // @[Rob.scala 113:28]
  wire  _GEN_1004 = io_exe_1_valid ? _GEN_876 : _GEN_748; // @[Rob.scala 113:28]
  wire  _GEN_1005 = io_exe_1_valid ? _GEN_877 : _GEN_749; // @[Rob.scala 113:28]
  wire  _GEN_1006 = io_exe_1_valid ? _GEN_878 : _GEN_750; // @[Rob.scala 113:28]
  wire  _GEN_1007 = io_exe_1_valid ? _GEN_879 : _GEN_751; // @[Rob.scala 113:28]
  wire  _GEN_1008 = io_exe_1_valid ? _GEN_880 : _GEN_752; // @[Rob.scala 113:28]
  wire  _GEN_1009 = io_exe_1_valid ? _GEN_881 : _GEN_753; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1010 = io_exe_1_valid ? _GEN_882 : _GEN_754; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1011 = io_exe_1_valid ? _GEN_883 : _GEN_755; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1012 = io_exe_1_valid ? _GEN_884 : _GEN_756; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1013 = io_exe_1_valid ? _GEN_885 : _GEN_757; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1014 = io_exe_1_valid ? _GEN_886 : _GEN_758; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1015 = io_exe_1_valid ? _GEN_887 : _GEN_759; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1016 = io_exe_1_valid ? _GEN_888 : _GEN_760; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1017 = io_exe_1_valid ? _GEN_889 : _GEN_761; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1018 = io_exe_1_valid ? _GEN_890 : _GEN_762; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1019 = io_exe_1_valid ? _GEN_891 : _GEN_763; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1020 = io_exe_1_valid ? _GEN_892 : _GEN_764; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1021 = io_exe_1_valid ? _GEN_893 : _GEN_765; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1022 = io_exe_1_valid ? _GEN_894 : _GEN_766; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1023 = io_exe_1_valid ? _GEN_895 : _GEN_767; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1024 = io_exe_1_valid ? _GEN_896 : _GEN_768; // @[Rob.scala 113:28]
  wire [31:0] _GEN_1025 = io_exe_1_valid ? _GEN_897 : _GEN_769; // @[Rob.scala 113:28]
  wire  _GEN_1026 = io_exe_1_valid ? _GEN_898 : _GEN_770; // @[Rob.scala 113:28]
  wire  _GEN_1027 = io_exe_1_valid ? _GEN_899 : _GEN_771; // @[Rob.scala 113:28]
  wire  _GEN_1028 = io_exe_1_valid ? _GEN_900 : _GEN_772; // @[Rob.scala 113:28]
  wire  _GEN_1029 = io_exe_1_valid ? _GEN_901 : _GEN_773; // @[Rob.scala 113:28]
  wire  _GEN_1030 = io_exe_1_valid ? _GEN_902 : _GEN_774; // @[Rob.scala 113:28]
  wire  _GEN_1031 = io_exe_1_valid ? _GEN_903 : _GEN_775; // @[Rob.scala 113:28]
  wire  _GEN_1032 = io_exe_1_valid ? _GEN_904 : _GEN_776; // @[Rob.scala 113:28]
  wire  _GEN_1033 = io_exe_1_valid ? _GEN_905 : _GEN_777; // @[Rob.scala 113:28]
  wire  _GEN_1034 = io_exe_1_valid ? _GEN_906 : _GEN_778; // @[Rob.scala 113:28]
  wire  _GEN_1035 = io_exe_1_valid ? _GEN_907 : _GEN_779; // @[Rob.scala 113:28]
  wire  _GEN_1036 = io_exe_1_valid ? _GEN_908 : _GEN_780; // @[Rob.scala 113:28]
  wire  _GEN_1037 = io_exe_1_valid ? _GEN_909 : _GEN_781; // @[Rob.scala 113:28]
  wire  _GEN_1038 = io_exe_1_valid ? _GEN_910 : _GEN_782; // @[Rob.scala 113:28]
  wire  _GEN_1039 = io_exe_1_valid ? _GEN_911 : _GEN_783; // @[Rob.scala 113:28]
  wire  _GEN_1040 = io_exe_1_valid ? _GEN_912 : _GEN_784; // @[Rob.scala 113:28]
  wire  _GEN_1041 = io_exe_1_valid ? _GEN_913 : _GEN_785; // @[Rob.scala 113:28]
  wire  _GEN_1042 = io_exe_1_valid ? _GEN_914 : _GEN_786; // @[Rob.scala 113:28]
  wire  _GEN_1043 = io_exe_1_valid ? _GEN_915 : _GEN_787; // @[Rob.scala 113:28]
  wire  _GEN_1044 = io_exe_1_valid ? _GEN_916 : _GEN_788; // @[Rob.scala 113:28]
  wire  _GEN_1045 = io_exe_1_valid ? _GEN_917 : _GEN_789; // @[Rob.scala 113:28]
  wire  _GEN_1046 = io_exe_1_valid ? _GEN_918 : _GEN_790; // @[Rob.scala 113:28]
  wire  _GEN_1047 = io_exe_1_valid ? _GEN_919 : _GEN_791; // @[Rob.scala 113:28]
  wire  _GEN_1048 = io_exe_1_valid ? _GEN_920 : _GEN_792; // @[Rob.scala 113:28]
  wire  _GEN_1049 = io_exe_1_valid ? _GEN_921 : _GEN_793; // @[Rob.scala 113:28]
  wire  _GEN_1050 = io_exe_1_valid ? _GEN_922 : _GEN_794; // @[Rob.scala 113:28]
  wire  _GEN_1051 = io_exe_1_valid ? _GEN_923 : _GEN_795; // @[Rob.scala 113:28]
  wire  _GEN_1052 = io_exe_1_valid ? _GEN_924 : _GEN_796; // @[Rob.scala 113:28]
  wire  _GEN_1053 = io_exe_1_valid ? _GEN_925 : _GEN_797; // @[Rob.scala 113:28]
  wire  _GEN_1054 = io_exe_1_valid ? _GEN_926 : _GEN_798; // @[Rob.scala 113:28]
  wire  _GEN_1055 = io_exe_1_valid ? _GEN_927 : _GEN_799; // @[Rob.scala 113:28]
  wire  _GEN_1056 = io_exe_1_valid ? _GEN_928 : _GEN_800; // @[Rob.scala 113:28]
  wire  _GEN_1057 = io_exe_1_valid ? _GEN_929 : _GEN_801; // @[Rob.scala 113:28]
  wire  _GEN_1074 = io_exe_1_valid ? _GEN_946 : _GEN_818; // @[Rob.scala 113:28]
  wire  _GEN_1075 = io_exe_1_valid ? _GEN_947 : _GEN_819; // @[Rob.scala 113:28]
  wire  _GEN_1076 = io_exe_1_valid ? _GEN_948 : _GEN_820; // @[Rob.scala 113:28]
  wire  _GEN_1077 = io_exe_1_valid ? _GEN_949 : _GEN_821; // @[Rob.scala 113:28]
  wire  _GEN_1078 = io_exe_1_valid ? _GEN_950 : _GEN_822; // @[Rob.scala 113:28]
  wire  _GEN_1079 = io_exe_1_valid ? _GEN_951 : _GEN_823; // @[Rob.scala 113:28]
  wire  _GEN_1080 = io_exe_1_valid ? _GEN_952 : _GEN_824; // @[Rob.scala 113:28]
  wire  _GEN_1081 = io_exe_1_valid ? _GEN_953 : _GEN_825; // @[Rob.scala 113:28]
  wire  _GEN_1082 = io_exe_1_valid ? _GEN_954 : _GEN_826; // @[Rob.scala 113:28]
  wire  _GEN_1083 = io_exe_1_valid ? _GEN_955 : _GEN_827; // @[Rob.scala 113:28]
  wire  _GEN_1084 = io_exe_1_valid ? _GEN_956 : _GEN_828; // @[Rob.scala 113:28]
  wire  _GEN_1085 = io_exe_1_valid ? _GEN_957 : _GEN_829; // @[Rob.scala 113:28]
  wire  _GEN_1086 = io_exe_1_valid ? _GEN_958 : _GEN_830; // @[Rob.scala 113:28]
  wire  _GEN_1087 = io_exe_1_valid ? _GEN_959 : _GEN_831; // @[Rob.scala 113:28]
  wire  _GEN_1088 = io_exe_1_valid ? _GEN_960 : _GEN_832; // @[Rob.scala 113:28]
  wire  _GEN_1089 = io_exe_1_valid ? _GEN_961 : _GEN_833; // @[Rob.scala 113:28]
  wire  _GEN_1090 = 4'h0 == io_exe_2_rob_addr | _GEN_962; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1091 = 4'h1 == io_exe_2_rob_addr | _GEN_963; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1092 = 4'h2 == io_exe_2_rob_addr | _GEN_964; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1093 = 4'h3 == io_exe_2_rob_addr | _GEN_965; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1094 = 4'h4 == io_exe_2_rob_addr | _GEN_966; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1095 = 4'h5 == io_exe_2_rob_addr | _GEN_967; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1096 = 4'h6 == io_exe_2_rob_addr | _GEN_968; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1097 = 4'h7 == io_exe_2_rob_addr | _GEN_969; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1098 = 4'h8 == io_exe_2_rob_addr | _GEN_970; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1099 = 4'h9 == io_exe_2_rob_addr | _GEN_971; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1100 = 4'ha == io_exe_2_rob_addr | _GEN_972; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1101 = 4'hb == io_exe_2_rob_addr | _GEN_973; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1102 = 4'hc == io_exe_2_rob_addr | _GEN_974; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1103 = 4'hd == io_exe_2_rob_addr | _GEN_975; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1104 = 4'he == io_exe_2_rob_addr | _GEN_976; // @[Rob.scala 114:{26,26}]
  wire  _GEN_1105 = 4'hf == io_exe_2_rob_addr | _GEN_977; // @[Rob.scala 114:{26,26}]
  wire [4:0] _GEN_2275 = {{3'd0}, num_deq}; // @[Rob.scala 122:44]
  wire [4:0] next_deq_vec_0 = deq_vec_0 + _GEN_2275; // @[Rob.scala 122:44]
  wire [4:0] next_deq_vec_1 = deq_vec_1 + _GEN_2275; // @[Rob.scala 122:44]
  reg  sys_in_flight; // @[Rob.scala 152:30]
  reg  intr_state; // @[Rob.scala 183:27]
  wire  intr_global_en = csr_mstatus_0[3]; // @[Rob.scala 187:36]
  wire  _T_49 = intr_global_en & csr_mie_mtie_0; // @[Rob.scala 192:28]
  wire  _GEN_1378 = intr_global_en & csr_mie_mtie_0 | intr_state; // @[Rob.scala 192:46 193:20 183:27]
  wire  _T_53 = ~sys_in_flight; // @[Rob.scala 198:51]
  wire  _T_54 = cm_0_valid & csr_mip_mtip_intr_0 & ~sys_in_flight; // @[Rob.scala 198:48]
  wire [63:0] _T_59 = {csr_mstatus_0[63:8],intr_global_en,csr_mstatus_0[6:4],1'h0,csr_mstatus_0[2:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_61 = {csr_mtvec_idx_0,2'h0}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_1379 = cm_0_valid & csr_mip_mtip_intr_0 & ~sys_in_flight ? _T_59 : 64'h1800; // @[Rob.scala 198:67 199:24]
  wire [31:0] deq_uop_0_pc = rob_pc_MPORT_2_data; // @[Rob.scala 156:21 229:16]
  wire [31:0] _GEN_1380 = cm_0_valid & csr_mip_mtip_intr_0 & ~sys_in_flight ? deq_uop_0_pc : 32'h0; // @[Rob.scala 198:67 200:21]
  wire [63:0] _GEN_1381 = cm_0_valid & csr_mip_mtip_intr_0 & ~sys_in_flight ? 64'h8000000000000007 : 64'h0; // @[Rob.scala 198:67 201:23]
  wire [31:0] _GEN_1383 = cm_0_valid & csr_mip_mtip_intr_0 & ~sys_in_flight ? _T_61 : 32'h0; // @[Rob.scala 198:67 203:23]
  wire  _GEN_1384 = cm_0_valid & csr_mip_mtip_intr_0 & ~sys_in_flight ? 1'h0 : intr_state; // @[Rob.scala 198:67 204:22 183:27]
  wire [63:0] _GEN_1385 = _T_49 ? _GEN_1379 : 64'h1800; // @[Rob.scala 197:46]
  wire [31:0] _GEN_1386 = _T_49 ? _GEN_1380 : 32'h0; // @[Rob.scala 197:46]
  wire [63:0] _GEN_1387 = _T_49 ? _GEN_1381 : 64'h0; // @[Rob.scala 197:46]
  wire  _GEN_1388 = _T_49 & _T_54; // @[Rob.scala 197:46]
  wire [31:0] _GEN_1389 = _T_49 ? _GEN_1383 : 32'h0; // @[Rob.scala 197:46]
  wire  _GEN_1390 = _T_49 & _GEN_1384; // @[Rob.scala 197:46 207:20]
  wire [63:0] _GEN_1391 = intr_state ? _GEN_1385 : 64'h1800; // @[Rob.scala 190:23]
  wire [31:0] _GEN_1392 = intr_state ? _GEN_1386 : 32'h0; // @[Rob.scala 190:23]
  wire [63:0] _GEN_1393 = intr_state ? _GEN_1387 : 64'h0; // @[Rob.scala 190:23]
  wire [31:0] _GEN_1395 = intr_state ? _GEN_1389 : 32'h0; // @[Rob.scala 190:23]
  wire [31:0] _GEN_1399 = ~intr_state ? 32'h0 : _GEN_1392; // @[Rob.scala 190:23]
  wire [31:0] intr_jmp_pc = ~intr_state ? 32'h0 : _GEN_1395; // @[Rob.scala 190:23]
  wire [31:0] _GEN_1440 = 4'h1 == deq_ptr ? ecp_1_jmp_pc : ecp_0_jmp_pc; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1441 = 4'h2 == deq_ptr ? ecp_2_jmp_pc : _GEN_1440; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1442 = 4'h3 == deq_ptr ? ecp_3_jmp_pc : _GEN_1441; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1443 = 4'h4 == deq_ptr ? ecp_4_jmp_pc : _GEN_1442; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1444 = 4'h5 == deq_ptr ? ecp_5_jmp_pc : _GEN_1443; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1445 = 4'h6 == deq_ptr ? ecp_6_jmp_pc : _GEN_1444; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1446 = 4'h7 == deq_ptr ? ecp_7_jmp_pc : _GEN_1445; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1447 = 4'h8 == deq_ptr ? ecp_8_jmp_pc : _GEN_1446; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1448 = 4'h9 == deq_ptr ? ecp_9_jmp_pc : _GEN_1447; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1449 = 4'ha == deq_ptr ? ecp_10_jmp_pc : _GEN_1448; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1450 = 4'hb == deq_ptr ? ecp_11_jmp_pc : _GEN_1449; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1451 = 4'hc == deq_ptr ? ecp_12_jmp_pc : _GEN_1450; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1452 = 4'hd == deq_ptr ? ecp_13_jmp_pc : _GEN_1451; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1453 = 4'he == deq_ptr ? ecp_14_jmp_pc : _GEN_1452; // @[Rob.scala 231:{16,16}]
  wire [31:0] deq_ecp_0_jmp_pc = 4'hf == deq_ptr ? ecp_15_jmp_pc : _GEN_1453; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1456 = 4'h1 == deq_ptr ? ecp_1_jmp : ecp_0_jmp; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1457 = 4'h2 == deq_ptr ? ecp_2_jmp : _GEN_1456; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1458 = 4'h3 == deq_ptr ? ecp_3_jmp : _GEN_1457; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1459 = 4'h4 == deq_ptr ? ecp_4_jmp : _GEN_1458; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1460 = 4'h5 == deq_ptr ? ecp_5_jmp : _GEN_1459; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1461 = 4'h6 == deq_ptr ? ecp_6_jmp : _GEN_1460; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1462 = 4'h7 == deq_ptr ? ecp_7_jmp : _GEN_1461; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1463 = 4'h8 == deq_ptr ? ecp_8_jmp : _GEN_1462; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1464 = 4'h9 == deq_ptr ? ecp_9_jmp : _GEN_1463; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1465 = 4'ha == deq_ptr ? ecp_10_jmp : _GEN_1464; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1466 = 4'hb == deq_ptr ? ecp_11_jmp : _GEN_1465; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1467 = 4'hc == deq_ptr ? ecp_12_jmp : _GEN_1466; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1468 = 4'hd == deq_ptr ? ecp_13_jmp : _GEN_1467; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1469 = 4'he == deq_ptr ? ecp_14_jmp : _GEN_1468; // @[Rob.scala 231:{16,16}]
  wire  deq_ecp_0_jmp = 4'hf == deq_ptr ? ecp_15_jmp : _GEN_1469; // @[Rob.scala 231:{16,16}]
  wire [2:0] deq_uop_0_fu_code = rob_fu_code_MPORT_2_data; // @[Rob.scala 156:21 229:16]
  wire  _T_66 = deq_uop_0_fu_code == 3'h3; // @[Rob.scala 233:32]
  wire  _GEN_1520 = deq_uop_0_fu_code == 3'h3 & _T_53 & ~rob_empty | sys_in_flight; // @[Rob.scala 233:83 235:23 152:30]
  wire  jmp_1h_0 = deq_ecp_0_jmp_valid & cm_0_valid; // @[Rob.scala 275:31]
  wire [2:0] deq_uop_0_sys_code = rob_sys_code_MPORT_2_data; // @[Rob.scala 156:21 229:16]
  wire  _T_79 = deq_uop_0_sys_code == 3'h7; // @[Rob.scala 283:53]
  wire [31:0] _GEN_1527 = jmp_1h_0 ? deq_uop_0_pc : 32'h0; // @[Rob.scala 143:17 276:22 278:29]
  wire  _GEN_1528 = jmp_1h_0 & deq_ecp_0_jmp; // @[Rob.scala 143:17 276:22 279:29]
  wire [31:0] _GEN_1529 = jmp_1h_0 ? deq_ecp_0_jmp_pc : 32'h0; // @[Rob.scala 143:17 276:22 280:29]
  wire  _GEN_1530 = jmp_1h_0 & deq_ecp_0_mis; // @[Rob.scala 143:17 276:22 281:29]
  wire  _GEN_1531 = jmp_1h_0 & (_T_66 & _T_79); // @[Rob.scala 143:17 276:22 282:29]
  wire  _GEN_1554 = 4'h1 == deq_vec_1[3:0] ? ecp_1_mis : ecp_0_mis; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1555 = 4'h2 == deq_vec_1[3:0] ? ecp_2_mis : _GEN_1554; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1556 = 4'h3 == deq_vec_1[3:0] ? ecp_3_mis : _GEN_1555; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1557 = 4'h4 == deq_vec_1[3:0] ? ecp_4_mis : _GEN_1556; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1558 = 4'h5 == deq_vec_1[3:0] ? ecp_5_mis : _GEN_1557; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1559 = 4'h6 == deq_vec_1[3:0] ? ecp_6_mis : _GEN_1558; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1560 = 4'h7 == deq_vec_1[3:0] ? ecp_7_mis : _GEN_1559; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1561 = 4'h8 == deq_vec_1[3:0] ? ecp_8_mis : _GEN_1560; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1562 = 4'h9 == deq_vec_1[3:0] ? ecp_9_mis : _GEN_1561; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1563 = 4'ha == deq_vec_1[3:0] ? ecp_10_mis : _GEN_1562; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1564 = 4'hb == deq_vec_1[3:0] ? ecp_11_mis : _GEN_1563; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1565 = 4'hc == deq_vec_1[3:0] ? ecp_12_mis : _GEN_1564; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1566 = 4'hd == deq_vec_1[3:0] ? ecp_13_mis : _GEN_1565; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1567 = 4'he == deq_vec_1[3:0] ? ecp_14_mis : _GEN_1566; // @[Rob.scala 231:{16,16}]
  wire  deq_ecp_1_mis = 4'hf == deq_vec_1[3:0] ? ecp_15_mis : _GEN_1567; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1570 = 4'h1 == deq_vec_1[3:0] ? ecp_1_jmp_pc : ecp_0_jmp_pc; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1571 = 4'h2 == deq_vec_1[3:0] ? ecp_2_jmp_pc : _GEN_1570; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1572 = 4'h3 == deq_vec_1[3:0] ? ecp_3_jmp_pc : _GEN_1571; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1573 = 4'h4 == deq_vec_1[3:0] ? ecp_4_jmp_pc : _GEN_1572; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1574 = 4'h5 == deq_vec_1[3:0] ? ecp_5_jmp_pc : _GEN_1573; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1575 = 4'h6 == deq_vec_1[3:0] ? ecp_6_jmp_pc : _GEN_1574; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1576 = 4'h7 == deq_vec_1[3:0] ? ecp_7_jmp_pc : _GEN_1575; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1577 = 4'h8 == deq_vec_1[3:0] ? ecp_8_jmp_pc : _GEN_1576; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1578 = 4'h9 == deq_vec_1[3:0] ? ecp_9_jmp_pc : _GEN_1577; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1579 = 4'ha == deq_vec_1[3:0] ? ecp_10_jmp_pc : _GEN_1578; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1580 = 4'hb == deq_vec_1[3:0] ? ecp_11_jmp_pc : _GEN_1579; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1581 = 4'hc == deq_vec_1[3:0] ? ecp_12_jmp_pc : _GEN_1580; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1582 = 4'hd == deq_vec_1[3:0] ? ecp_13_jmp_pc : _GEN_1581; // @[Rob.scala 231:{16,16}]
  wire [31:0] _GEN_1583 = 4'he == deq_vec_1[3:0] ? ecp_14_jmp_pc : _GEN_1582; // @[Rob.scala 231:{16,16}]
  wire [31:0] deq_ecp_1_jmp_pc = 4'hf == deq_vec_1[3:0] ? ecp_15_jmp_pc : _GEN_1583; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1586 = 4'h1 == deq_vec_1[3:0] ? ecp_1_jmp : ecp_0_jmp; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1587 = 4'h2 == deq_vec_1[3:0] ? ecp_2_jmp : _GEN_1586; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1588 = 4'h3 == deq_vec_1[3:0] ? ecp_3_jmp : _GEN_1587; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1589 = 4'h4 == deq_vec_1[3:0] ? ecp_4_jmp : _GEN_1588; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1590 = 4'h5 == deq_vec_1[3:0] ? ecp_5_jmp : _GEN_1589; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1591 = 4'h6 == deq_vec_1[3:0] ? ecp_6_jmp : _GEN_1590; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1592 = 4'h7 == deq_vec_1[3:0] ? ecp_7_jmp : _GEN_1591; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1593 = 4'h8 == deq_vec_1[3:0] ? ecp_8_jmp : _GEN_1592; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1594 = 4'h9 == deq_vec_1[3:0] ? ecp_9_jmp : _GEN_1593; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1595 = 4'ha == deq_vec_1[3:0] ? ecp_10_jmp : _GEN_1594; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1596 = 4'hb == deq_vec_1[3:0] ? ecp_11_jmp : _GEN_1595; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1597 = 4'hc == deq_vec_1[3:0] ? ecp_12_jmp : _GEN_1596; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1598 = 4'hd == deq_vec_1[3:0] ? ecp_13_jmp : _GEN_1597; // @[Rob.scala 231:{16,16}]
  wire  _GEN_1599 = 4'he == deq_vec_1[3:0] ? ecp_14_jmp : _GEN_1598; // @[Rob.scala 231:{16,16}]
  wire  deq_ecp_1_jmp = 4'hf == deq_vec_1[3:0] ? ecp_15_jmp : _GEN_1599; // @[Rob.scala 231:{16,16}]
  wire  sq_deq_req = cm_1_valid & deq_ecp_1_store_valid | cm_0_valid & deq_ecp_0_store_valid; // @[Rob.scala 270:42 271:18]
  wire  jmp_1h_1 = deq_ecp_1_jmp_valid & cm_1_valid; // @[Rob.scala 275:31]
  wire [2:0] deq_uop_1_fu_code = rob_fu_code_MPORT_3_data; // @[Rob.scala 156:21 229:16]
  wire [2:0] deq_uop_1_sys_code = rob_sys_code_MPORT_3_data; // @[Rob.scala 156:21 229:16]
  wire  _T_121 = deq_uop_1_sys_code == 3'h7; // @[Rob.scala 283:53]
  wire  _GEN_1654 = jmp_1h_1 | jmp_1h_0; // @[Rob.scala 276:22 277:29]
  wire [31:0] deq_uop_1_pc = rob_pc_MPORT_3_data; // @[Rob.scala 156:21 229:16]
  wire [31:0] _GEN_1655 = jmp_1h_1 ? deq_uop_1_pc : _GEN_1527; // @[Rob.scala 276:22 278:29]
  wire  _GEN_1656 = jmp_1h_1 ? deq_ecp_1_jmp : _GEN_1528; // @[Rob.scala 276:22 279:29]
  wire [31:0] _GEN_1657 = jmp_1h_1 ? deq_ecp_1_jmp_pc : _GEN_1529; // @[Rob.scala 276:22 280:29]
  wire  _GEN_1658 = jmp_1h_1 ? deq_ecp_1_mis : _GEN_1530; // @[Rob.scala 276:22 281:29]
  wire  _GEN_1659 = jmp_1h_1 ? deq_uop_1_fu_code == 3'h3 & _T_121 : _GEN_1531; // @[Rob.scala 276:22 282:29]
  wire [63:0] intr_mepc = {{32'd0}, _GEN_1399};
  wire  intr = ~intr_state ? 1'h0 : intr_state & _GEN_1388; // @[Rob.scala 190:23]
  wire  _GEN_1671 = io_flush | 6'he >= next_valid_entry; // @[Rob.scala 332:19 333:15 66:13]
  wire  _T_142 = ~intr; // @[Rob.scala 352:38]
  wire [63:0] intr_mstatus = ~intr_state ? 64'h1800 : _GEN_1391; // @[Rob.scala 190:23]
  wire [63:0] intr_mcause = ~intr_state ? 64'h0 : _GEN_1393; // @[Rob.scala 190:23]
//   assign rob_pc_MPORT_2_en = rob_pc_MPORT_2_en_pipe_0;
  assign rob_pc_MPORT_2_addr = rob_pc_MPORT_2_addr_pipe_0;
  assign rob_pc_MPORT_2_data = rob_pc[rob_pc_MPORT_2_addr]; // @[Rob.scala 44:24]
//   assign rob_pc_MPORT_3_en = rob_pc_MPORT_3_en_pipe_0;
  assign rob_pc_MPORT_3_addr = rob_pc_MPORT_3_addr_pipe_0;
  assign rob_pc_MPORT_3_data = rob_pc[rob_pc_MPORT_3_addr]; // @[Rob.scala 44:24]
  assign rob_pc_MPORT_data = io_in_bits_vec_0_pc;
  assign rob_pc_MPORT_addr = enq_vec_0[3:0];
  assign rob_pc_MPORT_mask = 1'h1;
  assign rob_pc_MPORT_en = _T_20 & _T_21;
  assign rob_pc_MPORT_1_data = io_in_bits_vec_1_pc;
  assign rob_pc_MPORT_1_addr = _GEN_289[3:0];
  assign rob_pc_MPORT_1_mask = 1'h1;
  assign rob_pc_MPORT_1_en = _T_25 & _T_21;
  assign rob_pc_MPORT_4_data = 32'h0;
  assign rob_pc_MPORT_4_addr = 4'h0;
  assign rob_pc_MPORT_4_mask = 1'h1;
  assign rob_pc_MPORT_4_en = reset;
  assign rob_pc_MPORT_5_data = 32'h0;
  assign rob_pc_MPORT_5_addr = 4'h1;
  assign rob_pc_MPORT_5_mask = 1'h1;
  assign rob_pc_MPORT_5_en = reset;
  assign rob_pc_MPORT_6_data = 32'h0;
  assign rob_pc_MPORT_6_addr = 4'h2;
  assign rob_pc_MPORT_6_mask = 1'h1;
  assign rob_pc_MPORT_6_en = reset;
  assign rob_pc_MPORT_7_data = 32'h0;
  assign rob_pc_MPORT_7_addr = 4'h3;
  assign rob_pc_MPORT_7_mask = 1'h1;
  assign rob_pc_MPORT_7_en = reset;
  assign rob_pc_MPORT_8_data = 32'h0;
  assign rob_pc_MPORT_8_addr = 4'h4;
  assign rob_pc_MPORT_8_mask = 1'h1;
  assign rob_pc_MPORT_8_en = reset;
  assign rob_pc_MPORT_9_data = 32'h0;
  assign rob_pc_MPORT_9_addr = 4'h5;
  assign rob_pc_MPORT_9_mask = 1'h1;
  assign rob_pc_MPORT_9_en = reset;
  assign rob_pc_MPORT_10_data = 32'h0;
  assign rob_pc_MPORT_10_addr = 4'h6;
  assign rob_pc_MPORT_10_mask = 1'h1;
  assign rob_pc_MPORT_10_en = reset;
  assign rob_pc_MPORT_11_data = 32'h0;
  assign rob_pc_MPORT_11_addr = 4'h7;
  assign rob_pc_MPORT_11_mask = 1'h1;
  assign rob_pc_MPORT_11_en = reset;
  assign rob_pc_MPORT_12_data = 32'h0;
  assign rob_pc_MPORT_12_addr = 4'h8;
  assign rob_pc_MPORT_12_mask = 1'h1;
  assign rob_pc_MPORT_12_en = reset;
  assign rob_pc_MPORT_13_data = 32'h0;
  assign rob_pc_MPORT_13_addr = 4'h9;
  assign rob_pc_MPORT_13_mask = 1'h1;
  assign rob_pc_MPORT_13_en = reset;
  assign rob_pc_MPORT_14_data = 32'h0;
  assign rob_pc_MPORT_14_addr = 4'ha;
  assign rob_pc_MPORT_14_mask = 1'h1;
  assign rob_pc_MPORT_14_en = reset;
  assign rob_pc_MPORT_15_data = 32'h0;
  assign rob_pc_MPORT_15_addr = 4'hb;
  assign rob_pc_MPORT_15_mask = 1'h1;
  assign rob_pc_MPORT_15_en = reset;
  assign rob_pc_MPORT_16_data = 32'h0;
  assign rob_pc_MPORT_16_addr = 4'hc;
  assign rob_pc_MPORT_16_mask = 1'h1;
  assign rob_pc_MPORT_16_en = reset;
  assign rob_pc_MPORT_17_data = 32'h0;
  assign rob_pc_MPORT_17_addr = 4'hd;
  assign rob_pc_MPORT_17_mask = 1'h1;
  assign rob_pc_MPORT_17_en = reset;
  assign rob_pc_MPORT_18_data = 32'h0;
  assign rob_pc_MPORT_18_addr = 4'he;
  assign rob_pc_MPORT_18_mask = 1'h1;
  assign rob_pc_MPORT_18_en = reset;
  assign rob_pc_MPORT_19_data = 32'h0;
  assign rob_pc_MPORT_19_addr = 4'hf;
  assign rob_pc_MPORT_19_mask = 1'h1;
  assign rob_pc_MPORT_19_en = reset;
//   assign rob_fu_code_MPORT_2_en = rob_fu_code_MPORT_2_en_pipe_0;
  assign rob_fu_code_MPORT_2_addr = rob_fu_code_MPORT_2_addr_pipe_0;
  assign rob_fu_code_MPORT_2_data = rob_fu_code[rob_fu_code_MPORT_2_addr]; // @[Rob.scala 44:24]
//   assign rob_fu_code_MPORT_3_en = rob_fu_code_MPORT_3_en_pipe_0;
  assign rob_fu_code_MPORT_3_addr = rob_fu_code_MPORT_3_addr_pipe_0;
  assign rob_fu_code_MPORT_3_data = rob_fu_code[rob_fu_code_MPORT_3_addr]; // @[Rob.scala 44:24]
  assign rob_fu_code_MPORT_data = io_in_bits_vec_0_fu_code;
  assign rob_fu_code_MPORT_addr = enq_vec_0[3:0];
  assign rob_fu_code_MPORT_mask = 1'h1;
  assign rob_fu_code_MPORT_en = _T_20 & _T_21;
  assign rob_fu_code_MPORT_1_data = io_in_bits_vec_1_fu_code;
  assign rob_fu_code_MPORT_1_addr = _GEN_289[3:0];
  assign rob_fu_code_MPORT_1_mask = 1'h1;
  assign rob_fu_code_MPORT_1_en = _T_25 & _T_21;
  assign rob_fu_code_MPORT_4_data = 3'h0;
  assign rob_fu_code_MPORT_4_addr = 4'h0;
  assign rob_fu_code_MPORT_4_mask = 1'h1;
  assign rob_fu_code_MPORT_4_en = reset;
  assign rob_fu_code_MPORT_5_data = 3'h0;
  assign rob_fu_code_MPORT_5_addr = 4'h1;
  assign rob_fu_code_MPORT_5_mask = 1'h1;
  assign rob_fu_code_MPORT_5_en = reset;
  assign rob_fu_code_MPORT_6_data = 3'h0;
  assign rob_fu_code_MPORT_6_addr = 4'h2;
  assign rob_fu_code_MPORT_6_mask = 1'h1;
  assign rob_fu_code_MPORT_6_en = reset;
  assign rob_fu_code_MPORT_7_data = 3'h0;
  assign rob_fu_code_MPORT_7_addr = 4'h3;
  assign rob_fu_code_MPORT_7_mask = 1'h1;
  assign rob_fu_code_MPORT_7_en = reset;
  assign rob_fu_code_MPORT_8_data = 3'h0;
  assign rob_fu_code_MPORT_8_addr = 4'h4;
  assign rob_fu_code_MPORT_8_mask = 1'h1;
  assign rob_fu_code_MPORT_8_en = reset;
  assign rob_fu_code_MPORT_9_data = 3'h0;
  assign rob_fu_code_MPORT_9_addr = 4'h5;
  assign rob_fu_code_MPORT_9_mask = 1'h1;
  assign rob_fu_code_MPORT_9_en = reset;
  assign rob_fu_code_MPORT_10_data = 3'h0;
  assign rob_fu_code_MPORT_10_addr = 4'h6;
  assign rob_fu_code_MPORT_10_mask = 1'h1;
  assign rob_fu_code_MPORT_10_en = reset;
  assign rob_fu_code_MPORT_11_data = 3'h0;
  assign rob_fu_code_MPORT_11_addr = 4'h7;
  assign rob_fu_code_MPORT_11_mask = 1'h1;
  assign rob_fu_code_MPORT_11_en = reset;
  assign rob_fu_code_MPORT_12_data = 3'h0;
  assign rob_fu_code_MPORT_12_addr = 4'h8;
  assign rob_fu_code_MPORT_12_mask = 1'h1;
  assign rob_fu_code_MPORT_12_en = reset;
  assign rob_fu_code_MPORT_13_data = 3'h0;
  assign rob_fu_code_MPORT_13_addr = 4'h9;
  assign rob_fu_code_MPORT_13_mask = 1'h1;
  assign rob_fu_code_MPORT_13_en = reset;
  assign rob_fu_code_MPORT_14_data = 3'h0;
  assign rob_fu_code_MPORT_14_addr = 4'ha;
  assign rob_fu_code_MPORT_14_mask = 1'h1;
  assign rob_fu_code_MPORT_14_en = reset;
  assign rob_fu_code_MPORT_15_data = 3'h0;
  assign rob_fu_code_MPORT_15_addr = 4'hb;
  assign rob_fu_code_MPORT_15_mask = 1'h1;
  assign rob_fu_code_MPORT_15_en = reset;
  assign rob_fu_code_MPORT_16_data = 3'h0;
  assign rob_fu_code_MPORT_16_addr = 4'hc;
  assign rob_fu_code_MPORT_16_mask = 1'h1;
  assign rob_fu_code_MPORT_16_en = reset;
  assign rob_fu_code_MPORT_17_data = 3'h0;
  assign rob_fu_code_MPORT_17_addr = 4'hd;
  assign rob_fu_code_MPORT_17_mask = 1'h1;
  assign rob_fu_code_MPORT_17_en = reset;
  assign rob_fu_code_MPORT_18_data = 3'h0;
  assign rob_fu_code_MPORT_18_addr = 4'he;
  assign rob_fu_code_MPORT_18_mask = 1'h1;
  assign rob_fu_code_MPORT_18_en = reset;
  assign rob_fu_code_MPORT_19_data = 3'h0;
  assign rob_fu_code_MPORT_19_addr = 4'hf;
  assign rob_fu_code_MPORT_19_mask = 1'h1;
  assign rob_fu_code_MPORT_19_en = reset;
//   assign rob_sys_code_MPORT_2_en = rob_sys_code_MPORT_2_en_pipe_0;
  assign rob_sys_code_MPORT_2_addr = rob_sys_code_MPORT_2_addr_pipe_0;
  assign rob_sys_code_MPORT_2_data = rob_sys_code[rob_sys_code_MPORT_2_addr]; // @[Rob.scala 44:24]
//   assign rob_sys_code_MPORT_3_en = rob_sys_code_MPORT_3_en_pipe_0;
  assign rob_sys_code_MPORT_3_addr = rob_sys_code_MPORT_3_addr_pipe_0;
  assign rob_sys_code_MPORT_3_data = rob_sys_code[rob_sys_code_MPORT_3_addr]; // @[Rob.scala 44:24]
  assign rob_sys_code_MPORT_data = io_in_bits_vec_0_sys_code;
  assign rob_sys_code_MPORT_addr = enq_vec_0[3:0];
  assign rob_sys_code_MPORT_mask = 1'h1;
  assign rob_sys_code_MPORT_en = _T_20 & _T_21;
  assign rob_sys_code_MPORT_1_data = io_in_bits_vec_1_sys_code;
  assign rob_sys_code_MPORT_1_addr = _GEN_289[3:0];
  assign rob_sys_code_MPORT_1_mask = 1'h1;
  assign rob_sys_code_MPORT_1_en = _T_25 & _T_21;
  assign rob_sys_code_MPORT_4_data = 3'h0;
  assign rob_sys_code_MPORT_4_addr = 4'h0;
  assign rob_sys_code_MPORT_4_mask = 1'h1;
  assign rob_sys_code_MPORT_4_en = reset;
  assign rob_sys_code_MPORT_5_data = 3'h0;
  assign rob_sys_code_MPORT_5_addr = 4'h1;
  assign rob_sys_code_MPORT_5_mask = 1'h1;
  assign rob_sys_code_MPORT_5_en = reset;
  assign rob_sys_code_MPORT_6_data = 3'h0;
  assign rob_sys_code_MPORT_6_addr = 4'h2;
  assign rob_sys_code_MPORT_6_mask = 1'h1;
  assign rob_sys_code_MPORT_6_en = reset;
  assign rob_sys_code_MPORT_7_data = 3'h0;
  assign rob_sys_code_MPORT_7_addr = 4'h3;
  assign rob_sys_code_MPORT_7_mask = 1'h1;
  assign rob_sys_code_MPORT_7_en = reset;
  assign rob_sys_code_MPORT_8_data = 3'h0;
  assign rob_sys_code_MPORT_8_addr = 4'h4;
  assign rob_sys_code_MPORT_8_mask = 1'h1;
  assign rob_sys_code_MPORT_8_en = reset;
  assign rob_sys_code_MPORT_9_data = 3'h0;
  assign rob_sys_code_MPORT_9_addr = 4'h5;
  assign rob_sys_code_MPORT_9_mask = 1'h1;
  assign rob_sys_code_MPORT_9_en = reset;
  assign rob_sys_code_MPORT_10_data = 3'h0;
  assign rob_sys_code_MPORT_10_addr = 4'h6;
  assign rob_sys_code_MPORT_10_mask = 1'h1;
  assign rob_sys_code_MPORT_10_en = reset;
  assign rob_sys_code_MPORT_11_data = 3'h0;
  assign rob_sys_code_MPORT_11_addr = 4'h7;
  assign rob_sys_code_MPORT_11_mask = 1'h1;
  assign rob_sys_code_MPORT_11_en = reset;
  assign rob_sys_code_MPORT_12_data = 3'h0;
  assign rob_sys_code_MPORT_12_addr = 4'h8;
  assign rob_sys_code_MPORT_12_mask = 1'h1;
  assign rob_sys_code_MPORT_12_en = reset;
  assign rob_sys_code_MPORT_13_data = 3'h0;
  assign rob_sys_code_MPORT_13_addr = 4'h9;
  assign rob_sys_code_MPORT_13_mask = 1'h1;
  assign rob_sys_code_MPORT_13_en = reset;
  assign rob_sys_code_MPORT_14_data = 3'h0;
  assign rob_sys_code_MPORT_14_addr = 4'ha;
  assign rob_sys_code_MPORT_14_mask = 1'h1;
  assign rob_sys_code_MPORT_14_en = reset;
  assign rob_sys_code_MPORT_15_data = 3'h0;
  assign rob_sys_code_MPORT_15_addr = 4'hb;
  assign rob_sys_code_MPORT_15_mask = 1'h1;
  assign rob_sys_code_MPORT_15_en = reset;
  assign rob_sys_code_MPORT_16_data = 3'h0;
  assign rob_sys_code_MPORT_16_addr = 4'hc;
  assign rob_sys_code_MPORT_16_mask = 1'h1;
  assign rob_sys_code_MPORT_16_en = reset;
  assign rob_sys_code_MPORT_17_data = 3'h0;
  assign rob_sys_code_MPORT_17_addr = 4'hd;
  assign rob_sys_code_MPORT_17_mask = 1'h1;
  assign rob_sys_code_MPORT_17_en = reset;
  assign rob_sys_code_MPORT_18_data = 3'h0;
  assign rob_sys_code_MPORT_18_addr = 4'he;
  assign rob_sys_code_MPORT_18_mask = 1'h1;
  assign rob_sys_code_MPORT_18_en = reset;
  assign rob_sys_code_MPORT_19_data = 3'h0;
  assign rob_sys_code_MPORT_19_addr = 4'hf;
  assign rob_sys_code_MPORT_19_mask = 1'h1;
  assign rob_sys_code_MPORT_19_en = reset;
//   assign rob_rd_addr_MPORT_2_en = rob_rd_addr_MPORT_2_en_pipe_0;
  assign rob_rd_addr_MPORT_2_addr = rob_rd_addr_MPORT_2_addr_pipe_0;
  assign rob_rd_addr_MPORT_2_data = rob_rd_addr[rob_rd_addr_MPORT_2_addr]; // @[Rob.scala 44:24]
//   assign rob_rd_addr_MPORT_3_en = rob_rd_addr_MPORT_3_en_pipe_0;
  assign rob_rd_addr_MPORT_3_addr = rob_rd_addr_MPORT_3_addr_pipe_0;
  assign rob_rd_addr_MPORT_3_data = rob_rd_addr[rob_rd_addr_MPORT_3_addr]; // @[Rob.scala 44:24]
  assign rob_rd_addr_MPORT_data = io_in_bits_vec_0_rd_addr;
  assign rob_rd_addr_MPORT_addr = enq_vec_0[3:0];
  assign rob_rd_addr_MPORT_mask = 1'h1;
  assign rob_rd_addr_MPORT_en = _T_20 & _T_21;
  assign rob_rd_addr_MPORT_1_data = io_in_bits_vec_1_rd_addr;
  assign rob_rd_addr_MPORT_1_addr = _GEN_289[3:0];
  assign rob_rd_addr_MPORT_1_mask = 1'h1;
  assign rob_rd_addr_MPORT_1_en = _T_25 & _T_21;
  assign rob_rd_addr_MPORT_4_data = 5'h0;
  assign rob_rd_addr_MPORT_4_addr = 4'h0;
  assign rob_rd_addr_MPORT_4_mask = 1'h1;
  assign rob_rd_addr_MPORT_4_en = reset;
  assign rob_rd_addr_MPORT_5_data = 5'h0;
  assign rob_rd_addr_MPORT_5_addr = 4'h1;
  assign rob_rd_addr_MPORT_5_mask = 1'h1;
  assign rob_rd_addr_MPORT_5_en = reset;
  assign rob_rd_addr_MPORT_6_data = 5'h0;
  assign rob_rd_addr_MPORT_6_addr = 4'h2;
  assign rob_rd_addr_MPORT_6_mask = 1'h1;
  assign rob_rd_addr_MPORT_6_en = reset;
  assign rob_rd_addr_MPORT_7_data = 5'h0;
  assign rob_rd_addr_MPORT_7_addr = 4'h3;
  assign rob_rd_addr_MPORT_7_mask = 1'h1;
  assign rob_rd_addr_MPORT_7_en = reset;
  assign rob_rd_addr_MPORT_8_data = 5'h0;
  assign rob_rd_addr_MPORT_8_addr = 4'h4;
  assign rob_rd_addr_MPORT_8_mask = 1'h1;
  assign rob_rd_addr_MPORT_8_en = reset;
  assign rob_rd_addr_MPORT_9_data = 5'h0;
  assign rob_rd_addr_MPORT_9_addr = 4'h5;
  assign rob_rd_addr_MPORT_9_mask = 1'h1;
  assign rob_rd_addr_MPORT_9_en = reset;
  assign rob_rd_addr_MPORT_10_data = 5'h0;
  assign rob_rd_addr_MPORT_10_addr = 4'h6;
  assign rob_rd_addr_MPORT_10_mask = 1'h1;
  assign rob_rd_addr_MPORT_10_en = reset;
  assign rob_rd_addr_MPORT_11_data = 5'h0;
  assign rob_rd_addr_MPORT_11_addr = 4'h7;
  assign rob_rd_addr_MPORT_11_mask = 1'h1;
  assign rob_rd_addr_MPORT_11_en = reset;
  assign rob_rd_addr_MPORT_12_data = 5'h0;
  assign rob_rd_addr_MPORT_12_addr = 4'h8;
  assign rob_rd_addr_MPORT_12_mask = 1'h1;
  assign rob_rd_addr_MPORT_12_en = reset;
  assign rob_rd_addr_MPORT_13_data = 5'h0;
  assign rob_rd_addr_MPORT_13_addr = 4'h9;
  assign rob_rd_addr_MPORT_13_mask = 1'h1;
  assign rob_rd_addr_MPORT_13_en = reset;
  assign rob_rd_addr_MPORT_14_data = 5'h0;
  assign rob_rd_addr_MPORT_14_addr = 4'ha;
  assign rob_rd_addr_MPORT_14_mask = 1'h1;
  assign rob_rd_addr_MPORT_14_en = reset;
  assign rob_rd_addr_MPORT_15_data = 5'h0;
  assign rob_rd_addr_MPORT_15_addr = 4'hb;
  assign rob_rd_addr_MPORT_15_mask = 1'h1;
  assign rob_rd_addr_MPORT_15_en = reset;
  assign rob_rd_addr_MPORT_16_data = 5'h0;
  assign rob_rd_addr_MPORT_16_addr = 4'hc;
  assign rob_rd_addr_MPORT_16_mask = 1'h1;
  assign rob_rd_addr_MPORT_16_en = reset;
  assign rob_rd_addr_MPORT_17_data = 5'h0;
  assign rob_rd_addr_MPORT_17_addr = 4'hd;
  assign rob_rd_addr_MPORT_17_mask = 1'h1;
  assign rob_rd_addr_MPORT_17_en = reset;
  assign rob_rd_addr_MPORT_18_data = 5'h0;
  assign rob_rd_addr_MPORT_18_addr = 4'he;
  assign rob_rd_addr_MPORT_18_mask = 1'h1;
  assign rob_rd_addr_MPORT_18_en = reset;
  assign rob_rd_addr_MPORT_19_data = 5'h0;
  assign rob_rd_addr_MPORT_19_addr = 4'hf;
  assign rob_rd_addr_MPORT_19_mask = 1'h1;
  assign rob_rd_addr_MPORT_19_en = reset;
//   assign rob_rd_en_MPORT_2_en = rob_rd_en_MPORT_2_en_pipe_0;
  assign rob_rd_en_MPORT_2_addr = rob_rd_en_MPORT_2_addr_pipe_0;
  assign rob_rd_en_MPORT_2_data = rob_rd_en[rob_rd_en_MPORT_2_addr]; // @[Rob.scala 44:24]
//   assign rob_rd_en_MPORT_3_en = rob_rd_en_MPORT_3_en_pipe_0;
  assign rob_rd_en_MPORT_3_addr = rob_rd_en_MPORT_3_addr_pipe_0;
  assign rob_rd_en_MPORT_3_data = rob_rd_en[rob_rd_en_MPORT_3_addr]; // @[Rob.scala 44:24]
  assign rob_rd_en_MPORT_data = io_in_bits_vec_0_rd_en;
  assign rob_rd_en_MPORT_addr = enq_vec_0[3:0];
  assign rob_rd_en_MPORT_mask = 1'h1;
  assign rob_rd_en_MPORT_en = _T_20 & _T_21;
  assign rob_rd_en_MPORT_1_data = io_in_bits_vec_1_rd_en;
  assign rob_rd_en_MPORT_1_addr = _GEN_289[3:0];
  assign rob_rd_en_MPORT_1_mask = 1'h1;
  assign rob_rd_en_MPORT_1_en = _T_25 & _T_21;
  assign rob_rd_en_MPORT_4_data = 1'h0;
  assign rob_rd_en_MPORT_4_addr = 4'h0;
  assign rob_rd_en_MPORT_4_mask = 1'h1;
  assign rob_rd_en_MPORT_4_en = reset;
  assign rob_rd_en_MPORT_5_data = 1'h0;
  assign rob_rd_en_MPORT_5_addr = 4'h1;
  assign rob_rd_en_MPORT_5_mask = 1'h1;
  assign rob_rd_en_MPORT_5_en = reset;
  assign rob_rd_en_MPORT_6_data = 1'h0;
  assign rob_rd_en_MPORT_6_addr = 4'h2;
  assign rob_rd_en_MPORT_6_mask = 1'h1;
  assign rob_rd_en_MPORT_6_en = reset;
  assign rob_rd_en_MPORT_7_data = 1'h0;
  assign rob_rd_en_MPORT_7_addr = 4'h3;
  assign rob_rd_en_MPORT_7_mask = 1'h1;
  assign rob_rd_en_MPORT_7_en = reset;
  assign rob_rd_en_MPORT_8_data = 1'h0;
  assign rob_rd_en_MPORT_8_addr = 4'h4;
  assign rob_rd_en_MPORT_8_mask = 1'h1;
  assign rob_rd_en_MPORT_8_en = reset;
  assign rob_rd_en_MPORT_9_data = 1'h0;
  assign rob_rd_en_MPORT_9_addr = 4'h5;
  assign rob_rd_en_MPORT_9_mask = 1'h1;
  assign rob_rd_en_MPORT_9_en = reset;
  assign rob_rd_en_MPORT_10_data = 1'h0;
  assign rob_rd_en_MPORT_10_addr = 4'h6;
  assign rob_rd_en_MPORT_10_mask = 1'h1;
  assign rob_rd_en_MPORT_10_en = reset;
  assign rob_rd_en_MPORT_11_data = 1'h0;
  assign rob_rd_en_MPORT_11_addr = 4'h7;
  assign rob_rd_en_MPORT_11_mask = 1'h1;
  assign rob_rd_en_MPORT_11_en = reset;
  assign rob_rd_en_MPORT_12_data = 1'h0;
  assign rob_rd_en_MPORT_12_addr = 4'h8;
  assign rob_rd_en_MPORT_12_mask = 1'h1;
  assign rob_rd_en_MPORT_12_en = reset;
  assign rob_rd_en_MPORT_13_data = 1'h0;
  assign rob_rd_en_MPORT_13_addr = 4'h9;
  assign rob_rd_en_MPORT_13_mask = 1'h1;
  assign rob_rd_en_MPORT_13_en = reset;
  assign rob_rd_en_MPORT_14_data = 1'h0;
  assign rob_rd_en_MPORT_14_addr = 4'ha;
  assign rob_rd_en_MPORT_14_mask = 1'h1;
  assign rob_rd_en_MPORT_14_en = reset;
  assign rob_rd_en_MPORT_15_data = 1'h0;
  assign rob_rd_en_MPORT_15_addr = 4'hb;
  assign rob_rd_en_MPORT_15_mask = 1'h1;
  assign rob_rd_en_MPORT_15_en = reset;
  assign rob_rd_en_MPORT_16_data = 1'h0;
  assign rob_rd_en_MPORT_16_addr = 4'hc;
  assign rob_rd_en_MPORT_16_mask = 1'h1;
  assign rob_rd_en_MPORT_16_en = reset;
  assign rob_rd_en_MPORT_17_data = 1'h0;
  assign rob_rd_en_MPORT_17_addr = 4'hd;
  assign rob_rd_en_MPORT_17_mask = 1'h1;
  assign rob_rd_en_MPORT_17_en = reset;
  assign rob_rd_en_MPORT_18_data = 1'h0;
  assign rob_rd_en_MPORT_18_addr = 4'he;
  assign rob_rd_en_MPORT_18_mask = 1'h1;
  assign rob_rd_en_MPORT_18_en = reset;
  assign rob_rd_en_MPORT_19_data = 1'h0;
  assign rob_rd_en_MPORT_19_addr = 4'hf;
  assign rob_rd_en_MPORT_19_mask = 1'h1;
  assign rob_rd_en_MPORT_19_en = reset;
//   assign rob_rd_paddr_MPORT_2_en = rob_rd_paddr_MPORT_2_en_pipe_0;
  assign rob_rd_paddr_MPORT_2_addr = rob_rd_paddr_MPORT_2_addr_pipe_0;
  assign rob_rd_paddr_MPORT_2_data = rob_rd_paddr[rob_rd_paddr_MPORT_2_addr]; // @[Rob.scala 44:24]
//   assign rob_rd_paddr_MPORT_3_en = rob_rd_paddr_MPORT_3_en_pipe_0;
  assign rob_rd_paddr_MPORT_3_addr = rob_rd_paddr_MPORT_3_addr_pipe_0;
  assign rob_rd_paddr_MPORT_3_data = rob_rd_paddr[rob_rd_paddr_MPORT_3_addr]; // @[Rob.scala 44:24]
  assign rob_rd_paddr_MPORT_data = io_in_bits_vec_0_rd_paddr;
  assign rob_rd_paddr_MPORT_addr = enq_vec_0[3:0];
  assign rob_rd_paddr_MPORT_mask = 1'h1;
  assign rob_rd_paddr_MPORT_en = _T_20 & _T_21;
  assign rob_rd_paddr_MPORT_1_data = io_in_bits_vec_1_rd_paddr;
  assign rob_rd_paddr_MPORT_1_addr = _GEN_289[3:0];
  assign rob_rd_paddr_MPORT_1_mask = 1'h1;
  assign rob_rd_paddr_MPORT_1_en = _T_25 & _T_21;
  assign rob_rd_paddr_MPORT_4_data = 6'h0;
  assign rob_rd_paddr_MPORT_4_addr = 4'h0;
  assign rob_rd_paddr_MPORT_4_mask = 1'h1;
  assign rob_rd_paddr_MPORT_4_en = reset;
  assign rob_rd_paddr_MPORT_5_data = 6'h0;
  assign rob_rd_paddr_MPORT_5_addr = 4'h1;
  assign rob_rd_paddr_MPORT_5_mask = 1'h1;
  assign rob_rd_paddr_MPORT_5_en = reset;
  assign rob_rd_paddr_MPORT_6_data = 6'h0;
  assign rob_rd_paddr_MPORT_6_addr = 4'h2;
  assign rob_rd_paddr_MPORT_6_mask = 1'h1;
  assign rob_rd_paddr_MPORT_6_en = reset;
  assign rob_rd_paddr_MPORT_7_data = 6'h0;
  assign rob_rd_paddr_MPORT_7_addr = 4'h3;
  assign rob_rd_paddr_MPORT_7_mask = 1'h1;
  assign rob_rd_paddr_MPORT_7_en = reset;
  assign rob_rd_paddr_MPORT_8_data = 6'h0;
  assign rob_rd_paddr_MPORT_8_addr = 4'h4;
  assign rob_rd_paddr_MPORT_8_mask = 1'h1;
  assign rob_rd_paddr_MPORT_8_en = reset;
  assign rob_rd_paddr_MPORT_9_data = 6'h0;
  assign rob_rd_paddr_MPORT_9_addr = 4'h5;
  assign rob_rd_paddr_MPORT_9_mask = 1'h1;
  assign rob_rd_paddr_MPORT_9_en = reset;
  assign rob_rd_paddr_MPORT_10_data = 6'h0;
  assign rob_rd_paddr_MPORT_10_addr = 4'h6;
  assign rob_rd_paddr_MPORT_10_mask = 1'h1;
  assign rob_rd_paddr_MPORT_10_en = reset;
  assign rob_rd_paddr_MPORT_11_data = 6'h0;
  assign rob_rd_paddr_MPORT_11_addr = 4'h7;
  assign rob_rd_paddr_MPORT_11_mask = 1'h1;
  assign rob_rd_paddr_MPORT_11_en = reset;
  assign rob_rd_paddr_MPORT_12_data = 6'h0;
  assign rob_rd_paddr_MPORT_12_addr = 4'h8;
  assign rob_rd_paddr_MPORT_12_mask = 1'h1;
  assign rob_rd_paddr_MPORT_12_en = reset;
  assign rob_rd_paddr_MPORT_13_data = 6'h0;
  assign rob_rd_paddr_MPORT_13_addr = 4'h9;
  assign rob_rd_paddr_MPORT_13_mask = 1'h1;
  assign rob_rd_paddr_MPORT_13_en = reset;
  assign rob_rd_paddr_MPORT_14_data = 6'h0;
  assign rob_rd_paddr_MPORT_14_addr = 4'ha;
  assign rob_rd_paddr_MPORT_14_mask = 1'h1;
  assign rob_rd_paddr_MPORT_14_en = reset;
  assign rob_rd_paddr_MPORT_15_data = 6'h0;
  assign rob_rd_paddr_MPORT_15_addr = 4'hb;
  assign rob_rd_paddr_MPORT_15_mask = 1'h1;
  assign rob_rd_paddr_MPORT_15_en = reset;
  assign rob_rd_paddr_MPORT_16_data = 6'h0;
  assign rob_rd_paddr_MPORT_16_addr = 4'hc;
  assign rob_rd_paddr_MPORT_16_mask = 1'h1;
  assign rob_rd_paddr_MPORT_16_en = reset;
  assign rob_rd_paddr_MPORT_17_data = 6'h0;
  assign rob_rd_paddr_MPORT_17_addr = 4'hd;
  assign rob_rd_paddr_MPORT_17_mask = 1'h1;
  assign rob_rd_paddr_MPORT_17_en = reset;
  assign rob_rd_paddr_MPORT_18_data = 6'h0;
  assign rob_rd_paddr_MPORT_18_addr = 4'he;
  assign rob_rd_paddr_MPORT_18_mask = 1'h1;
  assign rob_rd_paddr_MPORT_18_en = reset;
  assign rob_rd_paddr_MPORT_19_data = 6'h0;
  assign rob_rd_paddr_MPORT_19_addr = 4'hf;
  assign rob_rd_paddr_MPORT_19_mask = 1'h1;
  assign rob_rd_paddr_MPORT_19_en = reset;
//   assign rob_rd_ppaddr_MPORT_2_en = rob_rd_ppaddr_MPORT_2_en_pipe_0;
  assign rob_rd_ppaddr_MPORT_2_addr = rob_rd_ppaddr_MPORT_2_addr_pipe_0;
  assign rob_rd_ppaddr_MPORT_2_data = rob_rd_ppaddr[rob_rd_ppaddr_MPORT_2_addr]; // @[Rob.scala 44:24]
//   assign rob_rd_ppaddr_MPORT_3_en = rob_rd_ppaddr_MPORT_3_en_pipe_0;
  assign rob_rd_ppaddr_MPORT_3_addr = rob_rd_ppaddr_MPORT_3_addr_pipe_0;
  assign rob_rd_ppaddr_MPORT_3_data = rob_rd_ppaddr[rob_rd_ppaddr_MPORT_3_addr]; // @[Rob.scala 44:24]
  assign rob_rd_ppaddr_MPORT_data = io_in_bits_vec_0_rd_ppaddr;
  assign rob_rd_ppaddr_MPORT_addr = enq_vec_0[3:0];
  assign rob_rd_ppaddr_MPORT_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_en = _T_20 & _T_21;
  assign rob_rd_ppaddr_MPORT_1_data = io_in_bits_vec_1_rd_ppaddr;
  assign rob_rd_ppaddr_MPORT_1_addr = _GEN_289[3:0];
  assign rob_rd_ppaddr_MPORT_1_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_1_en = _T_25 & _T_21;
  assign rob_rd_ppaddr_MPORT_4_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_4_addr = 4'h0;
  assign rob_rd_ppaddr_MPORT_4_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_4_en = reset;
  assign rob_rd_ppaddr_MPORT_5_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_5_addr = 4'h1;
  assign rob_rd_ppaddr_MPORT_5_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_5_en = reset;
  assign rob_rd_ppaddr_MPORT_6_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_6_addr = 4'h2;
  assign rob_rd_ppaddr_MPORT_6_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_6_en = reset;
  assign rob_rd_ppaddr_MPORT_7_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_7_addr = 4'h3;
  assign rob_rd_ppaddr_MPORT_7_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_7_en = reset;
  assign rob_rd_ppaddr_MPORT_8_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_8_addr = 4'h4;
  assign rob_rd_ppaddr_MPORT_8_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_8_en = reset;
  assign rob_rd_ppaddr_MPORT_9_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_9_addr = 4'h5;
  assign rob_rd_ppaddr_MPORT_9_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_9_en = reset;
  assign rob_rd_ppaddr_MPORT_10_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_10_addr = 4'h6;
  assign rob_rd_ppaddr_MPORT_10_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_10_en = reset;
  assign rob_rd_ppaddr_MPORT_11_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_11_addr = 4'h7;
  assign rob_rd_ppaddr_MPORT_11_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_11_en = reset;
  assign rob_rd_ppaddr_MPORT_12_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_12_addr = 4'h8;
  assign rob_rd_ppaddr_MPORT_12_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_12_en = reset;
  assign rob_rd_ppaddr_MPORT_13_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_13_addr = 4'h9;
  assign rob_rd_ppaddr_MPORT_13_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_13_en = reset;
  assign rob_rd_ppaddr_MPORT_14_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_14_addr = 4'ha;
  assign rob_rd_ppaddr_MPORT_14_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_14_en = reset;
  assign rob_rd_ppaddr_MPORT_15_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_15_addr = 4'hb;
  assign rob_rd_ppaddr_MPORT_15_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_15_en = reset;
  assign rob_rd_ppaddr_MPORT_16_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_16_addr = 4'hc;
  assign rob_rd_ppaddr_MPORT_16_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_16_en = reset;
  assign rob_rd_ppaddr_MPORT_17_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_17_addr = 4'hd;
  assign rob_rd_ppaddr_MPORT_17_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_17_en = reset;
  assign rob_rd_ppaddr_MPORT_18_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_18_addr = 4'he;
  assign rob_rd_ppaddr_MPORT_18_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_18_en = reset;
  assign rob_rd_ppaddr_MPORT_19_data = 6'h0;
  assign rob_rd_ppaddr_MPORT_19_addr = 4'hf;
  assign rob_rd_ppaddr_MPORT_19_mask = 1'h1;
  assign rob_rd_ppaddr_MPORT_19_en = reset;
  assign io_in_ready = enq_ready; // @[Rob.scala 107:15]
  assign io_rob_addr_0 = io_in_bits_vec_0_valid & _T_11 & ~io_flush ? enq_ptr : 4'h0; // @[Rob.scala 91:65 95:22 97:22]
  assign io_rob_addr_1 = io_in_bits_vec_1_valid & _T_11 & ~io_flush ? _GEN_289[3:0] : 4'h0; // @[Rob.scala 91:65 95:22 97:22]
  assign io_cm_0_valid = cm_0_valid & ~intr; // @[Rob.scala 352:35]
  assign io_cm_0_rd_addr = rob_rd_addr_MPORT_2_data; // @[Rob.scala 156:21 229:16]
  assign io_cm_0_rd_en = rob_rd_en_MPORT_2_data; // @[Rob.scala 156:21 229:16]
  assign io_cm_0_rd_paddr = rob_rd_paddr_MPORT_2_data; // @[Rob.scala 156:21 229:16]
  assign io_cm_0_rd_ppaddr = rob_rd_ppaddr_MPORT_2_data; // @[Rob.scala 156:21 229:16]
  assign io_cm_1_valid = cm_1_valid & ~intr; // @[Rob.scala 352:35]
  assign io_cm_1_rd_addr = rob_rd_addr_MPORT_3_data; // @[Rob.scala 156:21 229:16]
  assign io_cm_1_rd_en = rob_rd_en_MPORT_3_data; // @[Rob.scala 156:21 229:16]
  assign io_cm_1_rd_paddr = rob_rd_paddr_MPORT_3_data; // @[Rob.scala 156:21 229:16]
  assign io_cm_1_rd_ppaddr = rob_rd_ppaddr_MPORT_3_data; // @[Rob.scala 156:21 229:16]
  assign io_jmp_packet_valid = intr | _GEN_1654; // @[Rob.scala 311:15 312:27]
  assign io_jmp_packet_inst_pc = intr ? intr_mepc[31:0] : _GEN_1655; // @[Rob.scala 311:15 313:27]
  assign io_jmp_packet_jmp = intr | _GEN_1656; // @[Rob.scala 311:15 314:27]
  assign io_jmp_packet_jmp_pc = intr ? intr_jmp_pc : _GEN_1657; // @[Rob.scala 311:15 315:27]
  assign io_jmp_packet_mis = intr | _GEN_1658; // @[Rob.scala 311:15 316:27]
  assign io_jmp_packet_sys = intr | _GEN_1659; // @[Rob.scala 311:15 317:27]
  assign io_sq_deq_req = sq_deq_req & _T_142; // @[Rob.scala 356:31]
  assign io_sys_ready = deq_uop_0_fu_code == 3'h3 & _T_53 & ~rob_empty; // @[Rob.scala 233:68]
  assign intr_mcause_0 = intr_mcause;
  assign intr_mstatus_0 = intr_mstatus;
  assign intr_0 = intr;
  assign intr_mepc_0 = intr_mepc;
  always @(posedge clock) begin
    if (rob_pc_MPORT_en & rob_pc_MPORT_mask) begin
      rob_pc[rob_pc_MPORT_addr] <= rob_pc_MPORT_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_1_en & rob_pc_MPORT_1_mask) begin
      rob_pc[rob_pc_MPORT_1_addr] <= rob_pc_MPORT_1_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_4_en & rob_pc_MPORT_4_mask) begin
      rob_pc[rob_pc_MPORT_4_addr] <= rob_pc_MPORT_4_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_5_en & rob_pc_MPORT_5_mask) begin
      rob_pc[rob_pc_MPORT_5_addr] <= rob_pc_MPORT_5_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_6_en & rob_pc_MPORT_6_mask) begin
      rob_pc[rob_pc_MPORT_6_addr] <= rob_pc_MPORT_6_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_7_en & rob_pc_MPORT_7_mask) begin
      rob_pc[rob_pc_MPORT_7_addr] <= rob_pc_MPORT_7_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_8_en & rob_pc_MPORT_8_mask) begin
      rob_pc[rob_pc_MPORT_8_addr] <= rob_pc_MPORT_8_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_9_en & rob_pc_MPORT_9_mask) begin
      rob_pc[rob_pc_MPORT_9_addr] <= rob_pc_MPORT_9_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_10_en & rob_pc_MPORT_10_mask) begin
      rob_pc[rob_pc_MPORT_10_addr] <= rob_pc_MPORT_10_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_11_en & rob_pc_MPORT_11_mask) begin
      rob_pc[rob_pc_MPORT_11_addr] <= rob_pc_MPORT_11_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_12_en & rob_pc_MPORT_12_mask) begin
      rob_pc[rob_pc_MPORT_12_addr] <= rob_pc_MPORT_12_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_13_en & rob_pc_MPORT_13_mask) begin
      rob_pc[rob_pc_MPORT_13_addr] <= rob_pc_MPORT_13_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_14_en & rob_pc_MPORT_14_mask) begin
      rob_pc[rob_pc_MPORT_14_addr] <= rob_pc_MPORT_14_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_15_en & rob_pc_MPORT_15_mask) begin
      rob_pc[rob_pc_MPORT_15_addr] <= rob_pc_MPORT_15_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_16_en & rob_pc_MPORT_16_mask) begin
      rob_pc[rob_pc_MPORT_16_addr] <= rob_pc_MPORT_16_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_17_en & rob_pc_MPORT_17_mask) begin
      rob_pc[rob_pc_MPORT_17_addr] <= rob_pc_MPORT_17_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_18_en & rob_pc_MPORT_18_mask) begin
      rob_pc[rob_pc_MPORT_18_addr] <= rob_pc_MPORT_18_data; // @[Rob.scala 44:24]
    end
    if (rob_pc_MPORT_19_en & rob_pc_MPORT_19_mask) begin
      rob_pc[rob_pc_MPORT_19_addr] <= rob_pc_MPORT_19_data; // @[Rob.scala 44:24]
    end
//     rob_pc_MPORT_2_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      rob_pc_MPORT_2_addr_pipe_0 <= next_deq_vec_0[3:0];
    end
//     rob_pc_MPORT_3_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      rob_pc_MPORT_3_addr_pipe_0 <= next_deq_vec_1[3:0];
    end
    if (rob_fu_code_MPORT_en & rob_fu_code_MPORT_mask) begin
      rob_fu_code[rob_fu_code_MPORT_addr] <= rob_fu_code_MPORT_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_1_en & rob_fu_code_MPORT_1_mask) begin
      rob_fu_code[rob_fu_code_MPORT_1_addr] <= rob_fu_code_MPORT_1_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_4_en & rob_fu_code_MPORT_4_mask) begin
      rob_fu_code[rob_fu_code_MPORT_4_addr] <= rob_fu_code_MPORT_4_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_5_en & rob_fu_code_MPORT_5_mask) begin
      rob_fu_code[rob_fu_code_MPORT_5_addr] <= rob_fu_code_MPORT_5_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_6_en & rob_fu_code_MPORT_6_mask) begin
      rob_fu_code[rob_fu_code_MPORT_6_addr] <= rob_fu_code_MPORT_6_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_7_en & rob_fu_code_MPORT_7_mask) begin
      rob_fu_code[rob_fu_code_MPORT_7_addr] <= rob_fu_code_MPORT_7_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_8_en & rob_fu_code_MPORT_8_mask) begin
      rob_fu_code[rob_fu_code_MPORT_8_addr] <= rob_fu_code_MPORT_8_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_9_en & rob_fu_code_MPORT_9_mask) begin
      rob_fu_code[rob_fu_code_MPORT_9_addr] <= rob_fu_code_MPORT_9_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_10_en & rob_fu_code_MPORT_10_mask) begin
      rob_fu_code[rob_fu_code_MPORT_10_addr] <= rob_fu_code_MPORT_10_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_11_en & rob_fu_code_MPORT_11_mask) begin
      rob_fu_code[rob_fu_code_MPORT_11_addr] <= rob_fu_code_MPORT_11_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_12_en & rob_fu_code_MPORT_12_mask) begin
      rob_fu_code[rob_fu_code_MPORT_12_addr] <= rob_fu_code_MPORT_12_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_13_en & rob_fu_code_MPORT_13_mask) begin
      rob_fu_code[rob_fu_code_MPORT_13_addr] <= rob_fu_code_MPORT_13_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_14_en & rob_fu_code_MPORT_14_mask) begin
      rob_fu_code[rob_fu_code_MPORT_14_addr] <= rob_fu_code_MPORT_14_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_15_en & rob_fu_code_MPORT_15_mask) begin
      rob_fu_code[rob_fu_code_MPORT_15_addr] <= rob_fu_code_MPORT_15_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_16_en & rob_fu_code_MPORT_16_mask) begin
      rob_fu_code[rob_fu_code_MPORT_16_addr] <= rob_fu_code_MPORT_16_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_17_en & rob_fu_code_MPORT_17_mask) begin
      rob_fu_code[rob_fu_code_MPORT_17_addr] <= rob_fu_code_MPORT_17_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_18_en & rob_fu_code_MPORT_18_mask) begin
      rob_fu_code[rob_fu_code_MPORT_18_addr] <= rob_fu_code_MPORT_18_data; // @[Rob.scala 44:24]
    end
    if (rob_fu_code_MPORT_19_en & rob_fu_code_MPORT_19_mask) begin
      rob_fu_code[rob_fu_code_MPORT_19_addr] <= rob_fu_code_MPORT_19_data; // @[Rob.scala 44:24]
    end
//     rob_fu_code_MPORT_2_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      rob_fu_code_MPORT_2_addr_pipe_0 <= next_deq_vec_0[3:0];
    end
//     rob_fu_code_MPORT_3_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      rob_fu_code_MPORT_3_addr_pipe_0 <= next_deq_vec_1[3:0];
    end
    if (rob_sys_code_MPORT_en & rob_sys_code_MPORT_mask) begin
      rob_sys_code[rob_sys_code_MPORT_addr] <= rob_sys_code_MPORT_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_1_en & rob_sys_code_MPORT_1_mask) begin
      rob_sys_code[rob_sys_code_MPORT_1_addr] <= rob_sys_code_MPORT_1_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_4_en & rob_sys_code_MPORT_4_mask) begin
      rob_sys_code[rob_sys_code_MPORT_4_addr] <= rob_sys_code_MPORT_4_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_5_en & rob_sys_code_MPORT_5_mask) begin
      rob_sys_code[rob_sys_code_MPORT_5_addr] <= rob_sys_code_MPORT_5_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_6_en & rob_sys_code_MPORT_6_mask) begin
      rob_sys_code[rob_sys_code_MPORT_6_addr] <= rob_sys_code_MPORT_6_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_7_en & rob_sys_code_MPORT_7_mask) begin
      rob_sys_code[rob_sys_code_MPORT_7_addr] <= rob_sys_code_MPORT_7_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_8_en & rob_sys_code_MPORT_8_mask) begin
      rob_sys_code[rob_sys_code_MPORT_8_addr] <= rob_sys_code_MPORT_8_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_9_en & rob_sys_code_MPORT_9_mask) begin
      rob_sys_code[rob_sys_code_MPORT_9_addr] <= rob_sys_code_MPORT_9_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_10_en & rob_sys_code_MPORT_10_mask) begin
      rob_sys_code[rob_sys_code_MPORT_10_addr] <= rob_sys_code_MPORT_10_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_11_en & rob_sys_code_MPORT_11_mask) begin
      rob_sys_code[rob_sys_code_MPORT_11_addr] <= rob_sys_code_MPORT_11_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_12_en & rob_sys_code_MPORT_12_mask) begin
      rob_sys_code[rob_sys_code_MPORT_12_addr] <= rob_sys_code_MPORT_12_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_13_en & rob_sys_code_MPORT_13_mask) begin
      rob_sys_code[rob_sys_code_MPORT_13_addr] <= rob_sys_code_MPORT_13_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_14_en & rob_sys_code_MPORT_14_mask) begin
      rob_sys_code[rob_sys_code_MPORT_14_addr] <= rob_sys_code_MPORT_14_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_15_en & rob_sys_code_MPORT_15_mask) begin
      rob_sys_code[rob_sys_code_MPORT_15_addr] <= rob_sys_code_MPORT_15_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_16_en & rob_sys_code_MPORT_16_mask) begin
      rob_sys_code[rob_sys_code_MPORT_16_addr] <= rob_sys_code_MPORT_16_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_17_en & rob_sys_code_MPORT_17_mask) begin
      rob_sys_code[rob_sys_code_MPORT_17_addr] <= rob_sys_code_MPORT_17_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_18_en & rob_sys_code_MPORT_18_mask) begin
      rob_sys_code[rob_sys_code_MPORT_18_addr] <= rob_sys_code_MPORT_18_data; // @[Rob.scala 44:24]
    end
    if (rob_sys_code_MPORT_19_en & rob_sys_code_MPORT_19_mask) begin
      rob_sys_code[rob_sys_code_MPORT_19_addr] <= rob_sys_code_MPORT_19_data; // @[Rob.scala 44:24]
    end
//     rob_sys_code_MPORT_2_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      rob_sys_code_MPORT_2_addr_pipe_0 <= next_deq_vec_0[3:0];
    end
//     rob_sys_code_MPORT_3_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      rob_sys_code_MPORT_3_addr_pipe_0 <= next_deq_vec_1[3:0];
    end
    if (rob_rd_addr_MPORT_en & rob_rd_addr_MPORT_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_addr] <= rob_rd_addr_MPORT_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_1_en & rob_rd_addr_MPORT_1_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_1_addr] <= rob_rd_addr_MPORT_1_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_4_en & rob_rd_addr_MPORT_4_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_4_addr] <= rob_rd_addr_MPORT_4_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_5_en & rob_rd_addr_MPORT_5_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_5_addr] <= rob_rd_addr_MPORT_5_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_6_en & rob_rd_addr_MPORT_6_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_6_addr] <= rob_rd_addr_MPORT_6_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_7_en & rob_rd_addr_MPORT_7_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_7_addr] <= rob_rd_addr_MPORT_7_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_8_en & rob_rd_addr_MPORT_8_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_8_addr] <= rob_rd_addr_MPORT_8_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_9_en & rob_rd_addr_MPORT_9_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_9_addr] <= rob_rd_addr_MPORT_9_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_10_en & rob_rd_addr_MPORT_10_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_10_addr] <= rob_rd_addr_MPORT_10_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_11_en & rob_rd_addr_MPORT_11_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_11_addr] <= rob_rd_addr_MPORT_11_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_12_en & rob_rd_addr_MPORT_12_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_12_addr] <= rob_rd_addr_MPORT_12_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_13_en & rob_rd_addr_MPORT_13_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_13_addr] <= rob_rd_addr_MPORT_13_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_14_en & rob_rd_addr_MPORT_14_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_14_addr] <= rob_rd_addr_MPORT_14_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_15_en & rob_rd_addr_MPORT_15_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_15_addr] <= rob_rd_addr_MPORT_15_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_16_en & rob_rd_addr_MPORT_16_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_16_addr] <= rob_rd_addr_MPORT_16_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_17_en & rob_rd_addr_MPORT_17_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_17_addr] <= rob_rd_addr_MPORT_17_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_18_en & rob_rd_addr_MPORT_18_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_18_addr] <= rob_rd_addr_MPORT_18_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_addr_MPORT_19_en & rob_rd_addr_MPORT_19_mask) begin
      rob_rd_addr[rob_rd_addr_MPORT_19_addr] <= rob_rd_addr_MPORT_19_data; // @[Rob.scala 44:24]
    end
//     rob_rd_addr_MPORT_2_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      rob_rd_addr_MPORT_2_addr_pipe_0 <= next_deq_vec_0[3:0];
    end
//     rob_rd_addr_MPORT_3_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      rob_rd_addr_MPORT_3_addr_pipe_0 <= next_deq_vec_1[3:0];
    end
    if (rob_rd_en_MPORT_en & rob_rd_en_MPORT_mask) begin
      rob_rd_en[rob_rd_en_MPORT_addr] <= rob_rd_en_MPORT_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_1_en & rob_rd_en_MPORT_1_mask) begin
      rob_rd_en[rob_rd_en_MPORT_1_addr] <= rob_rd_en_MPORT_1_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_4_en & rob_rd_en_MPORT_4_mask) begin
      rob_rd_en[rob_rd_en_MPORT_4_addr] <= rob_rd_en_MPORT_4_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_5_en & rob_rd_en_MPORT_5_mask) begin
      rob_rd_en[rob_rd_en_MPORT_5_addr] <= rob_rd_en_MPORT_5_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_6_en & rob_rd_en_MPORT_6_mask) begin
      rob_rd_en[rob_rd_en_MPORT_6_addr] <= rob_rd_en_MPORT_6_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_7_en & rob_rd_en_MPORT_7_mask) begin
      rob_rd_en[rob_rd_en_MPORT_7_addr] <= rob_rd_en_MPORT_7_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_8_en & rob_rd_en_MPORT_8_mask) begin
      rob_rd_en[rob_rd_en_MPORT_8_addr] <= rob_rd_en_MPORT_8_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_9_en & rob_rd_en_MPORT_9_mask) begin
      rob_rd_en[rob_rd_en_MPORT_9_addr] <= rob_rd_en_MPORT_9_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_10_en & rob_rd_en_MPORT_10_mask) begin
      rob_rd_en[rob_rd_en_MPORT_10_addr] <= rob_rd_en_MPORT_10_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_11_en & rob_rd_en_MPORT_11_mask) begin
      rob_rd_en[rob_rd_en_MPORT_11_addr] <= rob_rd_en_MPORT_11_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_12_en & rob_rd_en_MPORT_12_mask) begin
      rob_rd_en[rob_rd_en_MPORT_12_addr] <= rob_rd_en_MPORT_12_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_13_en & rob_rd_en_MPORT_13_mask) begin
      rob_rd_en[rob_rd_en_MPORT_13_addr] <= rob_rd_en_MPORT_13_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_14_en & rob_rd_en_MPORT_14_mask) begin
      rob_rd_en[rob_rd_en_MPORT_14_addr] <= rob_rd_en_MPORT_14_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_15_en & rob_rd_en_MPORT_15_mask) begin
      rob_rd_en[rob_rd_en_MPORT_15_addr] <= rob_rd_en_MPORT_15_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_16_en & rob_rd_en_MPORT_16_mask) begin
      rob_rd_en[rob_rd_en_MPORT_16_addr] <= rob_rd_en_MPORT_16_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_17_en & rob_rd_en_MPORT_17_mask) begin
      rob_rd_en[rob_rd_en_MPORT_17_addr] <= rob_rd_en_MPORT_17_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_18_en & rob_rd_en_MPORT_18_mask) begin
      rob_rd_en[rob_rd_en_MPORT_18_addr] <= rob_rd_en_MPORT_18_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_en_MPORT_19_en & rob_rd_en_MPORT_19_mask) begin
      rob_rd_en[rob_rd_en_MPORT_19_addr] <= rob_rd_en_MPORT_19_data; // @[Rob.scala 44:24]
    end
//     rob_rd_en_MPORT_2_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      rob_rd_en_MPORT_2_addr_pipe_0 <= next_deq_vec_0[3:0];
    end
//     rob_rd_en_MPORT_3_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      rob_rd_en_MPORT_3_addr_pipe_0 <= next_deq_vec_1[3:0];
    end
    if (rob_rd_paddr_MPORT_en & rob_rd_paddr_MPORT_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_addr] <= rob_rd_paddr_MPORT_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_1_en & rob_rd_paddr_MPORT_1_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_1_addr] <= rob_rd_paddr_MPORT_1_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_4_en & rob_rd_paddr_MPORT_4_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_4_addr] <= rob_rd_paddr_MPORT_4_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_5_en & rob_rd_paddr_MPORT_5_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_5_addr] <= rob_rd_paddr_MPORT_5_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_6_en & rob_rd_paddr_MPORT_6_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_6_addr] <= rob_rd_paddr_MPORT_6_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_7_en & rob_rd_paddr_MPORT_7_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_7_addr] <= rob_rd_paddr_MPORT_7_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_8_en & rob_rd_paddr_MPORT_8_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_8_addr] <= rob_rd_paddr_MPORT_8_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_9_en & rob_rd_paddr_MPORT_9_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_9_addr] <= rob_rd_paddr_MPORT_9_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_10_en & rob_rd_paddr_MPORT_10_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_10_addr] <= rob_rd_paddr_MPORT_10_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_11_en & rob_rd_paddr_MPORT_11_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_11_addr] <= rob_rd_paddr_MPORT_11_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_12_en & rob_rd_paddr_MPORT_12_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_12_addr] <= rob_rd_paddr_MPORT_12_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_13_en & rob_rd_paddr_MPORT_13_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_13_addr] <= rob_rd_paddr_MPORT_13_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_14_en & rob_rd_paddr_MPORT_14_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_14_addr] <= rob_rd_paddr_MPORT_14_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_15_en & rob_rd_paddr_MPORT_15_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_15_addr] <= rob_rd_paddr_MPORT_15_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_16_en & rob_rd_paddr_MPORT_16_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_16_addr] <= rob_rd_paddr_MPORT_16_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_17_en & rob_rd_paddr_MPORT_17_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_17_addr] <= rob_rd_paddr_MPORT_17_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_18_en & rob_rd_paddr_MPORT_18_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_18_addr] <= rob_rd_paddr_MPORT_18_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_paddr_MPORT_19_en & rob_rd_paddr_MPORT_19_mask) begin
      rob_rd_paddr[rob_rd_paddr_MPORT_19_addr] <= rob_rd_paddr_MPORT_19_data; // @[Rob.scala 44:24]
    end
//     rob_rd_paddr_MPORT_2_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      rob_rd_paddr_MPORT_2_addr_pipe_0 <= next_deq_vec_0[3:0];
    end
//     rob_rd_paddr_MPORT_3_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      rob_rd_paddr_MPORT_3_addr_pipe_0 <= next_deq_vec_1[3:0];
    end
    if (rob_rd_ppaddr_MPORT_en & rob_rd_ppaddr_MPORT_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_addr] <= rob_rd_ppaddr_MPORT_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_1_en & rob_rd_ppaddr_MPORT_1_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_1_addr] <= rob_rd_ppaddr_MPORT_1_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_4_en & rob_rd_ppaddr_MPORT_4_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_4_addr] <= rob_rd_ppaddr_MPORT_4_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_5_en & rob_rd_ppaddr_MPORT_5_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_5_addr] <= rob_rd_ppaddr_MPORT_5_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_6_en & rob_rd_ppaddr_MPORT_6_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_6_addr] <= rob_rd_ppaddr_MPORT_6_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_7_en & rob_rd_ppaddr_MPORT_7_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_7_addr] <= rob_rd_ppaddr_MPORT_7_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_8_en & rob_rd_ppaddr_MPORT_8_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_8_addr] <= rob_rd_ppaddr_MPORT_8_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_9_en & rob_rd_ppaddr_MPORT_9_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_9_addr] <= rob_rd_ppaddr_MPORT_9_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_10_en & rob_rd_ppaddr_MPORT_10_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_10_addr] <= rob_rd_ppaddr_MPORT_10_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_11_en & rob_rd_ppaddr_MPORT_11_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_11_addr] <= rob_rd_ppaddr_MPORT_11_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_12_en & rob_rd_ppaddr_MPORT_12_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_12_addr] <= rob_rd_ppaddr_MPORT_12_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_13_en & rob_rd_ppaddr_MPORT_13_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_13_addr] <= rob_rd_ppaddr_MPORT_13_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_14_en & rob_rd_ppaddr_MPORT_14_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_14_addr] <= rob_rd_ppaddr_MPORT_14_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_15_en & rob_rd_ppaddr_MPORT_15_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_15_addr] <= rob_rd_ppaddr_MPORT_15_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_16_en & rob_rd_ppaddr_MPORT_16_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_16_addr] <= rob_rd_ppaddr_MPORT_16_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_17_en & rob_rd_ppaddr_MPORT_17_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_17_addr] <= rob_rd_ppaddr_MPORT_17_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_18_en & rob_rd_ppaddr_MPORT_18_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_18_addr] <= rob_rd_ppaddr_MPORT_18_data; // @[Rob.scala 44:24]
    end
    if (rob_rd_ppaddr_MPORT_19_en & rob_rd_ppaddr_MPORT_19_mask) begin
      rob_rd_ppaddr[rob_rd_ppaddr_MPORT_19_addr] <= rob_rd_ppaddr_MPORT_19_data; // @[Rob.scala 44:24]
    end
//     rob_rd_ppaddr_MPORT_2_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      rob_rd_ppaddr_MPORT_2_addr_pipe_0 <= next_deq_vec_0[3:0];
    end
//     rob_rd_ppaddr_MPORT_3_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      rob_rd_ppaddr_MPORT_3_addr_pipe_0 <= next_deq_vec_1[3:0];
    end
    if (reset) begin // @[Rob.scala 46:24]
      enq_vec_0 <= 5'h0; // @[Rob.scala 46:24]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      enq_vec_0 <= 5'h0; // @[Rob.scala 336:13]
    end else if (_T_11 & _T_21) begin // @[Rob.scala 103:36]
      enq_vec_0 <= next_enq_vec_0; // @[Rob.scala 104:13]
    end
    if (reset) begin // @[Rob.scala 46:24]
      enq_vec_1 <= 5'h1; // @[Rob.scala 46:24]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      enq_vec_1 <= 5'h1; // @[Rob.scala 336:13]
    end else if (_T_11 & _T_21) begin // @[Rob.scala 103:36]
      enq_vec_1 <= next_enq_vec_1; // @[Rob.scala 104:13]
    end
    if (reset) begin // @[Rob.scala 47:24]
      deq_vec_0 <= 5'h0; // @[Rob.scala 47:24]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      deq_vec_0 <= 5'h0; // @[Rob.scala 337:13]
    end else begin
      deq_vec_0 <= next_deq_vec_0; // @[Rob.scala 123:11]
    end
    if (reset) begin // @[Rob.scala 47:24]
      deq_vec_1 <= 5'h1; // @[Rob.scala 47:24]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      deq_vec_1 <= 5'h1; // @[Rob.scala 337:13]
    end else begin
      deq_vec_1 <= next_deq_vec_1; // @[Rob.scala 123:11]
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_15 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_15 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_15 <= _GEN_1105;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_15 <= _GEN_849;
    end else begin
      complete_15 <= _GEN_721;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_14 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_14 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_14 <= _GEN_1104;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_14 <= _GEN_848;
    end else begin
      complete_14 <= _GEN_720;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_13 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_13 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_13 <= _GEN_1103;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_13 <= _GEN_847;
    end else begin
      complete_13 <= _GEN_719;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_12 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_12 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_12 <= _GEN_1102;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_12 <= _GEN_846;
    end else begin
      complete_12 <= _GEN_718;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_11 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_11 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_11 <= _GEN_1101;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_11 <= _GEN_845;
    end else begin
      complete_11 <= _GEN_717;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_10 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_10 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_10 <= _GEN_1100;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_10 <= _GEN_844;
    end else begin
      complete_10 <= _GEN_716;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_9 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_9 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_9 <= _GEN_1099;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_9 <= _GEN_843;
    end else begin
      complete_9 <= _GEN_715;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_8 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_8 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_8 <= _GEN_1098;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_8 <= _GEN_842;
    end else begin
      complete_8 <= _GEN_714;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_7 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_7 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_7 <= _GEN_1097;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_7 <= _GEN_841;
    end else begin
      complete_7 <= _GEN_713;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_6 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_6 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_6 <= _GEN_1096;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_6 <= _GEN_840;
    end else begin
      complete_6 <= _GEN_712;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_5 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_5 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_5 <= _GEN_1095;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_5 <= _GEN_839;
    end else begin
      complete_5 <= _GEN_711;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_4 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_4 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_4 <= _GEN_1094;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_4 <= _GEN_838;
    end else begin
      complete_4 <= _GEN_710;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_3 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_3 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_3 <= _GEN_1093;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_3 <= _GEN_837;
    end else begin
      complete_3 <= _GEN_709;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_2 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_2 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_2 <= _GEN_1092;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_2 <= _GEN_836;
    end else begin
      complete_2 <= _GEN_708;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_1 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_1 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_1 <= _GEN_1091;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_1 <= _GEN_835;
    end else begin
      complete_1 <= _GEN_707;
    end
    if (reset) begin // @[Rob.scala 70:25]
      complete_0 <= 1'h0; // @[Rob.scala 70:25]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      complete_0 <= 1'h0; // @[Rob.scala 334:14]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      complete_0 <= _GEN_1090;
    end else if (io_exe_1_valid) begin // @[Rob.scala 113:28]
      complete_0 <= _GEN_834;
    end else begin
      complete_0 <= _GEN_706;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_15_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_15_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hf == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_15_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_15_jmp_valid <= _GEN_1057;
      end
    end else begin
      ecp_15_jmp_valid <= _GEN_1057;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_14_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_14_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'he == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_14_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_14_jmp_valid <= _GEN_1056;
      end
    end else begin
      ecp_14_jmp_valid <= _GEN_1056;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_13_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_13_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hd == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_13_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_13_jmp_valid <= _GEN_1055;
      end
    end else begin
      ecp_13_jmp_valid <= _GEN_1055;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_12_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_12_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hc == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_12_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_12_jmp_valid <= _GEN_1054;
      end
    end else begin
      ecp_12_jmp_valid <= _GEN_1054;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_11_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_11_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hb == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_11_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_11_jmp_valid <= _GEN_1053;
      end
    end else begin
      ecp_11_jmp_valid <= _GEN_1053;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_10_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_10_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'ha == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_10_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_10_jmp_valid <= _GEN_1052;
      end
    end else begin
      ecp_10_jmp_valid <= _GEN_1052;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_9_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_9_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h9 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_9_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_9_jmp_valid <= _GEN_1051;
      end
    end else begin
      ecp_9_jmp_valid <= _GEN_1051;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_8_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_8_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h8 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_8_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_8_jmp_valid <= _GEN_1050;
      end
    end else begin
      ecp_8_jmp_valid <= _GEN_1050;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_7_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_7_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h7 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_7_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_7_jmp_valid <= _GEN_1049;
      end
    end else begin
      ecp_7_jmp_valid <= _GEN_1049;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_6_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_6_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h6 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_6_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_6_jmp_valid <= _GEN_1048;
      end
    end else begin
      ecp_6_jmp_valid <= _GEN_1048;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_5_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_5_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h5 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_5_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_5_jmp_valid <= _GEN_1047;
      end
    end else begin
      ecp_5_jmp_valid <= _GEN_1047;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_4_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_4_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h4 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_4_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_4_jmp_valid <= _GEN_1046;
      end
    end else begin
      ecp_4_jmp_valid <= _GEN_1046;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_3_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_3_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h3 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_3_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_3_jmp_valid <= _GEN_1045;
      end
    end else begin
      ecp_3_jmp_valid <= _GEN_1045;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_2_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_2_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h2 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_2_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_2_jmp_valid <= _GEN_1044;
      end
    end else begin
      ecp_2_jmp_valid <= _GEN_1044;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_1_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_1_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h1 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_1_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_1_jmp_valid <= _GEN_1043;
      end
    end else begin
      ecp_1_jmp_valid <= _GEN_1043;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_0_jmp_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_0_jmp_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h0 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_0_jmp_valid <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_0_jmp_valid <= _GEN_1042;
      end
    end else begin
      ecp_0_jmp_valid <= _GEN_1042;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_15_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_15_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hf == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_15_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_15_mis <= _GEN_1009;
      end
    end else begin
      ecp_15_mis <= _GEN_1009;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_14_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_14_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'he == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_14_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_14_mis <= _GEN_1008;
      end
    end else begin
      ecp_14_mis <= _GEN_1008;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_13_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_13_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hd == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_13_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_13_mis <= _GEN_1007;
      end
    end else begin
      ecp_13_mis <= _GEN_1007;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_12_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_12_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hc == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_12_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_12_mis <= _GEN_1006;
      end
    end else begin
      ecp_12_mis <= _GEN_1006;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_11_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_11_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hb == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_11_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_11_mis <= _GEN_1005;
      end
    end else begin
      ecp_11_mis <= _GEN_1005;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_10_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_10_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'ha == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_10_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_10_mis <= _GEN_1004;
      end
    end else begin
      ecp_10_mis <= _GEN_1004;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_9_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_9_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h9 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_9_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_9_mis <= _GEN_1003;
      end
    end else begin
      ecp_9_mis <= _GEN_1003;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_8_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_8_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h8 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_8_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_8_mis <= _GEN_1002;
      end
    end else begin
      ecp_8_mis <= _GEN_1002;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_7_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_7_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h7 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_7_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_7_mis <= _GEN_1001;
      end
    end else begin
      ecp_7_mis <= _GEN_1001;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_6_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_6_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h6 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_6_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_6_mis <= _GEN_1000;
      end
    end else begin
      ecp_6_mis <= _GEN_1000;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_5_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_5_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h5 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_5_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_5_mis <= _GEN_999;
      end
    end else begin
      ecp_5_mis <= _GEN_999;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_4_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_4_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h4 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_4_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_4_mis <= _GEN_998;
      end
    end else begin
      ecp_4_mis <= _GEN_998;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_3_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_3_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h3 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_3_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_3_mis <= _GEN_997;
      end
    end else begin
      ecp_3_mis <= _GEN_997;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_2_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_2_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h2 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_2_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_2_mis <= _GEN_996;
      end
    end else begin
      ecp_2_mis <= _GEN_996;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_1_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_1_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h1 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_1_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_1_mis <= _GEN_995;
      end
    end else begin
      ecp_1_mis <= _GEN_995;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_0_mis <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_0_mis <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h0 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_0_mis <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_0_mis <= _GEN_994;
      end
    end else begin
      ecp_0_mis <= _GEN_994;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_15_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_15_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hf == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_15_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_15_store_valid <= _GEN_1089;
      end
    end else begin
      ecp_15_store_valid <= _GEN_1089;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_14_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_14_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'he == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_14_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_14_store_valid <= _GEN_1088;
      end
    end else begin
      ecp_14_store_valid <= _GEN_1088;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_13_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_13_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hd == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_13_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_13_store_valid <= _GEN_1087;
      end
    end else begin
      ecp_13_store_valid <= _GEN_1087;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_12_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_12_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hc == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_12_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_12_store_valid <= _GEN_1086;
      end
    end else begin
      ecp_12_store_valid <= _GEN_1086;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_11_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_11_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hb == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_11_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_11_store_valid <= _GEN_1085;
      end
    end else begin
      ecp_11_store_valid <= _GEN_1085;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_10_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_10_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'ha == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_10_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_10_store_valid <= _GEN_1084;
      end
    end else begin
      ecp_10_store_valid <= _GEN_1084;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_9_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_9_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h9 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_9_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_9_store_valid <= _GEN_1083;
      end
    end else begin
      ecp_9_store_valid <= _GEN_1083;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_8_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_8_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h8 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_8_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_8_store_valid <= _GEN_1082;
      end
    end else begin
      ecp_8_store_valid <= _GEN_1082;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_7_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_7_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h7 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_7_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_7_store_valid <= _GEN_1081;
      end
    end else begin
      ecp_7_store_valid <= _GEN_1081;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_6_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_6_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h6 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_6_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_6_store_valid <= _GEN_1080;
      end
    end else begin
      ecp_6_store_valid <= _GEN_1080;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_5_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_5_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h5 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_5_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_5_store_valid <= _GEN_1079;
      end
    end else begin
      ecp_5_store_valid <= _GEN_1079;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_4_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_4_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h4 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_4_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_4_store_valid <= _GEN_1078;
      end
    end else begin
      ecp_4_store_valid <= _GEN_1078;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_3_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_3_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h3 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_3_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_3_store_valid <= _GEN_1077;
      end
    end else begin
      ecp_3_store_valid <= _GEN_1077;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_2_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_2_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h2 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_2_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_2_store_valid <= _GEN_1076;
      end
    end else begin
      ecp_2_store_valid <= _GEN_1076;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_1_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_1_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h1 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_1_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_1_store_valid <= _GEN_1075;
      end
    end else begin
      ecp_1_store_valid <= _GEN_1075;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_0_store_valid <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_0_store_valid <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h0 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_0_store_valid <= io_exe_ecp_2_store_valid; // @[Rob.scala 115:21]
      end else begin
        ecp_0_store_valid <= _GEN_1074;
      end
    end else begin
      ecp_0_store_valid <= _GEN_1074;
    end
    enq_ready <= reset | _GEN_1671; // @[Rob.scala 65:{26,26}]
    if (reset) begin // @[Rob.scala 71:20]
      ecp_0_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_0_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h0 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_0_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_0_jmp <= _GEN_1026;
      end
    end else begin
      ecp_0_jmp <= _GEN_1026;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_0_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_0_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h0 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_0_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_0_jmp_pc <= _GEN_1010;
      end
    end else begin
      ecp_0_jmp_pc <= _GEN_1010;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_1_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_1_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h1 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_1_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_1_jmp <= _GEN_1027;
      end
    end else begin
      ecp_1_jmp <= _GEN_1027;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_1_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_1_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h1 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_1_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_1_jmp_pc <= _GEN_1011;
      end
    end else begin
      ecp_1_jmp_pc <= _GEN_1011;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_2_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_2_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h2 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_2_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_2_jmp <= _GEN_1028;
      end
    end else begin
      ecp_2_jmp <= _GEN_1028;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_2_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_2_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h2 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_2_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_2_jmp_pc <= _GEN_1012;
      end
    end else begin
      ecp_2_jmp_pc <= _GEN_1012;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_3_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_3_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h3 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_3_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_3_jmp <= _GEN_1029;
      end
    end else begin
      ecp_3_jmp <= _GEN_1029;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_3_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_3_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h3 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_3_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_3_jmp_pc <= _GEN_1013;
      end
    end else begin
      ecp_3_jmp_pc <= _GEN_1013;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_4_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_4_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h4 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_4_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_4_jmp <= _GEN_1030;
      end
    end else begin
      ecp_4_jmp <= _GEN_1030;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_4_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_4_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h4 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_4_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_4_jmp_pc <= _GEN_1014;
      end
    end else begin
      ecp_4_jmp_pc <= _GEN_1014;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_5_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_5_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h5 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_5_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_5_jmp <= _GEN_1031;
      end
    end else begin
      ecp_5_jmp <= _GEN_1031;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_5_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_5_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h5 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_5_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_5_jmp_pc <= _GEN_1015;
      end
    end else begin
      ecp_5_jmp_pc <= _GEN_1015;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_6_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_6_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h6 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_6_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_6_jmp <= _GEN_1032;
      end
    end else begin
      ecp_6_jmp <= _GEN_1032;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_6_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_6_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h6 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_6_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_6_jmp_pc <= _GEN_1016;
      end
    end else begin
      ecp_6_jmp_pc <= _GEN_1016;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_7_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_7_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h7 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_7_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_7_jmp <= _GEN_1033;
      end
    end else begin
      ecp_7_jmp <= _GEN_1033;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_7_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_7_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h7 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_7_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_7_jmp_pc <= _GEN_1017;
      end
    end else begin
      ecp_7_jmp_pc <= _GEN_1017;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_8_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_8_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h8 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_8_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_8_jmp <= _GEN_1034;
      end
    end else begin
      ecp_8_jmp <= _GEN_1034;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_8_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_8_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h8 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_8_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_8_jmp_pc <= _GEN_1018;
      end
    end else begin
      ecp_8_jmp_pc <= _GEN_1018;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_9_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_9_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h9 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_9_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_9_jmp <= _GEN_1035;
      end
    end else begin
      ecp_9_jmp <= _GEN_1035;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_9_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_9_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'h9 == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_9_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_9_jmp_pc <= _GEN_1019;
      end
    end else begin
      ecp_9_jmp_pc <= _GEN_1019;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_10_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_10_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'ha == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_10_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_10_jmp <= _GEN_1036;
      end
    end else begin
      ecp_10_jmp <= _GEN_1036;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_10_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_10_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'ha == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_10_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_10_jmp_pc <= _GEN_1020;
      end
    end else begin
      ecp_10_jmp_pc <= _GEN_1020;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_11_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_11_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hb == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_11_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_11_jmp <= _GEN_1037;
      end
    end else begin
      ecp_11_jmp <= _GEN_1037;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_11_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_11_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hb == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_11_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_11_jmp_pc <= _GEN_1021;
      end
    end else begin
      ecp_11_jmp_pc <= _GEN_1021;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_12_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_12_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hc == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_12_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_12_jmp <= _GEN_1038;
      end
    end else begin
      ecp_12_jmp <= _GEN_1038;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_12_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_12_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hc == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_12_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_12_jmp_pc <= _GEN_1022;
      end
    end else begin
      ecp_12_jmp_pc <= _GEN_1022;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_13_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_13_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hd == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_13_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_13_jmp <= _GEN_1039;
      end
    end else begin
      ecp_13_jmp <= _GEN_1039;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_13_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_13_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hd == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_13_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_13_jmp_pc <= _GEN_1023;
      end
    end else begin
      ecp_13_jmp_pc <= _GEN_1023;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_14_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_14_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'he == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_14_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_14_jmp <= _GEN_1040;
      end
    end else begin
      ecp_14_jmp <= _GEN_1040;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_14_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_14_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'he == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_14_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_14_jmp_pc <= _GEN_1024;
      end
    end else begin
      ecp_14_jmp_pc <= _GEN_1024;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_15_jmp <= 1'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_15_jmp <= 1'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hf == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_15_jmp <= 1'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_15_jmp <= _GEN_1041;
      end
    end else begin
      ecp_15_jmp <= _GEN_1041;
    end
    if (reset) begin // @[Rob.scala 71:20]
      ecp_15_jmp_pc <= 32'h0; // @[Rob.scala 71:20]
    end else if (io_flush) begin // @[Rob.scala 332:19]
      ecp_15_jmp_pc <= 32'h0; // @[Rob.scala 335:9]
    end else if (io_exe_2_valid) begin // @[Rob.scala 113:28]
      if (4'hf == io_exe_2_rob_addr) begin // @[Rob.scala 115:21]
        ecp_15_jmp_pc <= 32'h0; // @[Rob.scala 115:21]
      end else begin
        ecp_15_jmp_pc <= _GEN_1025;
      end
    end else begin
      ecp_15_jmp_pc <= _GEN_1025;
    end
    if (reset) begin // @[Rob.scala 152:30]
      sys_in_flight <= 1'h0; // @[Rob.scala 152:30]
    end else if (cm_1_valid & sys_in_flight) begin // @[Rob.scala 265:41]
      sys_in_flight <= 1'h0; // @[Rob.scala 266:21]
    end else if (cm_0_valid & sys_in_flight) begin // @[Rob.scala 265:41]
      sys_in_flight <= 1'h0; // @[Rob.scala 266:21]
    end else begin
      sys_in_flight <= _GEN_1520;
    end
    if (reset) begin // @[Rob.scala 183:27]
      intr_state <= 1'h0; // @[Rob.scala 183:27]
    end else if (~intr_state) begin // @[Rob.scala 190:23]
      intr_state <= _GEN_1378;
    end else if (intr_state) begin // @[Rob.scala 190:23]
      intr_state <= _GEN_1390;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    rob_pc[initvar] = _RAND_0[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    rob_fu_code[initvar] = _RAND_5[2:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    rob_sys_code[initvar] = _RAND_10[2:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    rob_rd_addr[initvar] = _RAND_15[4:0];
  _RAND_20 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    rob_rd_en[initvar] = _RAND_20[0:0];
  _RAND_25 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    rob_rd_paddr[initvar] = _RAND_25[5:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    rob_rd_ppaddr[initvar] = _RAND_30[5:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
//   rob_pc_MPORT_2_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  rob_pc_MPORT_2_addr_pipe_0 = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
//   rob_pc_MPORT_3_en_pipe_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  rob_pc_MPORT_3_addr_pipe_0 = _RAND_4[3:0];
  _RAND_6 = {1{`RANDOM}};
//   rob_fu_code_MPORT_2_en_pipe_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  rob_fu_code_MPORT_2_addr_pipe_0 = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
//   rob_fu_code_MPORT_3_en_pipe_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  rob_fu_code_MPORT_3_addr_pipe_0 = _RAND_9[3:0];
  _RAND_11 = {1{`RANDOM}};
//   rob_sys_code_MPORT_2_en_pipe_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  rob_sys_code_MPORT_2_addr_pipe_0 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
//   rob_sys_code_MPORT_3_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  rob_sys_code_MPORT_3_addr_pipe_0 = _RAND_14[3:0];
  _RAND_16 = {1{`RANDOM}};
//   rob_rd_addr_MPORT_2_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  rob_rd_addr_MPORT_2_addr_pipe_0 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
//   rob_rd_addr_MPORT_3_en_pipe_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  rob_rd_addr_MPORT_3_addr_pipe_0 = _RAND_19[3:0];
  _RAND_21 = {1{`RANDOM}};
//   rob_rd_en_MPORT_2_en_pipe_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  rob_rd_en_MPORT_2_addr_pipe_0 = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
//   rob_rd_en_MPORT_3_en_pipe_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  rob_rd_en_MPORT_3_addr_pipe_0 = _RAND_24[3:0];
  _RAND_26 = {1{`RANDOM}};
//   rob_rd_paddr_MPORT_2_en_pipe_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  rob_rd_paddr_MPORT_2_addr_pipe_0 = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
//   rob_rd_paddr_MPORT_3_en_pipe_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  rob_rd_paddr_MPORT_3_addr_pipe_0 = _RAND_29[3:0];
  _RAND_31 = {1{`RANDOM}};
//   rob_rd_ppaddr_MPORT_2_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  rob_rd_ppaddr_MPORT_2_addr_pipe_0 = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
//   rob_rd_ppaddr_MPORT_3_en_pipe_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  rob_rd_ppaddr_MPORT_3_addr_pipe_0 = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  enq_vec_0 = _RAND_35[4:0];
  _RAND_36 = {1{`RANDOM}};
  enq_vec_1 = _RAND_36[4:0];
  _RAND_37 = {1{`RANDOM}};
  deq_vec_0 = _RAND_37[4:0];
  _RAND_38 = {1{`RANDOM}};
  deq_vec_1 = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  complete_15 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  complete_14 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  complete_13 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  complete_12 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  complete_11 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  complete_10 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  complete_9 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  complete_8 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  complete_7 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  complete_6 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  complete_5 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  complete_4 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  complete_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  complete_2 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  complete_1 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  complete_0 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  ecp_15_jmp_valid = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  ecp_14_jmp_valid = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  ecp_13_jmp_valid = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  ecp_12_jmp_valid = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  ecp_11_jmp_valid = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  ecp_10_jmp_valid = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  ecp_9_jmp_valid = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  ecp_8_jmp_valid = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  ecp_7_jmp_valid = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  ecp_6_jmp_valid = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  ecp_5_jmp_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  ecp_4_jmp_valid = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  ecp_3_jmp_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  ecp_2_jmp_valid = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  ecp_1_jmp_valid = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  ecp_0_jmp_valid = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  ecp_15_mis = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  ecp_14_mis = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  ecp_13_mis = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  ecp_12_mis = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  ecp_11_mis = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  ecp_10_mis = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  ecp_9_mis = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  ecp_8_mis = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  ecp_7_mis = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  ecp_6_mis = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  ecp_5_mis = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  ecp_4_mis = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  ecp_3_mis = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  ecp_2_mis = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  ecp_1_mis = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  ecp_0_mis = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  ecp_15_store_valid = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  ecp_14_store_valid = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  ecp_13_store_valid = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  ecp_12_store_valid = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  ecp_11_store_valid = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  ecp_10_store_valid = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  ecp_9_store_valid = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  ecp_8_store_valid = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  ecp_7_store_valid = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  ecp_6_store_valid = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  ecp_5_store_valid = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  ecp_4_store_valid = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  ecp_3_store_valid = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  ecp_2_store_valid = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  ecp_1_store_valid = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  ecp_0_store_valid = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  enq_ready = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  ecp_0_jmp = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  ecp_0_jmp_pc = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  ecp_1_jmp = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  ecp_1_jmp_pc = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  ecp_2_jmp = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  ecp_2_jmp_pc = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  ecp_3_jmp = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  ecp_3_jmp_pc = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  ecp_4_jmp = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  ecp_4_jmp_pc = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  ecp_5_jmp = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  ecp_5_jmp_pc = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  ecp_6_jmp = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  ecp_6_jmp_pc = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  ecp_7_jmp = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  ecp_7_jmp_pc = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  ecp_8_jmp = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  ecp_8_jmp_pc = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  ecp_9_jmp = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  ecp_9_jmp_pc = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  ecp_10_jmp = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  ecp_10_jmp_pc = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  ecp_11_jmp = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  ecp_11_jmp_pc = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  ecp_12_jmp = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  ecp_12_jmp_pc = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  ecp_13_jmp = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  ecp_13_jmp_pc = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  ecp_14_jmp = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  ecp_14_jmp_pc = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  ecp_15_jmp = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  ecp_15_jmp_pc = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  sys_in_flight = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  intr_state = _RAND_137[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_IntIssueQueueOutOfOrder(
  input         clock,
  input         reset,
  input         io_flush,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_vec_0_valid,
  input  [31:0] io_in_bits_vec_0_pc,
  input  [31:0] io_in_bits_vec_0_npc,
  input  [31:0] io_in_bits_vec_0_inst,
  input  [2:0]  io_in_bits_vec_0_fu_code,
  input  [3:0]  io_in_bits_vec_0_alu_code,
  input  [3:0]  io_in_bits_vec_0_jmp_code,
  input  [2:0]  io_in_bits_vec_0_sys_code,
  input         io_in_bits_vec_0_w_type,
  input  [1:0]  io_in_bits_vec_0_rs1_src,
  input  [1:0]  io_in_bits_vec_0_rs2_src,
  input         io_in_bits_vec_0_rd_en,
  input  [31:0] io_in_bits_vec_0_imm,
  input         io_in_bits_vec_0_pred_br,
  input  [31:0] io_in_bits_vec_0_pred_bpc,
  input  [5:0]  io_in_bits_vec_0_rs1_paddr,
  input  [5:0]  io_in_bits_vec_0_rs2_paddr,
  input  [5:0]  io_in_bits_vec_0_rd_paddr,
  input         io_in_bits_vec_1_valid,
  input  [31:0] io_in_bits_vec_1_pc,
  input  [31:0] io_in_bits_vec_1_npc,
  input  [31:0] io_in_bits_vec_1_inst,
  input  [2:0]  io_in_bits_vec_1_fu_code,
  input  [3:0]  io_in_bits_vec_1_alu_code,
  input  [3:0]  io_in_bits_vec_1_jmp_code,
  input  [2:0]  io_in_bits_vec_1_sys_code,
  input         io_in_bits_vec_1_w_type,
  input  [1:0]  io_in_bits_vec_1_rs1_src,
  input  [1:0]  io_in_bits_vec_1_rs2_src,
  input         io_in_bits_vec_1_rd_en,
  input  [31:0] io_in_bits_vec_1_imm,
  input         io_in_bits_vec_1_pred_br,
  input  [31:0] io_in_bits_vec_1_pred_bpc,
  input  [5:0]  io_in_bits_vec_1_rs1_paddr,
  input  [5:0]  io_in_bits_vec_1_rs2_paddr,
  input  [5:0]  io_in_bits_vec_1_rd_paddr,
  input  [3:0]  io_rob_addr_0,
  input  [3:0]  io_rob_addr_1,
  output        io_out_0_valid,
  output [31:0] io_out_0_pc,
  output [31:0] io_out_0_npc,
  output [31:0] io_out_0_inst,
  output [2:0]  io_out_0_fu_code,
  output [3:0]  io_out_0_alu_code,
  output [3:0]  io_out_0_jmp_code,
  output [2:0]  io_out_0_sys_code,
  output        io_out_0_w_type,
  output [1:0]  io_out_0_rs1_src,
  output [1:0]  io_out_0_rs2_src,
  output        io_out_0_rd_en,
  output [31:0] io_out_0_imm,
  output        io_out_0_pred_br,
  output [31:0] io_out_0_pred_bpc,
  output [5:0]  io_out_0_rs1_paddr,
  output [5:0]  io_out_0_rs2_paddr,
  output [5:0]  io_out_0_rd_paddr,
  output [3:0]  io_out_0_rob_addr,
  output        io_out_1_valid,
  output [31:0] io_out_1_pc,
  output [31:0] io_out_1_npc,
  output [2:0]  io_out_1_fu_code,
  output [3:0]  io_out_1_alu_code,
  output [3:0]  io_out_1_jmp_code,
  output        io_out_1_w_type,
  output [1:0]  io_out_1_rs1_src,
  output [1:0]  io_out_1_rs2_src,
  output        io_out_1_rd_en,
  output [31:0] io_out_1_imm,
  output        io_out_1_pred_br,
  output [31:0] io_out_1_pred_bpc,
  output [5:0]  io_out_1_rs1_paddr,
  output [5:0]  io_out_1_rs2_paddr,
  output [5:0]  io_out_1_rd_paddr,
  output [3:0]  io_out_1_rob_addr,
  input         io_avail_list_0,
  input         io_avail_list_1,
  input         io_avail_list_2,
  input         io_avail_list_3,
  input         io_avail_list_4,
  input         io_avail_list_5,
  input         io_avail_list_6,
  input         io_avail_list_7,
  input         io_avail_list_8,
  input         io_avail_list_9,
  input         io_avail_list_10,
  input         io_avail_list_11,
  input         io_avail_list_12,
  input         io_avail_list_13,
  input         io_avail_list_14,
  input         io_avail_list_15,
  input         io_avail_list_16,
  input         io_avail_list_17,
  input         io_avail_list_18,
  input         io_avail_list_19,
  input         io_avail_list_20,
  input         io_avail_list_21,
  input         io_avail_list_22,
  input         io_avail_list_23,
  input         io_avail_list_24,
  input         io_avail_list_25,
  input         io_avail_list_26,
  input         io_avail_list_27,
  input         io_avail_list_28,
  input         io_avail_list_29,
  input         io_avail_list_30,
  input         io_avail_list_31,
  input         io_avail_list_32,
  input         io_avail_list_33,
  input         io_avail_list_34,
  input         io_avail_list_35,
  input         io_avail_list_36,
  input         io_avail_list_37,
  input         io_avail_list_38,
  input         io_avail_list_39,
  input         io_avail_list_40,
  input         io_avail_list_41,
  input         io_avail_list_42,
  input         io_avail_list_43,
  input         io_avail_list_44,
  input         io_avail_list_45,
  input         io_avail_list_46,
  input         io_avail_list_47,
  input         io_avail_list_48,
  input         io_avail_list_49,
  input         io_avail_list_50,
  input         io_avail_list_51,
  input         io_avail_list_52,
  input         io_avail_list_53,
  input         io_avail_list_54,
  input         io_avail_list_55,
  input         io_avail_list_56,
  input         io_avail_list_57,
  input         io_avail_list_58,
  input         io_avail_list_59,
  input         io_avail_list_60,
  input         io_avail_list_61,
  input         io_avail_list_62,
  input         io_avail_list_63,
  input         io_sys_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
`endif // RANDOMIZE_REG_INIT
  reg  buf_0_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_0_pc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_0_npc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_0_inst; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_0_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_0_alu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_0_jmp_code; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_0_sys_code; // @[IssueUnit.scala 97:20]
  reg  buf_0_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_0_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_0_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_0_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_0_imm; // @[IssueUnit.scala 97:20]
  reg  buf_0_pred_br; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_0_pred_bpc; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_0_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_0_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_0_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_0_rob_addr; // @[IssueUnit.scala 97:20]
  reg  buf_1_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_1_pc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_1_npc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_1_inst; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_1_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_1_alu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_1_jmp_code; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_1_sys_code; // @[IssueUnit.scala 97:20]
  reg  buf_1_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_1_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_1_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_1_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_1_imm; // @[IssueUnit.scala 97:20]
  reg  buf_1_pred_br; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_1_pred_bpc; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_1_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_1_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_1_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_1_rob_addr; // @[IssueUnit.scala 97:20]
  reg  buf_2_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_2_pc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_2_npc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_2_inst; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_2_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_2_alu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_2_jmp_code; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_2_sys_code; // @[IssueUnit.scala 97:20]
  reg  buf_2_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_2_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_2_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_2_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_2_imm; // @[IssueUnit.scala 97:20]
  reg  buf_2_pred_br; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_2_pred_bpc; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_2_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_2_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_2_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_2_rob_addr; // @[IssueUnit.scala 97:20]
  reg  buf_3_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_3_pc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_3_npc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_3_inst; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_3_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_3_alu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_3_jmp_code; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_3_sys_code; // @[IssueUnit.scala 97:20]
  reg  buf_3_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_3_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_3_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_3_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_3_imm; // @[IssueUnit.scala 97:20]
  reg  buf_3_pred_br; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_3_pred_bpc; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_3_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_3_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_3_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_3_rob_addr; // @[IssueUnit.scala 97:20]
  reg  buf_4_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_4_pc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_4_npc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_4_inst; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_4_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_4_alu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_4_jmp_code; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_4_sys_code; // @[IssueUnit.scala 97:20]
  reg  buf_4_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_4_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_4_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_4_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_4_imm; // @[IssueUnit.scala 97:20]
  reg  buf_4_pred_br; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_4_pred_bpc; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_4_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_4_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_4_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_4_rob_addr; // @[IssueUnit.scala 97:20]
  reg  buf_5_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_5_pc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_5_npc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_5_inst; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_5_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_5_alu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_5_jmp_code; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_5_sys_code; // @[IssueUnit.scala 97:20]
  reg  buf_5_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_5_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_5_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_5_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_5_imm; // @[IssueUnit.scala 97:20]
  reg  buf_5_pred_br; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_5_pred_bpc; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_5_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_5_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_5_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_5_rob_addr; // @[IssueUnit.scala 97:20]
  reg  buf_6_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_6_pc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_6_npc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_6_inst; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_6_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_6_alu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_6_jmp_code; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_6_sys_code; // @[IssueUnit.scala 97:20]
  reg  buf_6_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_6_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_6_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_6_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_6_imm; // @[IssueUnit.scala 97:20]
  reg  buf_6_pred_br; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_6_pred_bpc; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_6_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_6_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_6_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_6_rob_addr; // @[IssueUnit.scala 97:20]
  reg  buf_7_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_7_pc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_7_npc; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_7_inst; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_7_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_7_alu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_7_jmp_code; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_7_sys_code; // @[IssueUnit.scala 97:20]
  reg  buf_7_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_7_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_7_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_7_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_7_imm; // @[IssueUnit.scala 97:20]
  reg  buf_7_pred_br; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_7_pred_bpc; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_7_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_7_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_7_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_7_rob_addr; // @[IssueUnit.scala 97:20]
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_1 = io_in_bits_vec_0_valid + io_in_bits_vec_1_valid; // @[Bitwise.scala 47:55]
  wire [1:0] num_enq = _T ? _T_1 : 2'h0; // @[IssueUnit.scala 99:20]
  wire [1:0] num_deq = io_out_0_valid + io_out_1_valid; // @[Bitwise.scala 47:55]
  reg [3:0] enq_vec_0; // @[IssueUnit.scala 102:24]
  reg [3:0] enq_vec_1; // @[IssueUnit.scala 102:24]
  wire [3:0] _GEN_2848 = {{2'd0}, num_deq}; // @[IssueUnit.scala 103:44]
  wire [3:0] enq_vec_real_0 = enq_vec_0 - _GEN_2848; // @[IssueUnit.scala 103:44]
  wire [3:0] enq_vec_real_1 = enq_vec_1 - _GEN_2848; // @[IssueUnit.scala 103:44]
  wire  enq_ready = enq_vec_real_0 <= 4'h6; // @[IssueUnit.scala 106:27]
  wire  is_sys_0 = buf_0_fu_code == 3'h3; // @[IssueUnit.scala 115:34]
  wire  is_sys_1 = buf_1_fu_code == 3'h3; // @[IssueUnit.scala 115:34]
  wire  is_sys_2 = buf_2_fu_code == 3'h3; // @[IssueUnit.scala 115:34]
  wire  is_sys_3 = buf_3_fu_code == 3'h3; // @[IssueUnit.scala 115:34]
  wire  is_sys_4 = buf_4_fu_code == 3'h3; // @[IssueUnit.scala 115:34]
  wire  is_sys_5 = buf_5_fu_code == 3'h3; // @[IssueUnit.scala 115:34]
  wire  is_sys_6 = buf_6_fu_code == 3'h3; // @[IssueUnit.scala 115:34]
  wire  is_sys_7 = buf_7_fu_code == 3'h3; // @[IssueUnit.scala 115:34]
  wire [7:0] _T_16 = {is_sys_0,is_sys_1,is_sys_2,is_sys_3,is_sys_4,is_sys_5,is_sys_6,is_sys_7}; // @[Cat.scala 30:58]
  wire  has_sys = |_T_16; // @[IssueUnit.scala 117:29]
  wire  _GEN_1 = 6'h1 == buf_0_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_2 = 6'h2 == buf_0_rs1_paddr ? io_avail_list_2 : _GEN_1; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_3 = 6'h3 == buf_0_rs1_paddr ? io_avail_list_3 : _GEN_2; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_4 = 6'h4 == buf_0_rs1_paddr ? io_avail_list_4 : _GEN_3; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_5 = 6'h5 == buf_0_rs1_paddr ? io_avail_list_5 : _GEN_4; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_6 = 6'h6 == buf_0_rs1_paddr ? io_avail_list_6 : _GEN_5; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_7 = 6'h7 == buf_0_rs1_paddr ? io_avail_list_7 : _GEN_6; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_8 = 6'h8 == buf_0_rs1_paddr ? io_avail_list_8 : _GEN_7; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_9 = 6'h9 == buf_0_rs1_paddr ? io_avail_list_9 : _GEN_8; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_10 = 6'ha == buf_0_rs1_paddr ? io_avail_list_10 : _GEN_9; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_11 = 6'hb == buf_0_rs1_paddr ? io_avail_list_11 : _GEN_10; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_12 = 6'hc == buf_0_rs1_paddr ? io_avail_list_12 : _GEN_11; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_13 = 6'hd == buf_0_rs1_paddr ? io_avail_list_13 : _GEN_12; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_14 = 6'he == buf_0_rs1_paddr ? io_avail_list_14 : _GEN_13; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_15 = 6'hf == buf_0_rs1_paddr ? io_avail_list_15 : _GEN_14; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_16 = 6'h10 == buf_0_rs1_paddr ? io_avail_list_16 : _GEN_15; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_17 = 6'h11 == buf_0_rs1_paddr ? io_avail_list_17 : _GEN_16; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_18 = 6'h12 == buf_0_rs1_paddr ? io_avail_list_18 : _GEN_17; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_19 = 6'h13 == buf_0_rs1_paddr ? io_avail_list_19 : _GEN_18; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_20 = 6'h14 == buf_0_rs1_paddr ? io_avail_list_20 : _GEN_19; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_21 = 6'h15 == buf_0_rs1_paddr ? io_avail_list_21 : _GEN_20; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_22 = 6'h16 == buf_0_rs1_paddr ? io_avail_list_22 : _GEN_21; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_23 = 6'h17 == buf_0_rs1_paddr ? io_avail_list_23 : _GEN_22; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_24 = 6'h18 == buf_0_rs1_paddr ? io_avail_list_24 : _GEN_23; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_25 = 6'h19 == buf_0_rs1_paddr ? io_avail_list_25 : _GEN_24; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_26 = 6'h1a == buf_0_rs1_paddr ? io_avail_list_26 : _GEN_25; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_27 = 6'h1b == buf_0_rs1_paddr ? io_avail_list_27 : _GEN_26; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_28 = 6'h1c == buf_0_rs1_paddr ? io_avail_list_28 : _GEN_27; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_29 = 6'h1d == buf_0_rs1_paddr ? io_avail_list_29 : _GEN_28; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_30 = 6'h1e == buf_0_rs1_paddr ? io_avail_list_30 : _GEN_29; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_31 = 6'h1f == buf_0_rs1_paddr ? io_avail_list_31 : _GEN_30; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_32 = 6'h20 == buf_0_rs1_paddr ? io_avail_list_32 : _GEN_31; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_33 = 6'h21 == buf_0_rs1_paddr ? io_avail_list_33 : _GEN_32; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_34 = 6'h22 == buf_0_rs1_paddr ? io_avail_list_34 : _GEN_33; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_35 = 6'h23 == buf_0_rs1_paddr ? io_avail_list_35 : _GEN_34; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_36 = 6'h24 == buf_0_rs1_paddr ? io_avail_list_36 : _GEN_35; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_37 = 6'h25 == buf_0_rs1_paddr ? io_avail_list_37 : _GEN_36; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_38 = 6'h26 == buf_0_rs1_paddr ? io_avail_list_38 : _GEN_37; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_39 = 6'h27 == buf_0_rs1_paddr ? io_avail_list_39 : _GEN_38; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_40 = 6'h28 == buf_0_rs1_paddr ? io_avail_list_40 : _GEN_39; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_41 = 6'h29 == buf_0_rs1_paddr ? io_avail_list_41 : _GEN_40; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_42 = 6'h2a == buf_0_rs1_paddr ? io_avail_list_42 : _GEN_41; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_43 = 6'h2b == buf_0_rs1_paddr ? io_avail_list_43 : _GEN_42; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_44 = 6'h2c == buf_0_rs1_paddr ? io_avail_list_44 : _GEN_43; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_45 = 6'h2d == buf_0_rs1_paddr ? io_avail_list_45 : _GEN_44; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_46 = 6'h2e == buf_0_rs1_paddr ? io_avail_list_46 : _GEN_45; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_47 = 6'h2f == buf_0_rs1_paddr ? io_avail_list_47 : _GEN_46; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_48 = 6'h30 == buf_0_rs1_paddr ? io_avail_list_48 : _GEN_47; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_49 = 6'h31 == buf_0_rs1_paddr ? io_avail_list_49 : _GEN_48; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_50 = 6'h32 == buf_0_rs1_paddr ? io_avail_list_50 : _GEN_49; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_51 = 6'h33 == buf_0_rs1_paddr ? io_avail_list_51 : _GEN_50; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_52 = 6'h34 == buf_0_rs1_paddr ? io_avail_list_52 : _GEN_51; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_53 = 6'h35 == buf_0_rs1_paddr ? io_avail_list_53 : _GEN_52; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_54 = 6'h36 == buf_0_rs1_paddr ? io_avail_list_54 : _GEN_53; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_55 = 6'h37 == buf_0_rs1_paddr ? io_avail_list_55 : _GEN_54; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_56 = 6'h38 == buf_0_rs1_paddr ? io_avail_list_56 : _GEN_55; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_57 = 6'h39 == buf_0_rs1_paddr ? io_avail_list_57 : _GEN_56; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_58 = 6'h3a == buf_0_rs1_paddr ? io_avail_list_58 : _GEN_57; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_59 = 6'h3b == buf_0_rs1_paddr ? io_avail_list_59 : _GEN_58; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_60 = 6'h3c == buf_0_rs1_paddr ? io_avail_list_60 : _GEN_59; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_61 = 6'h3d == buf_0_rs1_paddr ? io_avail_list_61 : _GEN_60; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_62 = 6'h3e == buf_0_rs1_paddr ? io_avail_list_62 : _GEN_61; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_63 = 6'h3f == buf_0_rs1_paddr ? io_avail_list_63 : _GEN_62; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_65 = 6'h1 == buf_0_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_66 = 6'h2 == buf_0_rs2_paddr ? io_avail_list_2 : _GEN_65; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_67 = 6'h3 == buf_0_rs2_paddr ? io_avail_list_3 : _GEN_66; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_68 = 6'h4 == buf_0_rs2_paddr ? io_avail_list_4 : _GEN_67; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_69 = 6'h5 == buf_0_rs2_paddr ? io_avail_list_5 : _GEN_68; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_70 = 6'h6 == buf_0_rs2_paddr ? io_avail_list_6 : _GEN_69; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_71 = 6'h7 == buf_0_rs2_paddr ? io_avail_list_7 : _GEN_70; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_72 = 6'h8 == buf_0_rs2_paddr ? io_avail_list_8 : _GEN_71; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_73 = 6'h9 == buf_0_rs2_paddr ? io_avail_list_9 : _GEN_72; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_74 = 6'ha == buf_0_rs2_paddr ? io_avail_list_10 : _GEN_73; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_75 = 6'hb == buf_0_rs2_paddr ? io_avail_list_11 : _GEN_74; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_76 = 6'hc == buf_0_rs2_paddr ? io_avail_list_12 : _GEN_75; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_77 = 6'hd == buf_0_rs2_paddr ? io_avail_list_13 : _GEN_76; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_78 = 6'he == buf_0_rs2_paddr ? io_avail_list_14 : _GEN_77; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_79 = 6'hf == buf_0_rs2_paddr ? io_avail_list_15 : _GEN_78; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_80 = 6'h10 == buf_0_rs2_paddr ? io_avail_list_16 : _GEN_79; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_81 = 6'h11 == buf_0_rs2_paddr ? io_avail_list_17 : _GEN_80; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_82 = 6'h12 == buf_0_rs2_paddr ? io_avail_list_18 : _GEN_81; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_83 = 6'h13 == buf_0_rs2_paddr ? io_avail_list_19 : _GEN_82; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_84 = 6'h14 == buf_0_rs2_paddr ? io_avail_list_20 : _GEN_83; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_85 = 6'h15 == buf_0_rs2_paddr ? io_avail_list_21 : _GEN_84; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_86 = 6'h16 == buf_0_rs2_paddr ? io_avail_list_22 : _GEN_85; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_87 = 6'h17 == buf_0_rs2_paddr ? io_avail_list_23 : _GEN_86; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_88 = 6'h18 == buf_0_rs2_paddr ? io_avail_list_24 : _GEN_87; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_89 = 6'h19 == buf_0_rs2_paddr ? io_avail_list_25 : _GEN_88; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_90 = 6'h1a == buf_0_rs2_paddr ? io_avail_list_26 : _GEN_89; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_91 = 6'h1b == buf_0_rs2_paddr ? io_avail_list_27 : _GEN_90; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_92 = 6'h1c == buf_0_rs2_paddr ? io_avail_list_28 : _GEN_91; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_93 = 6'h1d == buf_0_rs2_paddr ? io_avail_list_29 : _GEN_92; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_94 = 6'h1e == buf_0_rs2_paddr ? io_avail_list_30 : _GEN_93; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_95 = 6'h1f == buf_0_rs2_paddr ? io_avail_list_31 : _GEN_94; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_96 = 6'h20 == buf_0_rs2_paddr ? io_avail_list_32 : _GEN_95; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_97 = 6'h21 == buf_0_rs2_paddr ? io_avail_list_33 : _GEN_96; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_98 = 6'h22 == buf_0_rs2_paddr ? io_avail_list_34 : _GEN_97; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_99 = 6'h23 == buf_0_rs2_paddr ? io_avail_list_35 : _GEN_98; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_100 = 6'h24 == buf_0_rs2_paddr ? io_avail_list_36 : _GEN_99; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_101 = 6'h25 == buf_0_rs2_paddr ? io_avail_list_37 : _GEN_100; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_102 = 6'h26 == buf_0_rs2_paddr ? io_avail_list_38 : _GEN_101; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_103 = 6'h27 == buf_0_rs2_paddr ? io_avail_list_39 : _GEN_102; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_104 = 6'h28 == buf_0_rs2_paddr ? io_avail_list_40 : _GEN_103; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_105 = 6'h29 == buf_0_rs2_paddr ? io_avail_list_41 : _GEN_104; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_106 = 6'h2a == buf_0_rs2_paddr ? io_avail_list_42 : _GEN_105; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_107 = 6'h2b == buf_0_rs2_paddr ? io_avail_list_43 : _GEN_106; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_108 = 6'h2c == buf_0_rs2_paddr ? io_avail_list_44 : _GEN_107; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_109 = 6'h2d == buf_0_rs2_paddr ? io_avail_list_45 : _GEN_108; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_110 = 6'h2e == buf_0_rs2_paddr ? io_avail_list_46 : _GEN_109; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_111 = 6'h2f == buf_0_rs2_paddr ? io_avail_list_47 : _GEN_110; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_112 = 6'h30 == buf_0_rs2_paddr ? io_avail_list_48 : _GEN_111; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_113 = 6'h31 == buf_0_rs2_paddr ? io_avail_list_49 : _GEN_112; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_114 = 6'h32 == buf_0_rs2_paddr ? io_avail_list_50 : _GEN_113; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_115 = 6'h33 == buf_0_rs2_paddr ? io_avail_list_51 : _GEN_114; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_116 = 6'h34 == buf_0_rs2_paddr ? io_avail_list_52 : _GEN_115; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_117 = 6'h35 == buf_0_rs2_paddr ? io_avail_list_53 : _GEN_116; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_118 = 6'h36 == buf_0_rs2_paddr ? io_avail_list_54 : _GEN_117; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_119 = 6'h37 == buf_0_rs2_paddr ? io_avail_list_55 : _GEN_118; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_120 = 6'h38 == buf_0_rs2_paddr ? io_avail_list_56 : _GEN_119; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_121 = 6'h39 == buf_0_rs2_paddr ? io_avail_list_57 : _GEN_120; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_122 = 6'h3a == buf_0_rs2_paddr ? io_avail_list_58 : _GEN_121; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_123 = 6'h3b == buf_0_rs2_paddr ? io_avail_list_59 : _GEN_122; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_124 = 6'h3c == buf_0_rs2_paddr ? io_avail_list_60 : _GEN_123; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_125 = 6'h3d == buf_0_rs2_paddr ? io_avail_list_61 : _GEN_124; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_126 = 6'h3e == buf_0_rs2_paddr ? io_avail_list_62 : _GEN_125; // @[IssueUnit.scala 131:{34,34}]
  wire  _GEN_127 = 6'h3f == buf_0_rs2_paddr ? io_avail_list_63 : _GEN_126; // @[IssueUnit.scala 131:{34,34}]
  wire  ready_list_0 = _GEN_63 & _GEN_127 & (~is_sys_0 | is_sys_0 & io_sys_ready); // @[IssueUnit.scala 131:59]
  wire  _GEN_129 = 6'h1 == buf_1_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_130 = 6'h2 == buf_1_rs1_paddr ? io_avail_list_2 : _GEN_129; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_131 = 6'h3 == buf_1_rs1_paddr ? io_avail_list_3 : _GEN_130; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_132 = 6'h4 == buf_1_rs1_paddr ? io_avail_list_4 : _GEN_131; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_133 = 6'h5 == buf_1_rs1_paddr ? io_avail_list_5 : _GEN_132; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_134 = 6'h6 == buf_1_rs1_paddr ? io_avail_list_6 : _GEN_133; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_135 = 6'h7 == buf_1_rs1_paddr ? io_avail_list_7 : _GEN_134; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_136 = 6'h8 == buf_1_rs1_paddr ? io_avail_list_8 : _GEN_135; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_137 = 6'h9 == buf_1_rs1_paddr ? io_avail_list_9 : _GEN_136; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_138 = 6'ha == buf_1_rs1_paddr ? io_avail_list_10 : _GEN_137; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_139 = 6'hb == buf_1_rs1_paddr ? io_avail_list_11 : _GEN_138; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_140 = 6'hc == buf_1_rs1_paddr ? io_avail_list_12 : _GEN_139; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_141 = 6'hd == buf_1_rs1_paddr ? io_avail_list_13 : _GEN_140; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_142 = 6'he == buf_1_rs1_paddr ? io_avail_list_14 : _GEN_141; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_143 = 6'hf == buf_1_rs1_paddr ? io_avail_list_15 : _GEN_142; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_144 = 6'h10 == buf_1_rs1_paddr ? io_avail_list_16 : _GEN_143; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_145 = 6'h11 == buf_1_rs1_paddr ? io_avail_list_17 : _GEN_144; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_146 = 6'h12 == buf_1_rs1_paddr ? io_avail_list_18 : _GEN_145; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_147 = 6'h13 == buf_1_rs1_paddr ? io_avail_list_19 : _GEN_146; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_148 = 6'h14 == buf_1_rs1_paddr ? io_avail_list_20 : _GEN_147; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_149 = 6'h15 == buf_1_rs1_paddr ? io_avail_list_21 : _GEN_148; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_150 = 6'h16 == buf_1_rs1_paddr ? io_avail_list_22 : _GEN_149; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_151 = 6'h17 == buf_1_rs1_paddr ? io_avail_list_23 : _GEN_150; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_152 = 6'h18 == buf_1_rs1_paddr ? io_avail_list_24 : _GEN_151; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_153 = 6'h19 == buf_1_rs1_paddr ? io_avail_list_25 : _GEN_152; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_154 = 6'h1a == buf_1_rs1_paddr ? io_avail_list_26 : _GEN_153; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_155 = 6'h1b == buf_1_rs1_paddr ? io_avail_list_27 : _GEN_154; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_156 = 6'h1c == buf_1_rs1_paddr ? io_avail_list_28 : _GEN_155; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_157 = 6'h1d == buf_1_rs1_paddr ? io_avail_list_29 : _GEN_156; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_158 = 6'h1e == buf_1_rs1_paddr ? io_avail_list_30 : _GEN_157; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_159 = 6'h1f == buf_1_rs1_paddr ? io_avail_list_31 : _GEN_158; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_160 = 6'h20 == buf_1_rs1_paddr ? io_avail_list_32 : _GEN_159; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_161 = 6'h21 == buf_1_rs1_paddr ? io_avail_list_33 : _GEN_160; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_162 = 6'h22 == buf_1_rs1_paddr ? io_avail_list_34 : _GEN_161; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_163 = 6'h23 == buf_1_rs1_paddr ? io_avail_list_35 : _GEN_162; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_164 = 6'h24 == buf_1_rs1_paddr ? io_avail_list_36 : _GEN_163; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_165 = 6'h25 == buf_1_rs1_paddr ? io_avail_list_37 : _GEN_164; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_166 = 6'h26 == buf_1_rs1_paddr ? io_avail_list_38 : _GEN_165; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_167 = 6'h27 == buf_1_rs1_paddr ? io_avail_list_39 : _GEN_166; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_168 = 6'h28 == buf_1_rs1_paddr ? io_avail_list_40 : _GEN_167; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_169 = 6'h29 == buf_1_rs1_paddr ? io_avail_list_41 : _GEN_168; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_170 = 6'h2a == buf_1_rs1_paddr ? io_avail_list_42 : _GEN_169; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_171 = 6'h2b == buf_1_rs1_paddr ? io_avail_list_43 : _GEN_170; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_172 = 6'h2c == buf_1_rs1_paddr ? io_avail_list_44 : _GEN_171; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_173 = 6'h2d == buf_1_rs1_paddr ? io_avail_list_45 : _GEN_172; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_174 = 6'h2e == buf_1_rs1_paddr ? io_avail_list_46 : _GEN_173; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_175 = 6'h2f == buf_1_rs1_paddr ? io_avail_list_47 : _GEN_174; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_176 = 6'h30 == buf_1_rs1_paddr ? io_avail_list_48 : _GEN_175; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_177 = 6'h31 == buf_1_rs1_paddr ? io_avail_list_49 : _GEN_176; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_178 = 6'h32 == buf_1_rs1_paddr ? io_avail_list_50 : _GEN_177; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_179 = 6'h33 == buf_1_rs1_paddr ? io_avail_list_51 : _GEN_178; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_180 = 6'h34 == buf_1_rs1_paddr ? io_avail_list_52 : _GEN_179; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_181 = 6'h35 == buf_1_rs1_paddr ? io_avail_list_53 : _GEN_180; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_182 = 6'h36 == buf_1_rs1_paddr ? io_avail_list_54 : _GEN_181; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_183 = 6'h37 == buf_1_rs1_paddr ? io_avail_list_55 : _GEN_182; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_184 = 6'h38 == buf_1_rs1_paddr ? io_avail_list_56 : _GEN_183; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_185 = 6'h39 == buf_1_rs1_paddr ? io_avail_list_57 : _GEN_184; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_186 = 6'h3a == buf_1_rs1_paddr ? io_avail_list_58 : _GEN_185; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_187 = 6'h3b == buf_1_rs1_paddr ? io_avail_list_59 : _GEN_186; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_188 = 6'h3c == buf_1_rs1_paddr ? io_avail_list_60 : _GEN_187; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_189 = 6'h3d == buf_1_rs1_paddr ? io_avail_list_61 : _GEN_188; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_190 = 6'h3e == buf_1_rs1_paddr ? io_avail_list_62 : _GEN_189; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_191 = 6'h3f == buf_1_rs1_paddr ? io_avail_list_63 : _GEN_190; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_193 = 6'h1 == buf_1_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_194 = 6'h2 == buf_1_rs2_paddr ? io_avail_list_2 : _GEN_193; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_195 = 6'h3 == buf_1_rs2_paddr ? io_avail_list_3 : _GEN_194; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_196 = 6'h4 == buf_1_rs2_paddr ? io_avail_list_4 : _GEN_195; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_197 = 6'h5 == buf_1_rs2_paddr ? io_avail_list_5 : _GEN_196; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_198 = 6'h6 == buf_1_rs2_paddr ? io_avail_list_6 : _GEN_197; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_199 = 6'h7 == buf_1_rs2_paddr ? io_avail_list_7 : _GEN_198; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_200 = 6'h8 == buf_1_rs2_paddr ? io_avail_list_8 : _GEN_199; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_201 = 6'h9 == buf_1_rs2_paddr ? io_avail_list_9 : _GEN_200; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_202 = 6'ha == buf_1_rs2_paddr ? io_avail_list_10 : _GEN_201; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_203 = 6'hb == buf_1_rs2_paddr ? io_avail_list_11 : _GEN_202; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_204 = 6'hc == buf_1_rs2_paddr ? io_avail_list_12 : _GEN_203; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_205 = 6'hd == buf_1_rs2_paddr ? io_avail_list_13 : _GEN_204; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_206 = 6'he == buf_1_rs2_paddr ? io_avail_list_14 : _GEN_205; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_207 = 6'hf == buf_1_rs2_paddr ? io_avail_list_15 : _GEN_206; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_208 = 6'h10 == buf_1_rs2_paddr ? io_avail_list_16 : _GEN_207; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_209 = 6'h11 == buf_1_rs2_paddr ? io_avail_list_17 : _GEN_208; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_210 = 6'h12 == buf_1_rs2_paddr ? io_avail_list_18 : _GEN_209; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_211 = 6'h13 == buf_1_rs2_paddr ? io_avail_list_19 : _GEN_210; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_212 = 6'h14 == buf_1_rs2_paddr ? io_avail_list_20 : _GEN_211; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_213 = 6'h15 == buf_1_rs2_paddr ? io_avail_list_21 : _GEN_212; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_214 = 6'h16 == buf_1_rs2_paddr ? io_avail_list_22 : _GEN_213; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_215 = 6'h17 == buf_1_rs2_paddr ? io_avail_list_23 : _GEN_214; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_216 = 6'h18 == buf_1_rs2_paddr ? io_avail_list_24 : _GEN_215; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_217 = 6'h19 == buf_1_rs2_paddr ? io_avail_list_25 : _GEN_216; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_218 = 6'h1a == buf_1_rs2_paddr ? io_avail_list_26 : _GEN_217; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_219 = 6'h1b == buf_1_rs2_paddr ? io_avail_list_27 : _GEN_218; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_220 = 6'h1c == buf_1_rs2_paddr ? io_avail_list_28 : _GEN_219; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_221 = 6'h1d == buf_1_rs2_paddr ? io_avail_list_29 : _GEN_220; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_222 = 6'h1e == buf_1_rs2_paddr ? io_avail_list_30 : _GEN_221; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_223 = 6'h1f == buf_1_rs2_paddr ? io_avail_list_31 : _GEN_222; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_224 = 6'h20 == buf_1_rs2_paddr ? io_avail_list_32 : _GEN_223; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_225 = 6'h21 == buf_1_rs2_paddr ? io_avail_list_33 : _GEN_224; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_226 = 6'h22 == buf_1_rs2_paddr ? io_avail_list_34 : _GEN_225; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_227 = 6'h23 == buf_1_rs2_paddr ? io_avail_list_35 : _GEN_226; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_228 = 6'h24 == buf_1_rs2_paddr ? io_avail_list_36 : _GEN_227; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_229 = 6'h25 == buf_1_rs2_paddr ? io_avail_list_37 : _GEN_228; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_230 = 6'h26 == buf_1_rs2_paddr ? io_avail_list_38 : _GEN_229; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_231 = 6'h27 == buf_1_rs2_paddr ? io_avail_list_39 : _GEN_230; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_232 = 6'h28 == buf_1_rs2_paddr ? io_avail_list_40 : _GEN_231; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_233 = 6'h29 == buf_1_rs2_paddr ? io_avail_list_41 : _GEN_232; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_234 = 6'h2a == buf_1_rs2_paddr ? io_avail_list_42 : _GEN_233; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_235 = 6'h2b == buf_1_rs2_paddr ? io_avail_list_43 : _GEN_234; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_236 = 6'h2c == buf_1_rs2_paddr ? io_avail_list_44 : _GEN_235; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_237 = 6'h2d == buf_1_rs2_paddr ? io_avail_list_45 : _GEN_236; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_238 = 6'h2e == buf_1_rs2_paddr ? io_avail_list_46 : _GEN_237; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_239 = 6'h2f == buf_1_rs2_paddr ? io_avail_list_47 : _GEN_238; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_240 = 6'h30 == buf_1_rs2_paddr ? io_avail_list_48 : _GEN_239; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_241 = 6'h31 == buf_1_rs2_paddr ? io_avail_list_49 : _GEN_240; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_242 = 6'h32 == buf_1_rs2_paddr ? io_avail_list_50 : _GEN_241; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_243 = 6'h33 == buf_1_rs2_paddr ? io_avail_list_51 : _GEN_242; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_244 = 6'h34 == buf_1_rs2_paddr ? io_avail_list_52 : _GEN_243; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_245 = 6'h35 == buf_1_rs2_paddr ? io_avail_list_53 : _GEN_244; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_246 = 6'h36 == buf_1_rs2_paddr ? io_avail_list_54 : _GEN_245; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_247 = 6'h37 == buf_1_rs2_paddr ? io_avail_list_55 : _GEN_246; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_248 = 6'h38 == buf_1_rs2_paddr ? io_avail_list_56 : _GEN_247; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_249 = 6'h39 == buf_1_rs2_paddr ? io_avail_list_57 : _GEN_248; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_250 = 6'h3a == buf_1_rs2_paddr ? io_avail_list_58 : _GEN_249; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_251 = 6'h3b == buf_1_rs2_paddr ? io_avail_list_59 : _GEN_250; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_252 = 6'h3c == buf_1_rs2_paddr ? io_avail_list_60 : _GEN_251; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_253 = 6'h3d == buf_1_rs2_paddr ? io_avail_list_61 : _GEN_252; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_254 = 6'h3e == buf_1_rs2_paddr ? io_avail_list_62 : _GEN_253; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_255 = 6'h3f == buf_1_rs2_paddr ? io_avail_list_63 : _GEN_254; // @[IssueUnit.scala 133:{34,34}]
  wire  ready_list_1 = _GEN_191 & _GEN_255 & ~is_sys_1; // @[IssueUnit.scala 133:59]
  wire  _GEN_257 = 6'h1 == buf_2_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_258 = 6'h2 == buf_2_rs1_paddr ? io_avail_list_2 : _GEN_257; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_259 = 6'h3 == buf_2_rs1_paddr ? io_avail_list_3 : _GEN_258; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_260 = 6'h4 == buf_2_rs1_paddr ? io_avail_list_4 : _GEN_259; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_261 = 6'h5 == buf_2_rs1_paddr ? io_avail_list_5 : _GEN_260; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_262 = 6'h6 == buf_2_rs1_paddr ? io_avail_list_6 : _GEN_261; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_263 = 6'h7 == buf_2_rs1_paddr ? io_avail_list_7 : _GEN_262; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_264 = 6'h8 == buf_2_rs1_paddr ? io_avail_list_8 : _GEN_263; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_265 = 6'h9 == buf_2_rs1_paddr ? io_avail_list_9 : _GEN_264; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_266 = 6'ha == buf_2_rs1_paddr ? io_avail_list_10 : _GEN_265; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_267 = 6'hb == buf_2_rs1_paddr ? io_avail_list_11 : _GEN_266; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_268 = 6'hc == buf_2_rs1_paddr ? io_avail_list_12 : _GEN_267; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_269 = 6'hd == buf_2_rs1_paddr ? io_avail_list_13 : _GEN_268; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_270 = 6'he == buf_2_rs1_paddr ? io_avail_list_14 : _GEN_269; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_271 = 6'hf == buf_2_rs1_paddr ? io_avail_list_15 : _GEN_270; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_272 = 6'h10 == buf_2_rs1_paddr ? io_avail_list_16 : _GEN_271; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_273 = 6'h11 == buf_2_rs1_paddr ? io_avail_list_17 : _GEN_272; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_274 = 6'h12 == buf_2_rs1_paddr ? io_avail_list_18 : _GEN_273; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_275 = 6'h13 == buf_2_rs1_paddr ? io_avail_list_19 : _GEN_274; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_276 = 6'h14 == buf_2_rs1_paddr ? io_avail_list_20 : _GEN_275; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_277 = 6'h15 == buf_2_rs1_paddr ? io_avail_list_21 : _GEN_276; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_278 = 6'h16 == buf_2_rs1_paddr ? io_avail_list_22 : _GEN_277; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_279 = 6'h17 == buf_2_rs1_paddr ? io_avail_list_23 : _GEN_278; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_280 = 6'h18 == buf_2_rs1_paddr ? io_avail_list_24 : _GEN_279; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_281 = 6'h19 == buf_2_rs1_paddr ? io_avail_list_25 : _GEN_280; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_282 = 6'h1a == buf_2_rs1_paddr ? io_avail_list_26 : _GEN_281; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_283 = 6'h1b == buf_2_rs1_paddr ? io_avail_list_27 : _GEN_282; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_284 = 6'h1c == buf_2_rs1_paddr ? io_avail_list_28 : _GEN_283; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_285 = 6'h1d == buf_2_rs1_paddr ? io_avail_list_29 : _GEN_284; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_286 = 6'h1e == buf_2_rs1_paddr ? io_avail_list_30 : _GEN_285; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_287 = 6'h1f == buf_2_rs1_paddr ? io_avail_list_31 : _GEN_286; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_288 = 6'h20 == buf_2_rs1_paddr ? io_avail_list_32 : _GEN_287; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_289 = 6'h21 == buf_2_rs1_paddr ? io_avail_list_33 : _GEN_288; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_290 = 6'h22 == buf_2_rs1_paddr ? io_avail_list_34 : _GEN_289; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_291 = 6'h23 == buf_2_rs1_paddr ? io_avail_list_35 : _GEN_290; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_292 = 6'h24 == buf_2_rs1_paddr ? io_avail_list_36 : _GEN_291; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_293 = 6'h25 == buf_2_rs1_paddr ? io_avail_list_37 : _GEN_292; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_294 = 6'h26 == buf_2_rs1_paddr ? io_avail_list_38 : _GEN_293; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_295 = 6'h27 == buf_2_rs1_paddr ? io_avail_list_39 : _GEN_294; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_296 = 6'h28 == buf_2_rs1_paddr ? io_avail_list_40 : _GEN_295; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_297 = 6'h29 == buf_2_rs1_paddr ? io_avail_list_41 : _GEN_296; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_298 = 6'h2a == buf_2_rs1_paddr ? io_avail_list_42 : _GEN_297; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_299 = 6'h2b == buf_2_rs1_paddr ? io_avail_list_43 : _GEN_298; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_300 = 6'h2c == buf_2_rs1_paddr ? io_avail_list_44 : _GEN_299; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_301 = 6'h2d == buf_2_rs1_paddr ? io_avail_list_45 : _GEN_300; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_302 = 6'h2e == buf_2_rs1_paddr ? io_avail_list_46 : _GEN_301; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_303 = 6'h2f == buf_2_rs1_paddr ? io_avail_list_47 : _GEN_302; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_304 = 6'h30 == buf_2_rs1_paddr ? io_avail_list_48 : _GEN_303; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_305 = 6'h31 == buf_2_rs1_paddr ? io_avail_list_49 : _GEN_304; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_306 = 6'h32 == buf_2_rs1_paddr ? io_avail_list_50 : _GEN_305; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_307 = 6'h33 == buf_2_rs1_paddr ? io_avail_list_51 : _GEN_306; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_308 = 6'h34 == buf_2_rs1_paddr ? io_avail_list_52 : _GEN_307; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_309 = 6'h35 == buf_2_rs1_paddr ? io_avail_list_53 : _GEN_308; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_310 = 6'h36 == buf_2_rs1_paddr ? io_avail_list_54 : _GEN_309; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_311 = 6'h37 == buf_2_rs1_paddr ? io_avail_list_55 : _GEN_310; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_312 = 6'h38 == buf_2_rs1_paddr ? io_avail_list_56 : _GEN_311; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_313 = 6'h39 == buf_2_rs1_paddr ? io_avail_list_57 : _GEN_312; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_314 = 6'h3a == buf_2_rs1_paddr ? io_avail_list_58 : _GEN_313; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_315 = 6'h3b == buf_2_rs1_paddr ? io_avail_list_59 : _GEN_314; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_316 = 6'h3c == buf_2_rs1_paddr ? io_avail_list_60 : _GEN_315; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_317 = 6'h3d == buf_2_rs1_paddr ? io_avail_list_61 : _GEN_316; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_318 = 6'h3e == buf_2_rs1_paddr ? io_avail_list_62 : _GEN_317; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_319 = 6'h3f == buf_2_rs1_paddr ? io_avail_list_63 : _GEN_318; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_321 = 6'h1 == buf_2_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_322 = 6'h2 == buf_2_rs2_paddr ? io_avail_list_2 : _GEN_321; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_323 = 6'h3 == buf_2_rs2_paddr ? io_avail_list_3 : _GEN_322; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_324 = 6'h4 == buf_2_rs2_paddr ? io_avail_list_4 : _GEN_323; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_325 = 6'h5 == buf_2_rs2_paddr ? io_avail_list_5 : _GEN_324; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_326 = 6'h6 == buf_2_rs2_paddr ? io_avail_list_6 : _GEN_325; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_327 = 6'h7 == buf_2_rs2_paddr ? io_avail_list_7 : _GEN_326; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_328 = 6'h8 == buf_2_rs2_paddr ? io_avail_list_8 : _GEN_327; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_329 = 6'h9 == buf_2_rs2_paddr ? io_avail_list_9 : _GEN_328; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_330 = 6'ha == buf_2_rs2_paddr ? io_avail_list_10 : _GEN_329; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_331 = 6'hb == buf_2_rs2_paddr ? io_avail_list_11 : _GEN_330; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_332 = 6'hc == buf_2_rs2_paddr ? io_avail_list_12 : _GEN_331; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_333 = 6'hd == buf_2_rs2_paddr ? io_avail_list_13 : _GEN_332; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_334 = 6'he == buf_2_rs2_paddr ? io_avail_list_14 : _GEN_333; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_335 = 6'hf == buf_2_rs2_paddr ? io_avail_list_15 : _GEN_334; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_336 = 6'h10 == buf_2_rs2_paddr ? io_avail_list_16 : _GEN_335; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_337 = 6'h11 == buf_2_rs2_paddr ? io_avail_list_17 : _GEN_336; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_338 = 6'h12 == buf_2_rs2_paddr ? io_avail_list_18 : _GEN_337; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_339 = 6'h13 == buf_2_rs2_paddr ? io_avail_list_19 : _GEN_338; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_340 = 6'h14 == buf_2_rs2_paddr ? io_avail_list_20 : _GEN_339; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_341 = 6'h15 == buf_2_rs2_paddr ? io_avail_list_21 : _GEN_340; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_342 = 6'h16 == buf_2_rs2_paddr ? io_avail_list_22 : _GEN_341; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_343 = 6'h17 == buf_2_rs2_paddr ? io_avail_list_23 : _GEN_342; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_344 = 6'h18 == buf_2_rs2_paddr ? io_avail_list_24 : _GEN_343; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_345 = 6'h19 == buf_2_rs2_paddr ? io_avail_list_25 : _GEN_344; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_346 = 6'h1a == buf_2_rs2_paddr ? io_avail_list_26 : _GEN_345; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_347 = 6'h1b == buf_2_rs2_paddr ? io_avail_list_27 : _GEN_346; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_348 = 6'h1c == buf_2_rs2_paddr ? io_avail_list_28 : _GEN_347; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_349 = 6'h1d == buf_2_rs2_paddr ? io_avail_list_29 : _GEN_348; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_350 = 6'h1e == buf_2_rs2_paddr ? io_avail_list_30 : _GEN_349; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_351 = 6'h1f == buf_2_rs2_paddr ? io_avail_list_31 : _GEN_350; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_352 = 6'h20 == buf_2_rs2_paddr ? io_avail_list_32 : _GEN_351; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_353 = 6'h21 == buf_2_rs2_paddr ? io_avail_list_33 : _GEN_352; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_354 = 6'h22 == buf_2_rs2_paddr ? io_avail_list_34 : _GEN_353; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_355 = 6'h23 == buf_2_rs2_paddr ? io_avail_list_35 : _GEN_354; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_356 = 6'h24 == buf_2_rs2_paddr ? io_avail_list_36 : _GEN_355; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_357 = 6'h25 == buf_2_rs2_paddr ? io_avail_list_37 : _GEN_356; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_358 = 6'h26 == buf_2_rs2_paddr ? io_avail_list_38 : _GEN_357; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_359 = 6'h27 == buf_2_rs2_paddr ? io_avail_list_39 : _GEN_358; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_360 = 6'h28 == buf_2_rs2_paddr ? io_avail_list_40 : _GEN_359; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_361 = 6'h29 == buf_2_rs2_paddr ? io_avail_list_41 : _GEN_360; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_362 = 6'h2a == buf_2_rs2_paddr ? io_avail_list_42 : _GEN_361; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_363 = 6'h2b == buf_2_rs2_paddr ? io_avail_list_43 : _GEN_362; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_364 = 6'h2c == buf_2_rs2_paddr ? io_avail_list_44 : _GEN_363; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_365 = 6'h2d == buf_2_rs2_paddr ? io_avail_list_45 : _GEN_364; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_366 = 6'h2e == buf_2_rs2_paddr ? io_avail_list_46 : _GEN_365; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_367 = 6'h2f == buf_2_rs2_paddr ? io_avail_list_47 : _GEN_366; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_368 = 6'h30 == buf_2_rs2_paddr ? io_avail_list_48 : _GEN_367; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_369 = 6'h31 == buf_2_rs2_paddr ? io_avail_list_49 : _GEN_368; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_370 = 6'h32 == buf_2_rs2_paddr ? io_avail_list_50 : _GEN_369; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_371 = 6'h33 == buf_2_rs2_paddr ? io_avail_list_51 : _GEN_370; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_372 = 6'h34 == buf_2_rs2_paddr ? io_avail_list_52 : _GEN_371; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_373 = 6'h35 == buf_2_rs2_paddr ? io_avail_list_53 : _GEN_372; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_374 = 6'h36 == buf_2_rs2_paddr ? io_avail_list_54 : _GEN_373; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_375 = 6'h37 == buf_2_rs2_paddr ? io_avail_list_55 : _GEN_374; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_376 = 6'h38 == buf_2_rs2_paddr ? io_avail_list_56 : _GEN_375; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_377 = 6'h39 == buf_2_rs2_paddr ? io_avail_list_57 : _GEN_376; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_378 = 6'h3a == buf_2_rs2_paddr ? io_avail_list_58 : _GEN_377; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_379 = 6'h3b == buf_2_rs2_paddr ? io_avail_list_59 : _GEN_378; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_380 = 6'h3c == buf_2_rs2_paddr ? io_avail_list_60 : _GEN_379; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_381 = 6'h3d == buf_2_rs2_paddr ? io_avail_list_61 : _GEN_380; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_382 = 6'h3e == buf_2_rs2_paddr ? io_avail_list_62 : _GEN_381; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_383 = 6'h3f == buf_2_rs2_paddr ? io_avail_list_63 : _GEN_382; // @[IssueUnit.scala 133:{34,34}]
  wire  ready_list_2 = _GEN_319 & _GEN_383 & ~is_sys_2; // @[IssueUnit.scala 133:59]
  wire  _GEN_385 = 6'h1 == buf_3_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_386 = 6'h2 == buf_3_rs1_paddr ? io_avail_list_2 : _GEN_385; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_387 = 6'h3 == buf_3_rs1_paddr ? io_avail_list_3 : _GEN_386; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_388 = 6'h4 == buf_3_rs1_paddr ? io_avail_list_4 : _GEN_387; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_389 = 6'h5 == buf_3_rs1_paddr ? io_avail_list_5 : _GEN_388; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_390 = 6'h6 == buf_3_rs1_paddr ? io_avail_list_6 : _GEN_389; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_391 = 6'h7 == buf_3_rs1_paddr ? io_avail_list_7 : _GEN_390; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_392 = 6'h8 == buf_3_rs1_paddr ? io_avail_list_8 : _GEN_391; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_393 = 6'h9 == buf_3_rs1_paddr ? io_avail_list_9 : _GEN_392; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_394 = 6'ha == buf_3_rs1_paddr ? io_avail_list_10 : _GEN_393; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_395 = 6'hb == buf_3_rs1_paddr ? io_avail_list_11 : _GEN_394; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_396 = 6'hc == buf_3_rs1_paddr ? io_avail_list_12 : _GEN_395; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_397 = 6'hd == buf_3_rs1_paddr ? io_avail_list_13 : _GEN_396; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_398 = 6'he == buf_3_rs1_paddr ? io_avail_list_14 : _GEN_397; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_399 = 6'hf == buf_3_rs1_paddr ? io_avail_list_15 : _GEN_398; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_400 = 6'h10 == buf_3_rs1_paddr ? io_avail_list_16 : _GEN_399; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_401 = 6'h11 == buf_3_rs1_paddr ? io_avail_list_17 : _GEN_400; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_402 = 6'h12 == buf_3_rs1_paddr ? io_avail_list_18 : _GEN_401; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_403 = 6'h13 == buf_3_rs1_paddr ? io_avail_list_19 : _GEN_402; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_404 = 6'h14 == buf_3_rs1_paddr ? io_avail_list_20 : _GEN_403; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_405 = 6'h15 == buf_3_rs1_paddr ? io_avail_list_21 : _GEN_404; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_406 = 6'h16 == buf_3_rs1_paddr ? io_avail_list_22 : _GEN_405; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_407 = 6'h17 == buf_3_rs1_paddr ? io_avail_list_23 : _GEN_406; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_408 = 6'h18 == buf_3_rs1_paddr ? io_avail_list_24 : _GEN_407; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_409 = 6'h19 == buf_3_rs1_paddr ? io_avail_list_25 : _GEN_408; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_410 = 6'h1a == buf_3_rs1_paddr ? io_avail_list_26 : _GEN_409; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_411 = 6'h1b == buf_3_rs1_paddr ? io_avail_list_27 : _GEN_410; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_412 = 6'h1c == buf_3_rs1_paddr ? io_avail_list_28 : _GEN_411; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_413 = 6'h1d == buf_3_rs1_paddr ? io_avail_list_29 : _GEN_412; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_414 = 6'h1e == buf_3_rs1_paddr ? io_avail_list_30 : _GEN_413; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_415 = 6'h1f == buf_3_rs1_paddr ? io_avail_list_31 : _GEN_414; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_416 = 6'h20 == buf_3_rs1_paddr ? io_avail_list_32 : _GEN_415; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_417 = 6'h21 == buf_3_rs1_paddr ? io_avail_list_33 : _GEN_416; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_418 = 6'h22 == buf_3_rs1_paddr ? io_avail_list_34 : _GEN_417; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_419 = 6'h23 == buf_3_rs1_paddr ? io_avail_list_35 : _GEN_418; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_420 = 6'h24 == buf_3_rs1_paddr ? io_avail_list_36 : _GEN_419; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_421 = 6'h25 == buf_3_rs1_paddr ? io_avail_list_37 : _GEN_420; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_422 = 6'h26 == buf_3_rs1_paddr ? io_avail_list_38 : _GEN_421; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_423 = 6'h27 == buf_3_rs1_paddr ? io_avail_list_39 : _GEN_422; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_424 = 6'h28 == buf_3_rs1_paddr ? io_avail_list_40 : _GEN_423; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_425 = 6'h29 == buf_3_rs1_paddr ? io_avail_list_41 : _GEN_424; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_426 = 6'h2a == buf_3_rs1_paddr ? io_avail_list_42 : _GEN_425; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_427 = 6'h2b == buf_3_rs1_paddr ? io_avail_list_43 : _GEN_426; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_428 = 6'h2c == buf_3_rs1_paddr ? io_avail_list_44 : _GEN_427; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_429 = 6'h2d == buf_3_rs1_paddr ? io_avail_list_45 : _GEN_428; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_430 = 6'h2e == buf_3_rs1_paddr ? io_avail_list_46 : _GEN_429; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_431 = 6'h2f == buf_3_rs1_paddr ? io_avail_list_47 : _GEN_430; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_432 = 6'h30 == buf_3_rs1_paddr ? io_avail_list_48 : _GEN_431; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_433 = 6'h31 == buf_3_rs1_paddr ? io_avail_list_49 : _GEN_432; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_434 = 6'h32 == buf_3_rs1_paddr ? io_avail_list_50 : _GEN_433; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_435 = 6'h33 == buf_3_rs1_paddr ? io_avail_list_51 : _GEN_434; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_436 = 6'h34 == buf_3_rs1_paddr ? io_avail_list_52 : _GEN_435; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_437 = 6'h35 == buf_3_rs1_paddr ? io_avail_list_53 : _GEN_436; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_438 = 6'h36 == buf_3_rs1_paddr ? io_avail_list_54 : _GEN_437; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_439 = 6'h37 == buf_3_rs1_paddr ? io_avail_list_55 : _GEN_438; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_440 = 6'h38 == buf_3_rs1_paddr ? io_avail_list_56 : _GEN_439; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_441 = 6'h39 == buf_3_rs1_paddr ? io_avail_list_57 : _GEN_440; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_442 = 6'h3a == buf_3_rs1_paddr ? io_avail_list_58 : _GEN_441; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_443 = 6'h3b == buf_3_rs1_paddr ? io_avail_list_59 : _GEN_442; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_444 = 6'h3c == buf_3_rs1_paddr ? io_avail_list_60 : _GEN_443; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_445 = 6'h3d == buf_3_rs1_paddr ? io_avail_list_61 : _GEN_444; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_446 = 6'h3e == buf_3_rs1_paddr ? io_avail_list_62 : _GEN_445; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_447 = 6'h3f == buf_3_rs1_paddr ? io_avail_list_63 : _GEN_446; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_449 = 6'h1 == buf_3_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_450 = 6'h2 == buf_3_rs2_paddr ? io_avail_list_2 : _GEN_449; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_451 = 6'h3 == buf_3_rs2_paddr ? io_avail_list_3 : _GEN_450; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_452 = 6'h4 == buf_3_rs2_paddr ? io_avail_list_4 : _GEN_451; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_453 = 6'h5 == buf_3_rs2_paddr ? io_avail_list_5 : _GEN_452; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_454 = 6'h6 == buf_3_rs2_paddr ? io_avail_list_6 : _GEN_453; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_455 = 6'h7 == buf_3_rs2_paddr ? io_avail_list_7 : _GEN_454; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_456 = 6'h8 == buf_3_rs2_paddr ? io_avail_list_8 : _GEN_455; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_457 = 6'h9 == buf_3_rs2_paddr ? io_avail_list_9 : _GEN_456; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_458 = 6'ha == buf_3_rs2_paddr ? io_avail_list_10 : _GEN_457; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_459 = 6'hb == buf_3_rs2_paddr ? io_avail_list_11 : _GEN_458; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_460 = 6'hc == buf_3_rs2_paddr ? io_avail_list_12 : _GEN_459; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_461 = 6'hd == buf_3_rs2_paddr ? io_avail_list_13 : _GEN_460; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_462 = 6'he == buf_3_rs2_paddr ? io_avail_list_14 : _GEN_461; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_463 = 6'hf == buf_3_rs2_paddr ? io_avail_list_15 : _GEN_462; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_464 = 6'h10 == buf_3_rs2_paddr ? io_avail_list_16 : _GEN_463; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_465 = 6'h11 == buf_3_rs2_paddr ? io_avail_list_17 : _GEN_464; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_466 = 6'h12 == buf_3_rs2_paddr ? io_avail_list_18 : _GEN_465; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_467 = 6'h13 == buf_3_rs2_paddr ? io_avail_list_19 : _GEN_466; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_468 = 6'h14 == buf_3_rs2_paddr ? io_avail_list_20 : _GEN_467; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_469 = 6'h15 == buf_3_rs2_paddr ? io_avail_list_21 : _GEN_468; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_470 = 6'h16 == buf_3_rs2_paddr ? io_avail_list_22 : _GEN_469; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_471 = 6'h17 == buf_3_rs2_paddr ? io_avail_list_23 : _GEN_470; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_472 = 6'h18 == buf_3_rs2_paddr ? io_avail_list_24 : _GEN_471; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_473 = 6'h19 == buf_3_rs2_paddr ? io_avail_list_25 : _GEN_472; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_474 = 6'h1a == buf_3_rs2_paddr ? io_avail_list_26 : _GEN_473; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_475 = 6'h1b == buf_3_rs2_paddr ? io_avail_list_27 : _GEN_474; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_476 = 6'h1c == buf_3_rs2_paddr ? io_avail_list_28 : _GEN_475; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_477 = 6'h1d == buf_3_rs2_paddr ? io_avail_list_29 : _GEN_476; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_478 = 6'h1e == buf_3_rs2_paddr ? io_avail_list_30 : _GEN_477; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_479 = 6'h1f == buf_3_rs2_paddr ? io_avail_list_31 : _GEN_478; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_480 = 6'h20 == buf_3_rs2_paddr ? io_avail_list_32 : _GEN_479; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_481 = 6'h21 == buf_3_rs2_paddr ? io_avail_list_33 : _GEN_480; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_482 = 6'h22 == buf_3_rs2_paddr ? io_avail_list_34 : _GEN_481; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_483 = 6'h23 == buf_3_rs2_paddr ? io_avail_list_35 : _GEN_482; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_484 = 6'h24 == buf_3_rs2_paddr ? io_avail_list_36 : _GEN_483; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_485 = 6'h25 == buf_3_rs2_paddr ? io_avail_list_37 : _GEN_484; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_486 = 6'h26 == buf_3_rs2_paddr ? io_avail_list_38 : _GEN_485; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_487 = 6'h27 == buf_3_rs2_paddr ? io_avail_list_39 : _GEN_486; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_488 = 6'h28 == buf_3_rs2_paddr ? io_avail_list_40 : _GEN_487; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_489 = 6'h29 == buf_3_rs2_paddr ? io_avail_list_41 : _GEN_488; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_490 = 6'h2a == buf_3_rs2_paddr ? io_avail_list_42 : _GEN_489; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_491 = 6'h2b == buf_3_rs2_paddr ? io_avail_list_43 : _GEN_490; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_492 = 6'h2c == buf_3_rs2_paddr ? io_avail_list_44 : _GEN_491; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_493 = 6'h2d == buf_3_rs2_paddr ? io_avail_list_45 : _GEN_492; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_494 = 6'h2e == buf_3_rs2_paddr ? io_avail_list_46 : _GEN_493; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_495 = 6'h2f == buf_3_rs2_paddr ? io_avail_list_47 : _GEN_494; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_496 = 6'h30 == buf_3_rs2_paddr ? io_avail_list_48 : _GEN_495; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_497 = 6'h31 == buf_3_rs2_paddr ? io_avail_list_49 : _GEN_496; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_498 = 6'h32 == buf_3_rs2_paddr ? io_avail_list_50 : _GEN_497; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_499 = 6'h33 == buf_3_rs2_paddr ? io_avail_list_51 : _GEN_498; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_500 = 6'h34 == buf_3_rs2_paddr ? io_avail_list_52 : _GEN_499; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_501 = 6'h35 == buf_3_rs2_paddr ? io_avail_list_53 : _GEN_500; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_502 = 6'h36 == buf_3_rs2_paddr ? io_avail_list_54 : _GEN_501; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_503 = 6'h37 == buf_3_rs2_paddr ? io_avail_list_55 : _GEN_502; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_504 = 6'h38 == buf_3_rs2_paddr ? io_avail_list_56 : _GEN_503; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_505 = 6'h39 == buf_3_rs2_paddr ? io_avail_list_57 : _GEN_504; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_506 = 6'h3a == buf_3_rs2_paddr ? io_avail_list_58 : _GEN_505; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_507 = 6'h3b == buf_3_rs2_paddr ? io_avail_list_59 : _GEN_506; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_508 = 6'h3c == buf_3_rs2_paddr ? io_avail_list_60 : _GEN_507; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_509 = 6'h3d == buf_3_rs2_paddr ? io_avail_list_61 : _GEN_508; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_510 = 6'h3e == buf_3_rs2_paddr ? io_avail_list_62 : _GEN_509; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_511 = 6'h3f == buf_3_rs2_paddr ? io_avail_list_63 : _GEN_510; // @[IssueUnit.scala 133:{34,34}]
  wire  ready_list_3 = _GEN_447 & _GEN_511 & ~is_sys_3; // @[IssueUnit.scala 133:59]
  wire  _GEN_513 = 6'h1 == buf_4_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_514 = 6'h2 == buf_4_rs1_paddr ? io_avail_list_2 : _GEN_513; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_515 = 6'h3 == buf_4_rs1_paddr ? io_avail_list_3 : _GEN_514; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_516 = 6'h4 == buf_4_rs1_paddr ? io_avail_list_4 : _GEN_515; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_517 = 6'h5 == buf_4_rs1_paddr ? io_avail_list_5 : _GEN_516; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_518 = 6'h6 == buf_4_rs1_paddr ? io_avail_list_6 : _GEN_517; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_519 = 6'h7 == buf_4_rs1_paddr ? io_avail_list_7 : _GEN_518; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_520 = 6'h8 == buf_4_rs1_paddr ? io_avail_list_8 : _GEN_519; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_521 = 6'h9 == buf_4_rs1_paddr ? io_avail_list_9 : _GEN_520; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_522 = 6'ha == buf_4_rs1_paddr ? io_avail_list_10 : _GEN_521; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_523 = 6'hb == buf_4_rs1_paddr ? io_avail_list_11 : _GEN_522; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_524 = 6'hc == buf_4_rs1_paddr ? io_avail_list_12 : _GEN_523; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_525 = 6'hd == buf_4_rs1_paddr ? io_avail_list_13 : _GEN_524; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_526 = 6'he == buf_4_rs1_paddr ? io_avail_list_14 : _GEN_525; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_527 = 6'hf == buf_4_rs1_paddr ? io_avail_list_15 : _GEN_526; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_528 = 6'h10 == buf_4_rs1_paddr ? io_avail_list_16 : _GEN_527; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_529 = 6'h11 == buf_4_rs1_paddr ? io_avail_list_17 : _GEN_528; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_530 = 6'h12 == buf_4_rs1_paddr ? io_avail_list_18 : _GEN_529; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_531 = 6'h13 == buf_4_rs1_paddr ? io_avail_list_19 : _GEN_530; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_532 = 6'h14 == buf_4_rs1_paddr ? io_avail_list_20 : _GEN_531; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_533 = 6'h15 == buf_4_rs1_paddr ? io_avail_list_21 : _GEN_532; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_534 = 6'h16 == buf_4_rs1_paddr ? io_avail_list_22 : _GEN_533; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_535 = 6'h17 == buf_4_rs1_paddr ? io_avail_list_23 : _GEN_534; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_536 = 6'h18 == buf_4_rs1_paddr ? io_avail_list_24 : _GEN_535; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_537 = 6'h19 == buf_4_rs1_paddr ? io_avail_list_25 : _GEN_536; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_538 = 6'h1a == buf_4_rs1_paddr ? io_avail_list_26 : _GEN_537; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_539 = 6'h1b == buf_4_rs1_paddr ? io_avail_list_27 : _GEN_538; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_540 = 6'h1c == buf_4_rs1_paddr ? io_avail_list_28 : _GEN_539; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_541 = 6'h1d == buf_4_rs1_paddr ? io_avail_list_29 : _GEN_540; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_542 = 6'h1e == buf_4_rs1_paddr ? io_avail_list_30 : _GEN_541; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_543 = 6'h1f == buf_4_rs1_paddr ? io_avail_list_31 : _GEN_542; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_544 = 6'h20 == buf_4_rs1_paddr ? io_avail_list_32 : _GEN_543; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_545 = 6'h21 == buf_4_rs1_paddr ? io_avail_list_33 : _GEN_544; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_546 = 6'h22 == buf_4_rs1_paddr ? io_avail_list_34 : _GEN_545; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_547 = 6'h23 == buf_4_rs1_paddr ? io_avail_list_35 : _GEN_546; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_548 = 6'h24 == buf_4_rs1_paddr ? io_avail_list_36 : _GEN_547; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_549 = 6'h25 == buf_4_rs1_paddr ? io_avail_list_37 : _GEN_548; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_550 = 6'h26 == buf_4_rs1_paddr ? io_avail_list_38 : _GEN_549; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_551 = 6'h27 == buf_4_rs1_paddr ? io_avail_list_39 : _GEN_550; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_552 = 6'h28 == buf_4_rs1_paddr ? io_avail_list_40 : _GEN_551; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_553 = 6'h29 == buf_4_rs1_paddr ? io_avail_list_41 : _GEN_552; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_554 = 6'h2a == buf_4_rs1_paddr ? io_avail_list_42 : _GEN_553; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_555 = 6'h2b == buf_4_rs1_paddr ? io_avail_list_43 : _GEN_554; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_556 = 6'h2c == buf_4_rs1_paddr ? io_avail_list_44 : _GEN_555; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_557 = 6'h2d == buf_4_rs1_paddr ? io_avail_list_45 : _GEN_556; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_558 = 6'h2e == buf_4_rs1_paddr ? io_avail_list_46 : _GEN_557; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_559 = 6'h2f == buf_4_rs1_paddr ? io_avail_list_47 : _GEN_558; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_560 = 6'h30 == buf_4_rs1_paddr ? io_avail_list_48 : _GEN_559; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_561 = 6'h31 == buf_4_rs1_paddr ? io_avail_list_49 : _GEN_560; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_562 = 6'h32 == buf_4_rs1_paddr ? io_avail_list_50 : _GEN_561; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_563 = 6'h33 == buf_4_rs1_paddr ? io_avail_list_51 : _GEN_562; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_564 = 6'h34 == buf_4_rs1_paddr ? io_avail_list_52 : _GEN_563; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_565 = 6'h35 == buf_4_rs1_paddr ? io_avail_list_53 : _GEN_564; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_566 = 6'h36 == buf_4_rs1_paddr ? io_avail_list_54 : _GEN_565; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_567 = 6'h37 == buf_4_rs1_paddr ? io_avail_list_55 : _GEN_566; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_568 = 6'h38 == buf_4_rs1_paddr ? io_avail_list_56 : _GEN_567; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_569 = 6'h39 == buf_4_rs1_paddr ? io_avail_list_57 : _GEN_568; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_570 = 6'h3a == buf_4_rs1_paddr ? io_avail_list_58 : _GEN_569; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_571 = 6'h3b == buf_4_rs1_paddr ? io_avail_list_59 : _GEN_570; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_572 = 6'h3c == buf_4_rs1_paddr ? io_avail_list_60 : _GEN_571; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_573 = 6'h3d == buf_4_rs1_paddr ? io_avail_list_61 : _GEN_572; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_574 = 6'h3e == buf_4_rs1_paddr ? io_avail_list_62 : _GEN_573; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_575 = 6'h3f == buf_4_rs1_paddr ? io_avail_list_63 : _GEN_574; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_577 = 6'h1 == buf_4_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_578 = 6'h2 == buf_4_rs2_paddr ? io_avail_list_2 : _GEN_577; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_579 = 6'h3 == buf_4_rs2_paddr ? io_avail_list_3 : _GEN_578; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_580 = 6'h4 == buf_4_rs2_paddr ? io_avail_list_4 : _GEN_579; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_581 = 6'h5 == buf_4_rs2_paddr ? io_avail_list_5 : _GEN_580; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_582 = 6'h6 == buf_4_rs2_paddr ? io_avail_list_6 : _GEN_581; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_583 = 6'h7 == buf_4_rs2_paddr ? io_avail_list_7 : _GEN_582; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_584 = 6'h8 == buf_4_rs2_paddr ? io_avail_list_8 : _GEN_583; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_585 = 6'h9 == buf_4_rs2_paddr ? io_avail_list_9 : _GEN_584; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_586 = 6'ha == buf_4_rs2_paddr ? io_avail_list_10 : _GEN_585; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_587 = 6'hb == buf_4_rs2_paddr ? io_avail_list_11 : _GEN_586; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_588 = 6'hc == buf_4_rs2_paddr ? io_avail_list_12 : _GEN_587; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_589 = 6'hd == buf_4_rs2_paddr ? io_avail_list_13 : _GEN_588; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_590 = 6'he == buf_4_rs2_paddr ? io_avail_list_14 : _GEN_589; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_591 = 6'hf == buf_4_rs2_paddr ? io_avail_list_15 : _GEN_590; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_592 = 6'h10 == buf_4_rs2_paddr ? io_avail_list_16 : _GEN_591; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_593 = 6'h11 == buf_4_rs2_paddr ? io_avail_list_17 : _GEN_592; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_594 = 6'h12 == buf_4_rs2_paddr ? io_avail_list_18 : _GEN_593; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_595 = 6'h13 == buf_4_rs2_paddr ? io_avail_list_19 : _GEN_594; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_596 = 6'h14 == buf_4_rs2_paddr ? io_avail_list_20 : _GEN_595; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_597 = 6'h15 == buf_4_rs2_paddr ? io_avail_list_21 : _GEN_596; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_598 = 6'h16 == buf_4_rs2_paddr ? io_avail_list_22 : _GEN_597; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_599 = 6'h17 == buf_4_rs2_paddr ? io_avail_list_23 : _GEN_598; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_600 = 6'h18 == buf_4_rs2_paddr ? io_avail_list_24 : _GEN_599; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_601 = 6'h19 == buf_4_rs2_paddr ? io_avail_list_25 : _GEN_600; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_602 = 6'h1a == buf_4_rs2_paddr ? io_avail_list_26 : _GEN_601; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_603 = 6'h1b == buf_4_rs2_paddr ? io_avail_list_27 : _GEN_602; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_604 = 6'h1c == buf_4_rs2_paddr ? io_avail_list_28 : _GEN_603; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_605 = 6'h1d == buf_4_rs2_paddr ? io_avail_list_29 : _GEN_604; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_606 = 6'h1e == buf_4_rs2_paddr ? io_avail_list_30 : _GEN_605; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_607 = 6'h1f == buf_4_rs2_paddr ? io_avail_list_31 : _GEN_606; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_608 = 6'h20 == buf_4_rs2_paddr ? io_avail_list_32 : _GEN_607; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_609 = 6'h21 == buf_4_rs2_paddr ? io_avail_list_33 : _GEN_608; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_610 = 6'h22 == buf_4_rs2_paddr ? io_avail_list_34 : _GEN_609; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_611 = 6'h23 == buf_4_rs2_paddr ? io_avail_list_35 : _GEN_610; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_612 = 6'h24 == buf_4_rs2_paddr ? io_avail_list_36 : _GEN_611; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_613 = 6'h25 == buf_4_rs2_paddr ? io_avail_list_37 : _GEN_612; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_614 = 6'h26 == buf_4_rs2_paddr ? io_avail_list_38 : _GEN_613; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_615 = 6'h27 == buf_4_rs2_paddr ? io_avail_list_39 : _GEN_614; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_616 = 6'h28 == buf_4_rs2_paddr ? io_avail_list_40 : _GEN_615; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_617 = 6'h29 == buf_4_rs2_paddr ? io_avail_list_41 : _GEN_616; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_618 = 6'h2a == buf_4_rs2_paddr ? io_avail_list_42 : _GEN_617; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_619 = 6'h2b == buf_4_rs2_paddr ? io_avail_list_43 : _GEN_618; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_620 = 6'h2c == buf_4_rs2_paddr ? io_avail_list_44 : _GEN_619; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_621 = 6'h2d == buf_4_rs2_paddr ? io_avail_list_45 : _GEN_620; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_622 = 6'h2e == buf_4_rs2_paddr ? io_avail_list_46 : _GEN_621; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_623 = 6'h2f == buf_4_rs2_paddr ? io_avail_list_47 : _GEN_622; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_624 = 6'h30 == buf_4_rs2_paddr ? io_avail_list_48 : _GEN_623; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_625 = 6'h31 == buf_4_rs2_paddr ? io_avail_list_49 : _GEN_624; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_626 = 6'h32 == buf_4_rs2_paddr ? io_avail_list_50 : _GEN_625; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_627 = 6'h33 == buf_4_rs2_paddr ? io_avail_list_51 : _GEN_626; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_628 = 6'h34 == buf_4_rs2_paddr ? io_avail_list_52 : _GEN_627; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_629 = 6'h35 == buf_4_rs2_paddr ? io_avail_list_53 : _GEN_628; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_630 = 6'h36 == buf_4_rs2_paddr ? io_avail_list_54 : _GEN_629; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_631 = 6'h37 == buf_4_rs2_paddr ? io_avail_list_55 : _GEN_630; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_632 = 6'h38 == buf_4_rs2_paddr ? io_avail_list_56 : _GEN_631; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_633 = 6'h39 == buf_4_rs2_paddr ? io_avail_list_57 : _GEN_632; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_634 = 6'h3a == buf_4_rs2_paddr ? io_avail_list_58 : _GEN_633; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_635 = 6'h3b == buf_4_rs2_paddr ? io_avail_list_59 : _GEN_634; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_636 = 6'h3c == buf_4_rs2_paddr ? io_avail_list_60 : _GEN_635; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_637 = 6'h3d == buf_4_rs2_paddr ? io_avail_list_61 : _GEN_636; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_638 = 6'h3e == buf_4_rs2_paddr ? io_avail_list_62 : _GEN_637; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_639 = 6'h3f == buf_4_rs2_paddr ? io_avail_list_63 : _GEN_638; // @[IssueUnit.scala 133:{34,34}]
  wire  ready_list_4 = _GEN_575 & _GEN_639 & ~is_sys_4; // @[IssueUnit.scala 133:59]
  wire  _GEN_641 = 6'h1 == buf_5_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_642 = 6'h2 == buf_5_rs1_paddr ? io_avail_list_2 : _GEN_641; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_643 = 6'h3 == buf_5_rs1_paddr ? io_avail_list_3 : _GEN_642; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_644 = 6'h4 == buf_5_rs1_paddr ? io_avail_list_4 : _GEN_643; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_645 = 6'h5 == buf_5_rs1_paddr ? io_avail_list_5 : _GEN_644; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_646 = 6'h6 == buf_5_rs1_paddr ? io_avail_list_6 : _GEN_645; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_647 = 6'h7 == buf_5_rs1_paddr ? io_avail_list_7 : _GEN_646; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_648 = 6'h8 == buf_5_rs1_paddr ? io_avail_list_8 : _GEN_647; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_649 = 6'h9 == buf_5_rs1_paddr ? io_avail_list_9 : _GEN_648; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_650 = 6'ha == buf_5_rs1_paddr ? io_avail_list_10 : _GEN_649; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_651 = 6'hb == buf_5_rs1_paddr ? io_avail_list_11 : _GEN_650; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_652 = 6'hc == buf_5_rs1_paddr ? io_avail_list_12 : _GEN_651; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_653 = 6'hd == buf_5_rs1_paddr ? io_avail_list_13 : _GEN_652; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_654 = 6'he == buf_5_rs1_paddr ? io_avail_list_14 : _GEN_653; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_655 = 6'hf == buf_5_rs1_paddr ? io_avail_list_15 : _GEN_654; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_656 = 6'h10 == buf_5_rs1_paddr ? io_avail_list_16 : _GEN_655; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_657 = 6'h11 == buf_5_rs1_paddr ? io_avail_list_17 : _GEN_656; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_658 = 6'h12 == buf_5_rs1_paddr ? io_avail_list_18 : _GEN_657; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_659 = 6'h13 == buf_5_rs1_paddr ? io_avail_list_19 : _GEN_658; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_660 = 6'h14 == buf_5_rs1_paddr ? io_avail_list_20 : _GEN_659; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_661 = 6'h15 == buf_5_rs1_paddr ? io_avail_list_21 : _GEN_660; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_662 = 6'h16 == buf_5_rs1_paddr ? io_avail_list_22 : _GEN_661; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_663 = 6'h17 == buf_5_rs1_paddr ? io_avail_list_23 : _GEN_662; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_664 = 6'h18 == buf_5_rs1_paddr ? io_avail_list_24 : _GEN_663; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_665 = 6'h19 == buf_5_rs1_paddr ? io_avail_list_25 : _GEN_664; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_666 = 6'h1a == buf_5_rs1_paddr ? io_avail_list_26 : _GEN_665; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_667 = 6'h1b == buf_5_rs1_paddr ? io_avail_list_27 : _GEN_666; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_668 = 6'h1c == buf_5_rs1_paddr ? io_avail_list_28 : _GEN_667; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_669 = 6'h1d == buf_5_rs1_paddr ? io_avail_list_29 : _GEN_668; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_670 = 6'h1e == buf_5_rs1_paddr ? io_avail_list_30 : _GEN_669; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_671 = 6'h1f == buf_5_rs1_paddr ? io_avail_list_31 : _GEN_670; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_672 = 6'h20 == buf_5_rs1_paddr ? io_avail_list_32 : _GEN_671; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_673 = 6'h21 == buf_5_rs1_paddr ? io_avail_list_33 : _GEN_672; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_674 = 6'h22 == buf_5_rs1_paddr ? io_avail_list_34 : _GEN_673; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_675 = 6'h23 == buf_5_rs1_paddr ? io_avail_list_35 : _GEN_674; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_676 = 6'h24 == buf_5_rs1_paddr ? io_avail_list_36 : _GEN_675; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_677 = 6'h25 == buf_5_rs1_paddr ? io_avail_list_37 : _GEN_676; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_678 = 6'h26 == buf_5_rs1_paddr ? io_avail_list_38 : _GEN_677; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_679 = 6'h27 == buf_5_rs1_paddr ? io_avail_list_39 : _GEN_678; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_680 = 6'h28 == buf_5_rs1_paddr ? io_avail_list_40 : _GEN_679; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_681 = 6'h29 == buf_5_rs1_paddr ? io_avail_list_41 : _GEN_680; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_682 = 6'h2a == buf_5_rs1_paddr ? io_avail_list_42 : _GEN_681; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_683 = 6'h2b == buf_5_rs1_paddr ? io_avail_list_43 : _GEN_682; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_684 = 6'h2c == buf_5_rs1_paddr ? io_avail_list_44 : _GEN_683; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_685 = 6'h2d == buf_5_rs1_paddr ? io_avail_list_45 : _GEN_684; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_686 = 6'h2e == buf_5_rs1_paddr ? io_avail_list_46 : _GEN_685; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_687 = 6'h2f == buf_5_rs1_paddr ? io_avail_list_47 : _GEN_686; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_688 = 6'h30 == buf_5_rs1_paddr ? io_avail_list_48 : _GEN_687; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_689 = 6'h31 == buf_5_rs1_paddr ? io_avail_list_49 : _GEN_688; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_690 = 6'h32 == buf_5_rs1_paddr ? io_avail_list_50 : _GEN_689; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_691 = 6'h33 == buf_5_rs1_paddr ? io_avail_list_51 : _GEN_690; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_692 = 6'h34 == buf_5_rs1_paddr ? io_avail_list_52 : _GEN_691; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_693 = 6'h35 == buf_5_rs1_paddr ? io_avail_list_53 : _GEN_692; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_694 = 6'h36 == buf_5_rs1_paddr ? io_avail_list_54 : _GEN_693; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_695 = 6'h37 == buf_5_rs1_paddr ? io_avail_list_55 : _GEN_694; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_696 = 6'h38 == buf_5_rs1_paddr ? io_avail_list_56 : _GEN_695; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_697 = 6'h39 == buf_5_rs1_paddr ? io_avail_list_57 : _GEN_696; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_698 = 6'h3a == buf_5_rs1_paddr ? io_avail_list_58 : _GEN_697; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_699 = 6'h3b == buf_5_rs1_paddr ? io_avail_list_59 : _GEN_698; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_700 = 6'h3c == buf_5_rs1_paddr ? io_avail_list_60 : _GEN_699; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_701 = 6'h3d == buf_5_rs1_paddr ? io_avail_list_61 : _GEN_700; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_702 = 6'h3e == buf_5_rs1_paddr ? io_avail_list_62 : _GEN_701; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_703 = 6'h3f == buf_5_rs1_paddr ? io_avail_list_63 : _GEN_702; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_705 = 6'h1 == buf_5_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_706 = 6'h2 == buf_5_rs2_paddr ? io_avail_list_2 : _GEN_705; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_707 = 6'h3 == buf_5_rs2_paddr ? io_avail_list_3 : _GEN_706; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_708 = 6'h4 == buf_5_rs2_paddr ? io_avail_list_4 : _GEN_707; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_709 = 6'h5 == buf_5_rs2_paddr ? io_avail_list_5 : _GEN_708; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_710 = 6'h6 == buf_5_rs2_paddr ? io_avail_list_6 : _GEN_709; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_711 = 6'h7 == buf_5_rs2_paddr ? io_avail_list_7 : _GEN_710; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_712 = 6'h8 == buf_5_rs2_paddr ? io_avail_list_8 : _GEN_711; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_713 = 6'h9 == buf_5_rs2_paddr ? io_avail_list_9 : _GEN_712; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_714 = 6'ha == buf_5_rs2_paddr ? io_avail_list_10 : _GEN_713; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_715 = 6'hb == buf_5_rs2_paddr ? io_avail_list_11 : _GEN_714; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_716 = 6'hc == buf_5_rs2_paddr ? io_avail_list_12 : _GEN_715; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_717 = 6'hd == buf_5_rs2_paddr ? io_avail_list_13 : _GEN_716; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_718 = 6'he == buf_5_rs2_paddr ? io_avail_list_14 : _GEN_717; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_719 = 6'hf == buf_5_rs2_paddr ? io_avail_list_15 : _GEN_718; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_720 = 6'h10 == buf_5_rs2_paddr ? io_avail_list_16 : _GEN_719; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_721 = 6'h11 == buf_5_rs2_paddr ? io_avail_list_17 : _GEN_720; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_722 = 6'h12 == buf_5_rs2_paddr ? io_avail_list_18 : _GEN_721; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_723 = 6'h13 == buf_5_rs2_paddr ? io_avail_list_19 : _GEN_722; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_724 = 6'h14 == buf_5_rs2_paddr ? io_avail_list_20 : _GEN_723; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_725 = 6'h15 == buf_5_rs2_paddr ? io_avail_list_21 : _GEN_724; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_726 = 6'h16 == buf_5_rs2_paddr ? io_avail_list_22 : _GEN_725; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_727 = 6'h17 == buf_5_rs2_paddr ? io_avail_list_23 : _GEN_726; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_728 = 6'h18 == buf_5_rs2_paddr ? io_avail_list_24 : _GEN_727; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_729 = 6'h19 == buf_5_rs2_paddr ? io_avail_list_25 : _GEN_728; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_730 = 6'h1a == buf_5_rs2_paddr ? io_avail_list_26 : _GEN_729; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_731 = 6'h1b == buf_5_rs2_paddr ? io_avail_list_27 : _GEN_730; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_732 = 6'h1c == buf_5_rs2_paddr ? io_avail_list_28 : _GEN_731; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_733 = 6'h1d == buf_5_rs2_paddr ? io_avail_list_29 : _GEN_732; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_734 = 6'h1e == buf_5_rs2_paddr ? io_avail_list_30 : _GEN_733; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_735 = 6'h1f == buf_5_rs2_paddr ? io_avail_list_31 : _GEN_734; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_736 = 6'h20 == buf_5_rs2_paddr ? io_avail_list_32 : _GEN_735; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_737 = 6'h21 == buf_5_rs2_paddr ? io_avail_list_33 : _GEN_736; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_738 = 6'h22 == buf_5_rs2_paddr ? io_avail_list_34 : _GEN_737; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_739 = 6'h23 == buf_5_rs2_paddr ? io_avail_list_35 : _GEN_738; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_740 = 6'h24 == buf_5_rs2_paddr ? io_avail_list_36 : _GEN_739; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_741 = 6'h25 == buf_5_rs2_paddr ? io_avail_list_37 : _GEN_740; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_742 = 6'h26 == buf_5_rs2_paddr ? io_avail_list_38 : _GEN_741; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_743 = 6'h27 == buf_5_rs2_paddr ? io_avail_list_39 : _GEN_742; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_744 = 6'h28 == buf_5_rs2_paddr ? io_avail_list_40 : _GEN_743; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_745 = 6'h29 == buf_5_rs2_paddr ? io_avail_list_41 : _GEN_744; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_746 = 6'h2a == buf_5_rs2_paddr ? io_avail_list_42 : _GEN_745; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_747 = 6'h2b == buf_5_rs2_paddr ? io_avail_list_43 : _GEN_746; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_748 = 6'h2c == buf_5_rs2_paddr ? io_avail_list_44 : _GEN_747; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_749 = 6'h2d == buf_5_rs2_paddr ? io_avail_list_45 : _GEN_748; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_750 = 6'h2e == buf_5_rs2_paddr ? io_avail_list_46 : _GEN_749; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_751 = 6'h2f == buf_5_rs2_paddr ? io_avail_list_47 : _GEN_750; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_752 = 6'h30 == buf_5_rs2_paddr ? io_avail_list_48 : _GEN_751; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_753 = 6'h31 == buf_5_rs2_paddr ? io_avail_list_49 : _GEN_752; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_754 = 6'h32 == buf_5_rs2_paddr ? io_avail_list_50 : _GEN_753; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_755 = 6'h33 == buf_5_rs2_paddr ? io_avail_list_51 : _GEN_754; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_756 = 6'h34 == buf_5_rs2_paddr ? io_avail_list_52 : _GEN_755; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_757 = 6'h35 == buf_5_rs2_paddr ? io_avail_list_53 : _GEN_756; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_758 = 6'h36 == buf_5_rs2_paddr ? io_avail_list_54 : _GEN_757; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_759 = 6'h37 == buf_5_rs2_paddr ? io_avail_list_55 : _GEN_758; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_760 = 6'h38 == buf_5_rs2_paddr ? io_avail_list_56 : _GEN_759; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_761 = 6'h39 == buf_5_rs2_paddr ? io_avail_list_57 : _GEN_760; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_762 = 6'h3a == buf_5_rs2_paddr ? io_avail_list_58 : _GEN_761; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_763 = 6'h3b == buf_5_rs2_paddr ? io_avail_list_59 : _GEN_762; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_764 = 6'h3c == buf_5_rs2_paddr ? io_avail_list_60 : _GEN_763; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_765 = 6'h3d == buf_5_rs2_paddr ? io_avail_list_61 : _GEN_764; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_766 = 6'h3e == buf_5_rs2_paddr ? io_avail_list_62 : _GEN_765; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_767 = 6'h3f == buf_5_rs2_paddr ? io_avail_list_63 : _GEN_766; // @[IssueUnit.scala 133:{34,34}]
  wire  ready_list_5 = _GEN_703 & _GEN_767 & ~is_sys_5; // @[IssueUnit.scala 133:59]
  wire  _GEN_769 = 6'h1 == buf_6_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_770 = 6'h2 == buf_6_rs1_paddr ? io_avail_list_2 : _GEN_769; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_771 = 6'h3 == buf_6_rs1_paddr ? io_avail_list_3 : _GEN_770; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_772 = 6'h4 == buf_6_rs1_paddr ? io_avail_list_4 : _GEN_771; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_773 = 6'h5 == buf_6_rs1_paddr ? io_avail_list_5 : _GEN_772; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_774 = 6'h6 == buf_6_rs1_paddr ? io_avail_list_6 : _GEN_773; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_775 = 6'h7 == buf_6_rs1_paddr ? io_avail_list_7 : _GEN_774; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_776 = 6'h8 == buf_6_rs1_paddr ? io_avail_list_8 : _GEN_775; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_777 = 6'h9 == buf_6_rs1_paddr ? io_avail_list_9 : _GEN_776; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_778 = 6'ha == buf_6_rs1_paddr ? io_avail_list_10 : _GEN_777; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_779 = 6'hb == buf_6_rs1_paddr ? io_avail_list_11 : _GEN_778; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_780 = 6'hc == buf_6_rs1_paddr ? io_avail_list_12 : _GEN_779; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_781 = 6'hd == buf_6_rs1_paddr ? io_avail_list_13 : _GEN_780; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_782 = 6'he == buf_6_rs1_paddr ? io_avail_list_14 : _GEN_781; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_783 = 6'hf == buf_6_rs1_paddr ? io_avail_list_15 : _GEN_782; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_784 = 6'h10 == buf_6_rs1_paddr ? io_avail_list_16 : _GEN_783; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_785 = 6'h11 == buf_6_rs1_paddr ? io_avail_list_17 : _GEN_784; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_786 = 6'h12 == buf_6_rs1_paddr ? io_avail_list_18 : _GEN_785; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_787 = 6'h13 == buf_6_rs1_paddr ? io_avail_list_19 : _GEN_786; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_788 = 6'h14 == buf_6_rs1_paddr ? io_avail_list_20 : _GEN_787; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_789 = 6'h15 == buf_6_rs1_paddr ? io_avail_list_21 : _GEN_788; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_790 = 6'h16 == buf_6_rs1_paddr ? io_avail_list_22 : _GEN_789; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_791 = 6'h17 == buf_6_rs1_paddr ? io_avail_list_23 : _GEN_790; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_792 = 6'h18 == buf_6_rs1_paddr ? io_avail_list_24 : _GEN_791; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_793 = 6'h19 == buf_6_rs1_paddr ? io_avail_list_25 : _GEN_792; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_794 = 6'h1a == buf_6_rs1_paddr ? io_avail_list_26 : _GEN_793; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_795 = 6'h1b == buf_6_rs1_paddr ? io_avail_list_27 : _GEN_794; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_796 = 6'h1c == buf_6_rs1_paddr ? io_avail_list_28 : _GEN_795; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_797 = 6'h1d == buf_6_rs1_paddr ? io_avail_list_29 : _GEN_796; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_798 = 6'h1e == buf_6_rs1_paddr ? io_avail_list_30 : _GEN_797; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_799 = 6'h1f == buf_6_rs1_paddr ? io_avail_list_31 : _GEN_798; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_800 = 6'h20 == buf_6_rs1_paddr ? io_avail_list_32 : _GEN_799; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_801 = 6'h21 == buf_6_rs1_paddr ? io_avail_list_33 : _GEN_800; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_802 = 6'h22 == buf_6_rs1_paddr ? io_avail_list_34 : _GEN_801; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_803 = 6'h23 == buf_6_rs1_paddr ? io_avail_list_35 : _GEN_802; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_804 = 6'h24 == buf_6_rs1_paddr ? io_avail_list_36 : _GEN_803; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_805 = 6'h25 == buf_6_rs1_paddr ? io_avail_list_37 : _GEN_804; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_806 = 6'h26 == buf_6_rs1_paddr ? io_avail_list_38 : _GEN_805; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_807 = 6'h27 == buf_6_rs1_paddr ? io_avail_list_39 : _GEN_806; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_808 = 6'h28 == buf_6_rs1_paddr ? io_avail_list_40 : _GEN_807; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_809 = 6'h29 == buf_6_rs1_paddr ? io_avail_list_41 : _GEN_808; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_810 = 6'h2a == buf_6_rs1_paddr ? io_avail_list_42 : _GEN_809; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_811 = 6'h2b == buf_6_rs1_paddr ? io_avail_list_43 : _GEN_810; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_812 = 6'h2c == buf_6_rs1_paddr ? io_avail_list_44 : _GEN_811; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_813 = 6'h2d == buf_6_rs1_paddr ? io_avail_list_45 : _GEN_812; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_814 = 6'h2e == buf_6_rs1_paddr ? io_avail_list_46 : _GEN_813; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_815 = 6'h2f == buf_6_rs1_paddr ? io_avail_list_47 : _GEN_814; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_816 = 6'h30 == buf_6_rs1_paddr ? io_avail_list_48 : _GEN_815; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_817 = 6'h31 == buf_6_rs1_paddr ? io_avail_list_49 : _GEN_816; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_818 = 6'h32 == buf_6_rs1_paddr ? io_avail_list_50 : _GEN_817; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_819 = 6'h33 == buf_6_rs1_paddr ? io_avail_list_51 : _GEN_818; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_820 = 6'h34 == buf_6_rs1_paddr ? io_avail_list_52 : _GEN_819; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_821 = 6'h35 == buf_6_rs1_paddr ? io_avail_list_53 : _GEN_820; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_822 = 6'h36 == buf_6_rs1_paddr ? io_avail_list_54 : _GEN_821; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_823 = 6'h37 == buf_6_rs1_paddr ? io_avail_list_55 : _GEN_822; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_824 = 6'h38 == buf_6_rs1_paddr ? io_avail_list_56 : _GEN_823; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_825 = 6'h39 == buf_6_rs1_paddr ? io_avail_list_57 : _GEN_824; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_826 = 6'h3a == buf_6_rs1_paddr ? io_avail_list_58 : _GEN_825; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_827 = 6'h3b == buf_6_rs1_paddr ? io_avail_list_59 : _GEN_826; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_828 = 6'h3c == buf_6_rs1_paddr ? io_avail_list_60 : _GEN_827; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_829 = 6'h3d == buf_6_rs1_paddr ? io_avail_list_61 : _GEN_828; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_830 = 6'h3e == buf_6_rs1_paddr ? io_avail_list_62 : _GEN_829; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_831 = 6'h3f == buf_6_rs1_paddr ? io_avail_list_63 : _GEN_830; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_833 = 6'h1 == buf_6_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_834 = 6'h2 == buf_6_rs2_paddr ? io_avail_list_2 : _GEN_833; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_835 = 6'h3 == buf_6_rs2_paddr ? io_avail_list_3 : _GEN_834; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_836 = 6'h4 == buf_6_rs2_paddr ? io_avail_list_4 : _GEN_835; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_837 = 6'h5 == buf_6_rs2_paddr ? io_avail_list_5 : _GEN_836; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_838 = 6'h6 == buf_6_rs2_paddr ? io_avail_list_6 : _GEN_837; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_839 = 6'h7 == buf_6_rs2_paddr ? io_avail_list_7 : _GEN_838; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_840 = 6'h8 == buf_6_rs2_paddr ? io_avail_list_8 : _GEN_839; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_841 = 6'h9 == buf_6_rs2_paddr ? io_avail_list_9 : _GEN_840; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_842 = 6'ha == buf_6_rs2_paddr ? io_avail_list_10 : _GEN_841; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_843 = 6'hb == buf_6_rs2_paddr ? io_avail_list_11 : _GEN_842; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_844 = 6'hc == buf_6_rs2_paddr ? io_avail_list_12 : _GEN_843; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_845 = 6'hd == buf_6_rs2_paddr ? io_avail_list_13 : _GEN_844; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_846 = 6'he == buf_6_rs2_paddr ? io_avail_list_14 : _GEN_845; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_847 = 6'hf == buf_6_rs2_paddr ? io_avail_list_15 : _GEN_846; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_848 = 6'h10 == buf_6_rs2_paddr ? io_avail_list_16 : _GEN_847; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_849 = 6'h11 == buf_6_rs2_paddr ? io_avail_list_17 : _GEN_848; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_850 = 6'h12 == buf_6_rs2_paddr ? io_avail_list_18 : _GEN_849; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_851 = 6'h13 == buf_6_rs2_paddr ? io_avail_list_19 : _GEN_850; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_852 = 6'h14 == buf_6_rs2_paddr ? io_avail_list_20 : _GEN_851; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_853 = 6'h15 == buf_6_rs2_paddr ? io_avail_list_21 : _GEN_852; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_854 = 6'h16 == buf_6_rs2_paddr ? io_avail_list_22 : _GEN_853; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_855 = 6'h17 == buf_6_rs2_paddr ? io_avail_list_23 : _GEN_854; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_856 = 6'h18 == buf_6_rs2_paddr ? io_avail_list_24 : _GEN_855; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_857 = 6'h19 == buf_6_rs2_paddr ? io_avail_list_25 : _GEN_856; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_858 = 6'h1a == buf_6_rs2_paddr ? io_avail_list_26 : _GEN_857; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_859 = 6'h1b == buf_6_rs2_paddr ? io_avail_list_27 : _GEN_858; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_860 = 6'h1c == buf_6_rs2_paddr ? io_avail_list_28 : _GEN_859; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_861 = 6'h1d == buf_6_rs2_paddr ? io_avail_list_29 : _GEN_860; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_862 = 6'h1e == buf_6_rs2_paddr ? io_avail_list_30 : _GEN_861; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_863 = 6'h1f == buf_6_rs2_paddr ? io_avail_list_31 : _GEN_862; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_864 = 6'h20 == buf_6_rs2_paddr ? io_avail_list_32 : _GEN_863; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_865 = 6'h21 == buf_6_rs2_paddr ? io_avail_list_33 : _GEN_864; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_866 = 6'h22 == buf_6_rs2_paddr ? io_avail_list_34 : _GEN_865; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_867 = 6'h23 == buf_6_rs2_paddr ? io_avail_list_35 : _GEN_866; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_868 = 6'h24 == buf_6_rs2_paddr ? io_avail_list_36 : _GEN_867; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_869 = 6'h25 == buf_6_rs2_paddr ? io_avail_list_37 : _GEN_868; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_870 = 6'h26 == buf_6_rs2_paddr ? io_avail_list_38 : _GEN_869; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_871 = 6'h27 == buf_6_rs2_paddr ? io_avail_list_39 : _GEN_870; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_872 = 6'h28 == buf_6_rs2_paddr ? io_avail_list_40 : _GEN_871; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_873 = 6'h29 == buf_6_rs2_paddr ? io_avail_list_41 : _GEN_872; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_874 = 6'h2a == buf_6_rs2_paddr ? io_avail_list_42 : _GEN_873; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_875 = 6'h2b == buf_6_rs2_paddr ? io_avail_list_43 : _GEN_874; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_876 = 6'h2c == buf_6_rs2_paddr ? io_avail_list_44 : _GEN_875; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_877 = 6'h2d == buf_6_rs2_paddr ? io_avail_list_45 : _GEN_876; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_878 = 6'h2e == buf_6_rs2_paddr ? io_avail_list_46 : _GEN_877; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_879 = 6'h2f == buf_6_rs2_paddr ? io_avail_list_47 : _GEN_878; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_880 = 6'h30 == buf_6_rs2_paddr ? io_avail_list_48 : _GEN_879; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_881 = 6'h31 == buf_6_rs2_paddr ? io_avail_list_49 : _GEN_880; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_882 = 6'h32 == buf_6_rs2_paddr ? io_avail_list_50 : _GEN_881; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_883 = 6'h33 == buf_6_rs2_paddr ? io_avail_list_51 : _GEN_882; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_884 = 6'h34 == buf_6_rs2_paddr ? io_avail_list_52 : _GEN_883; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_885 = 6'h35 == buf_6_rs2_paddr ? io_avail_list_53 : _GEN_884; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_886 = 6'h36 == buf_6_rs2_paddr ? io_avail_list_54 : _GEN_885; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_887 = 6'h37 == buf_6_rs2_paddr ? io_avail_list_55 : _GEN_886; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_888 = 6'h38 == buf_6_rs2_paddr ? io_avail_list_56 : _GEN_887; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_889 = 6'h39 == buf_6_rs2_paddr ? io_avail_list_57 : _GEN_888; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_890 = 6'h3a == buf_6_rs2_paddr ? io_avail_list_58 : _GEN_889; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_891 = 6'h3b == buf_6_rs2_paddr ? io_avail_list_59 : _GEN_890; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_892 = 6'h3c == buf_6_rs2_paddr ? io_avail_list_60 : _GEN_891; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_893 = 6'h3d == buf_6_rs2_paddr ? io_avail_list_61 : _GEN_892; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_894 = 6'h3e == buf_6_rs2_paddr ? io_avail_list_62 : _GEN_893; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_895 = 6'h3f == buf_6_rs2_paddr ? io_avail_list_63 : _GEN_894; // @[IssueUnit.scala 133:{34,34}]
  wire  ready_list_6 = _GEN_831 & _GEN_895 & ~is_sys_6; // @[IssueUnit.scala 133:59]
  wire  _GEN_897 = 6'h1 == buf_7_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_898 = 6'h2 == buf_7_rs1_paddr ? io_avail_list_2 : _GEN_897; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_899 = 6'h3 == buf_7_rs1_paddr ? io_avail_list_3 : _GEN_898; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_900 = 6'h4 == buf_7_rs1_paddr ? io_avail_list_4 : _GEN_899; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_901 = 6'h5 == buf_7_rs1_paddr ? io_avail_list_5 : _GEN_900; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_902 = 6'h6 == buf_7_rs1_paddr ? io_avail_list_6 : _GEN_901; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_903 = 6'h7 == buf_7_rs1_paddr ? io_avail_list_7 : _GEN_902; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_904 = 6'h8 == buf_7_rs1_paddr ? io_avail_list_8 : _GEN_903; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_905 = 6'h9 == buf_7_rs1_paddr ? io_avail_list_9 : _GEN_904; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_906 = 6'ha == buf_7_rs1_paddr ? io_avail_list_10 : _GEN_905; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_907 = 6'hb == buf_7_rs1_paddr ? io_avail_list_11 : _GEN_906; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_908 = 6'hc == buf_7_rs1_paddr ? io_avail_list_12 : _GEN_907; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_909 = 6'hd == buf_7_rs1_paddr ? io_avail_list_13 : _GEN_908; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_910 = 6'he == buf_7_rs1_paddr ? io_avail_list_14 : _GEN_909; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_911 = 6'hf == buf_7_rs1_paddr ? io_avail_list_15 : _GEN_910; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_912 = 6'h10 == buf_7_rs1_paddr ? io_avail_list_16 : _GEN_911; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_913 = 6'h11 == buf_7_rs1_paddr ? io_avail_list_17 : _GEN_912; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_914 = 6'h12 == buf_7_rs1_paddr ? io_avail_list_18 : _GEN_913; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_915 = 6'h13 == buf_7_rs1_paddr ? io_avail_list_19 : _GEN_914; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_916 = 6'h14 == buf_7_rs1_paddr ? io_avail_list_20 : _GEN_915; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_917 = 6'h15 == buf_7_rs1_paddr ? io_avail_list_21 : _GEN_916; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_918 = 6'h16 == buf_7_rs1_paddr ? io_avail_list_22 : _GEN_917; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_919 = 6'h17 == buf_7_rs1_paddr ? io_avail_list_23 : _GEN_918; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_920 = 6'h18 == buf_7_rs1_paddr ? io_avail_list_24 : _GEN_919; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_921 = 6'h19 == buf_7_rs1_paddr ? io_avail_list_25 : _GEN_920; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_922 = 6'h1a == buf_7_rs1_paddr ? io_avail_list_26 : _GEN_921; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_923 = 6'h1b == buf_7_rs1_paddr ? io_avail_list_27 : _GEN_922; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_924 = 6'h1c == buf_7_rs1_paddr ? io_avail_list_28 : _GEN_923; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_925 = 6'h1d == buf_7_rs1_paddr ? io_avail_list_29 : _GEN_924; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_926 = 6'h1e == buf_7_rs1_paddr ? io_avail_list_30 : _GEN_925; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_927 = 6'h1f == buf_7_rs1_paddr ? io_avail_list_31 : _GEN_926; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_928 = 6'h20 == buf_7_rs1_paddr ? io_avail_list_32 : _GEN_927; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_929 = 6'h21 == buf_7_rs1_paddr ? io_avail_list_33 : _GEN_928; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_930 = 6'h22 == buf_7_rs1_paddr ? io_avail_list_34 : _GEN_929; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_931 = 6'h23 == buf_7_rs1_paddr ? io_avail_list_35 : _GEN_930; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_932 = 6'h24 == buf_7_rs1_paddr ? io_avail_list_36 : _GEN_931; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_933 = 6'h25 == buf_7_rs1_paddr ? io_avail_list_37 : _GEN_932; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_934 = 6'h26 == buf_7_rs1_paddr ? io_avail_list_38 : _GEN_933; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_935 = 6'h27 == buf_7_rs1_paddr ? io_avail_list_39 : _GEN_934; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_936 = 6'h28 == buf_7_rs1_paddr ? io_avail_list_40 : _GEN_935; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_937 = 6'h29 == buf_7_rs1_paddr ? io_avail_list_41 : _GEN_936; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_938 = 6'h2a == buf_7_rs1_paddr ? io_avail_list_42 : _GEN_937; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_939 = 6'h2b == buf_7_rs1_paddr ? io_avail_list_43 : _GEN_938; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_940 = 6'h2c == buf_7_rs1_paddr ? io_avail_list_44 : _GEN_939; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_941 = 6'h2d == buf_7_rs1_paddr ? io_avail_list_45 : _GEN_940; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_942 = 6'h2e == buf_7_rs1_paddr ? io_avail_list_46 : _GEN_941; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_943 = 6'h2f == buf_7_rs1_paddr ? io_avail_list_47 : _GEN_942; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_944 = 6'h30 == buf_7_rs1_paddr ? io_avail_list_48 : _GEN_943; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_945 = 6'h31 == buf_7_rs1_paddr ? io_avail_list_49 : _GEN_944; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_946 = 6'h32 == buf_7_rs1_paddr ? io_avail_list_50 : _GEN_945; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_947 = 6'h33 == buf_7_rs1_paddr ? io_avail_list_51 : _GEN_946; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_948 = 6'h34 == buf_7_rs1_paddr ? io_avail_list_52 : _GEN_947; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_949 = 6'h35 == buf_7_rs1_paddr ? io_avail_list_53 : _GEN_948; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_950 = 6'h36 == buf_7_rs1_paddr ? io_avail_list_54 : _GEN_949; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_951 = 6'h37 == buf_7_rs1_paddr ? io_avail_list_55 : _GEN_950; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_952 = 6'h38 == buf_7_rs1_paddr ? io_avail_list_56 : _GEN_951; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_953 = 6'h39 == buf_7_rs1_paddr ? io_avail_list_57 : _GEN_952; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_954 = 6'h3a == buf_7_rs1_paddr ? io_avail_list_58 : _GEN_953; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_955 = 6'h3b == buf_7_rs1_paddr ? io_avail_list_59 : _GEN_954; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_956 = 6'h3c == buf_7_rs1_paddr ? io_avail_list_60 : _GEN_955; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_957 = 6'h3d == buf_7_rs1_paddr ? io_avail_list_61 : _GEN_956; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_958 = 6'h3e == buf_7_rs1_paddr ? io_avail_list_62 : _GEN_957; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_959 = 6'h3f == buf_7_rs1_paddr ? io_avail_list_63 : _GEN_958; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_961 = 6'h1 == buf_7_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_962 = 6'h2 == buf_7_rs2_paddr ? io_avail_list_2 : _GEN_961; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_963 = 6'h3 == buf_7_rs2_paddr ? io_avail_list_3 : _GEN_962; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_964 = 6'h4 == buf_7_rs2_paddr ? io_avail_list_4 : _GEN_963; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_965 = 6'h5 == buf_7_rs2_paddr ? io_avail_list_5 : _GEN_964; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_966 = 6'h6 == buf_7_rs2_paddr ? io_avail_list_6 : _GEN_965; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_967 = 6'h7 == buf_7_rs2_paddr ? io_avail_list_7 : _GEN_966; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_968 = 6'h8 == buf_7_rs2_paddr ? io_avail_list_8 : _GEN_967; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_969 = 6'h9 == buf_7_rs2_paddr ? io_avail_list_9 : _GEN_968; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_970 = 6'ha == buf_7_rs2_paddr ? io_avail_list_10 : _GEN_969; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_971 = 6'hb == buf_7_rs2_paddr ? io_avail_list_11 : _GEN_970; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_972 = 6'hc == buf_7_rs2_paddr ? io_avail_list_12 : _GEN_971; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_973 = 6'hd == buf_7_rs2_paddr ? io_avail_list_13 : _GEN_972; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_974 = 6'he == buf_7_rs2_paddr ? io_avail_list_14 : _GEN_973; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_975 = 6'hf == buf_7_rs2_paddr ? io_avail_list_15 : _GEN_974; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_976 = 6'h10 == buf_7_rs2_paddr ? io_avail_list_16 : _GEN_975; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_977 = 6'h11 == buf_7_rs2_paddr ? io_avail_list_17 : _GEN_976; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_978 = 6'h12 == buf_7_rs2_paddr ? io_avail_list_18 : _GEN_977; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_979 = 6'h13 == buf_7_rs2_paddr ? io_avail_list_19 : _GEN_978; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_980 = 6'h14 == buf_7_rs2_paddr ? io_avail_list_20 : _GEN_979; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_981 = 6'h15 == buf_7_rs2_paddr ? io_avail_list_21 : _GEN_980; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_982 = 6'h16 == buf_7_rs2_paddr ? io_avail_list_22 : _GEN_981; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_983 = 6'h17 == buf_7_rs2_paddr ? io_avail_list_23 : _GEN_982; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_984 = 6'h18 == buf_7_rs2_paddr ? io_avail_list_24 : _GEN_983; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_985 = 6'h19 == buf_7_rs2_paddr ? io_avail_list_25 : _GEN_984; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_986 = 6'h1a == buf_7_rs2_paddr ? io_avail_list_26 : _GEN_985; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_987 = 6'h1b == buf_7_rs2_paddr ? io_avail_list_27 : _GEN_986; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_988 = 6'h1c == buf_7_rs2_paddr ? io_avail_list_28 : _GEN_987; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_989 = 6'h1d == buf_7_rs2_paddr ? io_avail_list_29 : _GEN_988; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_990 = 6'h1e == buf_7_rs2_paddr ? io_avail_list_30 : _GEN_989; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_991 = 6'h1f == buf_7_rs2_paddr ? io_avail_list_31 : _GEN_990; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_992 = 6'h20 == buf_7_rs2_paddr ? io_avail_list_32 : _GEN_991; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_993 = 6'h21 == buf_7_rs2_paddr ? io_avail_list_33 : _GEN_992; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_994 = 6'h22 == buf_7_rs2_paddr ? io_avail_list_34 : _GEN_993; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_995 = 6'h23 == buf_7_rs2_paddr ? io_avail_list_35 : _GEN_994; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_996 = 6'h24 == buf_7_rs2_paddr ? io_avail_list_36 : _GEN_995; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_997 = 6'h25 == buf_7_rs2_paddr ? io_avail_list_37 : _GEN_996; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_998 = 6'h26 == buf_7_rs2_paddr ? io_avail_list_38 : _GEN_997; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_999 = 6'h27 == buf_7_rs2_paddr ? io_avail_list_39 : _GEN_998; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1000 = 6'h28 == buf_7_rs2_paddr ? io_avail_list_40 : _GEN_999; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1001 = 6'h29 == buf_7_rs2_paddr ? io_avail_list_41 : _GEN_1000; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1002 = 6'h2a == buf_7_rs2_paddr ? io_avail_list_42 : _GEN_1001; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1003 = 6'h2b == buf_7_rs2_paddr ? io_avail_list_43 : _GEN_1002; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1004 = 6'h2c == buf_7_rs2_paddr ? io_avail_list_44 : _GEN_1003; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1005 = 6'h2d == buf_7_rs2_paddr ? io_avail_list_45 : _GEN_1004; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1006 = 6'h2e == buf_7_rs2_paddr ? io_avail_list_46 : _GEN_1005; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1007 = 6'h2f == buf_7_rs2_paddr ? io_avail_list_47 : _GEN_1006; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1008 = 6'h30 == buf_7_rs2_paddr ? io_avail_list_48 : _GEN_1007; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1009 = 6'h31 == buf_7_rs2_paddr ? io_avail_list_49 : _GEN_1008; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1010 = 6'h32 == buf_7_rs2_paddr ? io_avail_list_50 : _GEN_1009; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1011 = 6'h33 == buf_7_rs2_paddr ? io_avail_list_51 : _GEN_1010; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1012 = 6'h34 == buf_7_rs2_paddr ? io_avail_list_52 : _GEN_1011; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1013 = 6'h35 == buf_7_rs2_paddr ? io_avail_list_53 : _GEN_1012; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1014 = 6'h36 == buf_7_rs2_paddr ? io_avail_list_54 : _GEN_1013; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1015 = 6'h37 == buf_7_rs2_paddr ? io_avail_list_55 : _GEN_1014; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1016 = 6'h38 == buf_7_rs2_paddr ? io_avail_list_56 : _GEN_1015; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1017 = 6'h39 == buf_7_rs2_paddr ? io_avail_list_57 : _GEN_1016; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1018 = 6'h3a == buf_7_rs2_paddr ? io_avail_list_58 : _GEN_1017; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1019 = 6'h3b == buf_7_rs2_paddr ? io_avail_list_59 : _GEN_1018; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1020 = 6'h3c == buf_7_rs2_paddr ? io_avail_list_60 : _GEN_1019; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1021 = 6'h3d == buf_7_rs2_paddr ? io_avail_list_61 : _GEN_1020; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1022 = 6'h3e == buf_7_rs2_paddr ? io_avail_list_62 : _GEN_1021; // @[IssueUnit.scala 133:{34,34}]
  wire  _GEN_1023 = 6'h3f == buf_7_rs2_paddr ? io_avail_list_63 : _GEN_1022; // @[IssueUnit.scala 133:{34,34}]
  wire  ready_list_7 = _GEN_959 & _GEN_1023 & ~is_sys_7; // @[IssueUnit.scala 133:59]
  wire [7:0] rl0 = {ready_list_7,ready_list_6,ready_list_5,ready_list_4,ready_list_3,ready_list_2,ready_list_1,
    ready_list_0}; // @[Cat.scala 30:58]
  wire [2:0] _T_59 = rl0[6] ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_60 = rl0[5] ? 3'h5 : _T_59; // @[Mux.scala 47:69]
  wire [2:0] _T_61 = rl0[4] ? 3'h4 : _T_60; // @[Mux.scala 47:69]
  wire [2:0] _T_62 = rl0[3] ? 3'h3 : _T_61; // @[Mux.scala 47:69]
  wire [2:0] _T_63 = rl0[2] ? 3'h2 : _T_62; // @[Mux.scala 47:69]
  wire [2:0] _T_64 = rl0[1] ? 3'h1 : _T_63; // @[Mux.scala 47:69]
  wire [2:0] deq_vec_0 = rl0[0] ? 3'h0 : _T_64; // @[Mux.scala 47:69]
  wire  _GEN_1025 = 3'h1 == deq_vec_0 ? ready_list_1 : ready_list_0; // @[IssueUnit.scala 140:{20,20}]
  wire  _GEN_1026 = 3'h2 == deq_vec_0 ? ready_list_2 : _GEN_1025; // @[IssueUnit.scala 140:{20,20}]
  wire  _GEN_1027 = 3'h3 == deq_vec_0 ? ready_list_3 : _GEN_1026; // @[IssueUnit.scala 140:{20,20}]
  wire  _GEN_1028 = 3'h4 == deq_vec_0 ? ready_list_4 : _GEN_1027; // @[IssueUnit.scala 140:{20,20}]
  wire  _GEN_1029 = 3'h5 == deq_vec_0 ? ready_list_5 : _GEN_1028; // @[IssueUnit.scala 140:{20,20}]
  wire  _GEN_1030 = 3'h6 == deq_vec_0 ? ready_list_6 : _GEN_1029; // @[IssueUnit.scala 140:{20,20}]
  wire  deq_vec_valid_0 = 3'h7 == deq_vec_0 ? ready_list_7 : _GEN_1030; // @[IssueUnit.scala 140:{20,20}]
  wire [7:0] _T_66 = 8'h1 << deq_vec_0; // @[OneHot.scala 65:12]
  wire [7:0] _T_68 = ~_T_66; // @[IssueUnit.scala 142:19]
  wire [7:0] rl1 = rl0 & _T_68; // @[IssueUnit.scala 142:17]
  wire [2:0] _T_77 = rl1[6] ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_78 = rl1[5] ? 3'h5 : _T_77; // @[Mux.scala 47:69]
  wire [2:0] _T_79 = rl1[4] ? 3'h4 : _T_78; // @[Mux.scala 47:69]
  wire [2:0] _T_80 = rl1[3] ? 3'h3 : _T_79; // @[Mux.scala 47:69]
  wire [2:0] _T_81 = rl1[2] ? 3'h2 : _T_80; // @[Mux.scala 47:69]
  wire [2:0] _T_82 = rl1[1] ? 3'h1 : _T_81; // @[Mux.scala 47:69]
  wire [2:0] deq_vec_1 = rl1[0] ? 3'h0 : _T_82; // @[Mux.scala 47:69]
  wire  _GEN_1033 = 3'h1 == deq_vec_1 ? ready_list_1 : ready_list_0; // @[IssueUnit.scala 144:{46,46}]
  wire  _GEN_1034 = 3'h2 == deq_vec_1 ? ready_list_2 : _GEN_1033; // @[IssueUnit.scala 144:{46,46}]
  wire  _GEN_1035 = 3'h3 == deq_vec_1 ? ready_list_3 : _GEN_1034; // @[IssueUnit.scala 144:{46,46}]
  wire  _GEN_1036 = 3'h4 == deq_vec_1 ? ready_list_4 : _GEN_1035; // @[IssueUnit.scala 144:{46,46}]
  wire  _GEN_1037 = 3'h5 == deq_vec_1 ? ready_list_5 : _GEN_1036; // @[IssueUnit.scala 144:{46,46}]
  wire  _GEN_1038 = 3'h6 == deq_vec_1 ? ready_list_6 : _GEN_1037; // @[IssueUnit.scala 144:{46,46}]
  wire  _GEN_1039 = 3'h7 == deq_vec_1 ? ready_list_7 : _GEN_1038; // @[IssueUnit.scala 144:{46,46}]
  wire  deq_vec_valid_1 = _GEN_1039 & deq_vec_1 != deq_vec_0; // @[IssueUnit.scala 144:46]
  wire [3:0] _GEN_1041 = 3'h1 == deq_vec_0 ? buf_1_rob_addr : buf_0_rob_addr; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1042 = 3'h2 == deq_vec_0 ? buf_2_rob_addr : _GEN_1041; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1043 = 3'h3 == deq_vec_0 ? buf_3_rob_addr : _GEN_1042; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1044 = 3'h4 == deq_vec_0 ? buf_4_rob_addr : _GEN_1043; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1045 = 3'h5 == deq_vec_0 ? buf_5_rob_addr : _GEN_1044; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1046 = 3'h6 == deq_vec_0 ? buf_6_rob_addr : _GEN_1045; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1057 = 3'h1 == deq_vec_0 ? buf_1_rd_paddr : buf_0_rd_paddr; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1058 = 3'h2 == deq_vec_0 ? buf_2_rd_paddr : _GEN_1057; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1059 = 3'h3 == deq_vec_0 ? buf_3_rd_paddr : _GEN_1058; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1060 = 3'h4 == deq_vec_0 ? buf_4_rd_paddr : _GEN_1059; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1061 = 3'h5 == deq_vec_0 ? buf_5_rd_paddr : _GEN_1060; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1062 = 3'h6 == deq_vec_0 ? buf_6_rd_paddr : _GEN_1061; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1065 = 3'h1 == deq_vec_0 ? buf_1_rs2_paddr : buf_0_rs2_paddr; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1066 = 3'h2 == deq_vec_0 ? buf_2_rs2_paddr : _GEN_1065; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1067 = 3'h3 == deq_vec_0 ? buf_3_rs2_paddr : _GEN_1066; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1068 = 3'h4 == deq_vec_0 ? buf_4_rs2_paddr : _GEN_1067; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1069 = 3'h5 == deq_vec_0 ? buf_5_rs2_paddr : _GEN_1068; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1070 = 3'h6 == deq_vec_0 ? buf_6_rs2_paddr : _GEN_1069; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1073 = 3'h1 == deq_vec_0 ? buf_1_rs1_paddr : buf_0_rs1_paddr; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1074 = 3'h2 == deq_vec_0 ? buf_2_rs1_paddr : _GEN_1073; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1075 = 3'h3 == deq_vec_0 ? buf_3_rs1_paddr : _GEN_1074; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1076 = 3'h4 == deq_vec_0 ? buf_4_rs1_paddr : _GEN_1075; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1077 = 3'h5 == deq_vec_0 ? buf_5_rs1_paddr : _GEN_1076; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1078 = 3'h6 == deq_vec_0 ? buf_6_rs1_paddr : _GEN_1077; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1081 = 3'h1 == deq_vec_0 ? buf_1_pred_bpc : buf_0_pred_bpc; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1082 = 3'h2 == deq_vec_0 ? buf_2_pred_bpc : _GEN_1081; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1083 = 3'h3 == deq_vec_0 ? buf_3_pred_bpc : _GEN_1082; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1084 = 3'h4 == deq_vec_0 ? buf_4_pred_bpc : _GEN_1083; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1085 = 3'h5 == deq_vec_0 ? buf_5_pred_bpc : _GEN_1084; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1086 = 3'h6 == deq_vec_0 ? buf_6_pred_bpc : _GEN_1085; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1089 = 3'h1 == deq_vec_0 ? buf_1_pred_br : buf_0_pred_br; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1090 = 3'h2 == deq_vec_0 ? buf_2_pred_br : _GEN_1089; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1091 = 3'h3 == deq_vec_0 ? buf_3_pred_br : _GEN_1090; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1092 = 3'h4 == deq_vec_0 ? buf_4_pred_br : _GEN_1091; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1093 = 3'h5 == deq_vec_0 ? buf_5_pred_br : _GEN_1092; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1094 = 3'h6 == deq_vec_0 ? buf_6_pred_br : _GEN_1093; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1097 = 3'h1 == deq_vec_0 ? buf_1_imm : buf_0_imm; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1098 = 3'h2 == deq_vec_0 ? buf_2_imm : _GEN_1097; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1099 = 3'h3 == deq_vec_0 ? buf_3_imm : _GEN_1098; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1100 = 3'h4 == deq_vec_0 ? buf_4_imm : _GEN_1099; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1101 = 3'h5 == deq_vec_0 ? buf_5_imm : _GEN_1100; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1102 = 3'h6 == deq_vec_0 ? buf_6_imm : _GEN_1101; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1105 = 3'h1 == deq_vec_0 ? buf_1_rd_en : buf_0_rd_en; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1106 = 3'h2 == deq_vec_0 ? buf_2_rd_en : _GEN_1105; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1107 = 3'h3 == deq_vec_0 ? buf_3_rd_en : _GEN_1106; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1108 = 3'h4 == deq_vec_0 ? buf_4_rd_en : _GEN_1107; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1109 = 3'h5 == deq_vec_0 ? buf_5_rd_en : _GEN_1108; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1110 = 3'h6 == deq_vec_0 ? buf_6_rd_en : _GEN_1109; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1137 = 3'h1 == deq_vec_0 ? buf_1_rs2_src : buf_0_rs2_src; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1138 = 3'h2 == deq_vec_0 ? buf_2_rs2_src : _GEN_1137; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1139 = 3'h3 == deq_vec_0 ? buf_3_rs2_src : _GEN_1138; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1140 = 3'h4 == deq_vec_0 ? buf_4_rs2_src : _GEN_1139; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1141 = 3'h5 == deq_vec_0 ? buf_5_rs2_src : _GEN_1140; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1142 = 3'h6 == deq_vec_0 ? buf_6_rs2_src : _GEN_1141; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1145 = 3'h1 == deq_vec_0 ? buf_1_rs1_src : buf_0_rs1_src; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1146 = 3'h2 == deq_vec_0 ? buf_2_rs1_src : _GEN_1145; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1147 = 3'h3 == deq_vec_0 ? buf_3_rs1_src : _GEN_1146; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1148 = 3'h4 == deq_vec_0 ? buf_4_rs1_src : _GEN_1147; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1149 = 3'h5 == deq_vec_0 ? buf_5_rs1_src : _GEN_1148; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1150 = 3'h6 == deq_vec_0 ? buf_6_rs1_src : _GEN_1149; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1153 = 3'h1 == deq_vec_0 ? buf_1_w_type : buf_0_w_type; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1154 = 3'h2 == deq_vec_0 ? buf_2_w_type : _GEN_1153; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1155 = 3'h3 == deq_vec_0 ? buf_3_w_type : _GEN_1154; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1156 = 3'h4 == deq_vec_0 ? buf_4_w_type : _GEN_1155; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1157 = 3'h5 == deq_vec_0 ? buf_5_w_type : _GEN_1156; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1158 = 3'h6 == deq_vec_0 ? buf_6_w_type : _GEN_1157; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1161 = 3'h1 == deq_vec_0 ? buf_1_sys_code : buf_0_sys_code; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1162 = 3'h2 == deq_vec_0 ? buf_2_sys_code : _GEN_1161; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1163 = 3'h3 == deq_vec_0 ? buf_3_sys_code : _GEN_1162; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1164 = 3'h4 == deq_vec_0 ? buf_4_sys_code : _GEN_1163; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1165 = 3'h5 == deq_vec_0 ? buf_5_sys_code : _GEN_1164; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1166 = 3'h6 == deq_vec_0 ? buf_6_sys_code : _GEN_1165; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1185 = 3'h1 == deq_vec_0 ? buf_1_jmp_code : buf_0_jmp_code; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1186 = 3'h2 == deq_vec_0 ? buf_2_jmp_code : _GEN_1185; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1187 = 3'h3 == deq_vec_0 ? buf_3_jmp_code : _GEN_1186; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1188 = 3'h4 == deq_vec_0 ? buf_4_jmp_code : _GEN_1187; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1189 = 3'h5 == deq_vec_0 ? buf_5_jmp_code : _GEN_1188; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1190 = 3'h6 == deq_vec_0 ? buf_6_jmp_code : _GEN_1189; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1193 = 3'h1 == deq_vec_0 ? buf_1_alu_code : buf_0_alu_code; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1194 = 3'h2 == deq_vec_0 ? buf_2_alu_code : _GEN_1193; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1195 = 3'h3 == deq_vec_0 ? buf_3_alu_code : _GEN_1194; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1196 = 3'h4 == deq_vec_0 ? buf_4_alu_code : _GEN_1195; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1197 = 3'h5 == deq_vec_0 ? buf_5_alu_code : _GEN_1196; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1198 = 3'h6 == deq_vec_0 ? buf_6_alu_code : _GEN_1197; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1201 = 3'h1 == deq_vec_0 ? buf_1_fu_code : buf_0_fu_code; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1202 = 3'h2 == deq_vec_0 ? buf_2_fu_code : _GEN_1201; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1203 = 3'h3 == deq_vec_0 ? buf_3_fu_code : _GEN_1202; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1204 = 3'h4 == deq_vec_0 ? buf_4_fu_code : _GEN_1203; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1205 = 3'h5 == deq_vec_0 ? buf_5_fu_code : _GEN_1204; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1206 = 3'h6 == deq_vec_0 ? buf_6_fu_code : _GEN_1205; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1209 = 3'h1 == deq_vec_0 ? buf_1_inst : buf_0_inst; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1210 = 3'h2 == deq_vec_0 ? buf_2_inst : _GEN_1209; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1211 = 3'h3 == deq_vec_0 ? buf_3_inst : _GEN_1210; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1212 = 3'h4 == deq_vec_0 ? buf_4_inst : _GEN_1211; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1213 = 3'h5 == deq_vec_0 ? buf_5_inst : _GEN_1212; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1214 = 3'h6 == deq_vec_0 ? buf_6_inst : _GEN_1213; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1217 = 3'h1 == deq_vec_0 ? buf_1_npc : buf_0_npc; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1218 = 3'h2 == deq_vec_0 ? buf_2_npc : _GEN_1217; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1219 = 3'h3 == deq_vec_0 ? buf_3_npc : _GEN_1218; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1220 = 3'h4 == deq_vec_0 ? buf_4_npc : _GEN_1219; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1221 = 3'h5 == deq_vec_0 ? buf_5_npc : _GEN_1220; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1222 = 3'h6 == deq_vec_0 ? buf_6_npc : _GEN_1221; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1225 = 3'h1 == deq_vec_0 ? buf_1_pc : buf_0_pc; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1226 = 3'h2 == deq_vec_0 ? buf_2_pc : _GEN_1225; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1227 = 3'h3 == deq_vec_0 ? buf_3_pc : _GEN_1226; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1228 = 3'h4 == deq_vec_0 ? buf_4_pc : _GEN_1227; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1229 = 3'h5 == deq_vec_0 ? buf_5_pc : _GEN_1228; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1230 = 3'h6 == deq_vec_0 ? buf_6_pc : _GEN_1229; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1233 = 3'h1 == deq_vec_0 ? buf_1_valid : buf_0_valid; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1234 = 3'h2 == deq_vec_0 ? buf_2_valid : _GEN_1233; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1235 = 3'h3 == deq_vec_0 ? buf_3_valid : _GEN_1234; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1236 = 3'h4 == deq_vec_0 ? buf_4_valid : _GEN_1235; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1237 = 3'h5 == deq_vec_0 ? buf_5_valid : _GEN_1236; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1238 = 3'h6 == deq_vec_0 ? buf_6_valid : _GEN_1237; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1239 = 3'h7 == deq_vec_0 ? buf_7_valid : _GEN_1238; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1241 = 3'h1 == deq_vec_1 ? buf_1_rob_addr : buf_0_rob_addr; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1242 = 3'h2 == deq_vec_1 ? buf_2_rob_addr : _GEN_1241; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1243 = 3'h3 == deq_vec_1 ? buf_3_rob_addr : _GEN_1242; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1244 = 3'h4 == deq_vec_1 ? buf_4_rob_addr : _GEN_1243; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1245 = 3'h5 == deq_vec_1 ? buf_5_rob_addr : _GEN_1244; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1246 = 3'h6 == deq_vec_1 ? buf_6_rob_addr : _GEN_1245; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1257 = 3'h1 == deq_vec_1 ? buf_1_rd_paddr : buf_0_rd_paddr; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1258 = 3'h2 == deq_vec_1 ? buf_2_rd_paddr : _GEN_1257; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1259 = 3'h3 == deq_vec_1 ? buf_3_rd_paddr : _GEN_1258; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1260 = 3'h4 == deq_vec_1 ? buf_4_rd_paddr : _GEN_1259; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1261 = 3'h5 == deq_vec_1 ? buf_5_rd_paddr : _GEN_1260; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1262 = 3'h6 == deq_vec_1 ? buf_6_rd_paddr : _GEN_1261; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1265 = 3'h1 == deq_vec_1 ? buf_1_rs2_paddr : buf_0_rs2_paddr; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1266 = 3'h2 == deq_vec_1 ? buf_2_rs2_paddr : _GEN_1265; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1267 = 3'h3 == deq_vec_1 ? buf_3_rs2_paddr : _GEN_1266; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1268 = 3'h4 == deq_vec_1 ? buf_4_rs2_paddr : _GEN_1267; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1269 = 3'h5 == deq_vec_1 ? buf_5_rs2_paddr : _GEN_1268; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1270 = 3'h6 == deq_vec_1 ? buf_6_rs2_paddr : _GEN_1269; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1273 = 3'h1 == deq_vec_1 ? buf_1_rs1_paddr : buf_0_rs1_paddr; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1274 = 3'h2 == deq_vec_1 ? buf_2_rs1_paddr : _GEN_1273; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1275 = 3'h3 == deq_vec_1 ? buf_3_rs1_paddr : _GEN_1274; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1276 = 3'h4 == deq_vec_1 ? buf_4_rs1_paddr : _GEN_1275; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1277 = 3'h5 == deq_vec_1 ? buf_5_rs1_paddr : _GEN_1276; // @[IssueUnit.scala 148:{15,15}]
  wire [5:0] _GEN_1278 = 3'h6 == deq_vec_1 ? buf_6_rs1_paddr : _GEN_1277; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1281 = 3'h1 == deq_vec_1 ? buf_1_pred_bpc : buf_0_pred_bpc; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1282 = 3'h2 == deq_vec_1 ? buf_2_pred_bpc : _GEN_1281; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1283 = 3'h3 == deq_vec_1 ? buf_3_pred_bpc : _GEN_1282; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1284 = 3'h4 == deq_vec_1 ? buf_4_pred_bpc : _GEN_1283; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1285 = 3'h5 == deq_vec_1 ? buf_5_pred_bpc : _GEN_1284; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1286 = 3'h6 == deq_vec_1 ? buf_6_pred_bpc : _GEN_1285; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1289 = 3'h1 == deq_vec_1 ? buf_1_pred_br : buf_0_pred_br; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1290 = 3'h2 == deq_vec_1 ? buf_2_pred_br : _GEN_1289; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1291 = 3'h3 == deq_vec_1 ? buf_3_pred_br : _GEN_1290; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1292 = 3'h4 == deq_vec_1 ? buf_4_pred_br : _GEN_1291; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1293 = 3'h5 == deq_vec_1 ? buf_5_pred_br : _GEN_1292; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1294 = 3'h6 == deq_vec_1 ? buf_6_pred_br : _GEN_1293; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1297 = 3'h1 == deq_vec_1 ? buf_1_imm : buf_0_imm; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1298 = 3'h2 == deq_vec_1 ? buf_2_imm : _GEN_1297; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1299 = 3'h3 == deq_vec_1 ? buf_3_imm : _GEN_1298; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1300 = 3'h4 == deq_vec_1 ? buf_4_imm : _GEN_1299; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1301 = 3'h5 == deq_vec_1 ? buf_5_imm : _GEN_1300; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1302 = 3'h6 == deq_vec_1 ? buf_6_imm : _GEN_1301; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1305 = 3'h1 == deq_vec_1 ? buf_1_rd_en : buf_0_rd_en; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1306 = 3'h2 == deq_vec_1 ? buf_2_rd_en : _GEN_1305; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1307 = 3'h3 == deq_vec_1 ? buf_3_rd_en : _GEN_1306; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1308 = 3'h4 == deq_vec_1 ? buf_4_rd_en : _GEN_1307; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1309 = 3'h5 == deq_vec_1 ? buf_5_rd_en : _GEN_1308; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1310 = 3'h6 == deq_vec_1 ? buf_6_rd_en : _GEN_1309; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1337 = 3'h1 == deq_vec_1 ? buf_1_rs2_src : buf_0_rs2_src; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1338 = 3'h2 == deq_vec_1 ? buf_2_rs2_src : _GEN_1337; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1339 = 3'h3 == deq_vec_1 ? buf_3_rs2_src : _GEN_1338; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1340 = 3'h4 == deq_vec_1 ? buf_4_rs2_src : _GEN_1339; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1341 = 3'h5 == deq_vec_1 ? buf_5_rs2_src : _GEN_1340; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1342 = 3'h6 == deq_vec_1 ? buf_6_rs2_src : _GEN_1341; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1345 = 3'h1 == deq_vec_1 ? buf_1_rs1_src : buf_0_rs1_src; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1346 = 3'h2 == deq_vec_1 ? buf_2_rs1_src : _GEN_1345; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1347 = 3'h3 == deq_vec_1 ? buf_3_rs1_src : _GEN_1346; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1348 = 3'h4 == deq_vec_1 ? buf_4_rs1_src : _GEN_1347; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1349 = 3'h5 == deq_vec_1 ? buf_5_rs1_src : _GEN_1348; // @[IssueUnit.scala 148:{15,15}]
  wire [1:0] _GEN_1350 = 3'h6 == deq_vec_1 ? buf_6_rs1_src : _GEN_1349; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1353 = 3'h1 == deq_vec_1 ? buf_1_w_type : buf_0_w_type; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1354 = 3'h2 == deq_vec_1 ? buf_2_w_type : _GEN_1353; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1355 = 3'h3 == deq_vec_1 ? buf_3_w_type : _GEN_1354; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1356 = 3'h4 == deq_vec_1 ? buf_4_w_type : _GEN_1355; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1357 = 3'h5 == deq_vec_1 ? buf_5_w_type : _GEN_1356; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1358 = 3'h6 == deq_vec_1 ? buf_6_w_type : _GEN_1357; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1385 = 3'h1 == deq_vec_1 ? buf_1_jmp_code : buf_0_jmp_code; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1386 = 3'h2 == deq_vec_1 ? buf_2_jmp_code : _GEN_1385; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1387 = 3'h3 == deq_vec_1 ? buf_3_jmp_code : _GEN_1386; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1388 = 3'h4 == deq_vec_1 ? buf_4_jmp_code : _GEN_1387; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1389 = 3'h5 == deq_vec_1 ? buf_5_jmp_code : _GEN_1388; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1390 = 3'h6 == deq_vec_1 ? buf_6_jmp_code : _GEN_1389; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1393 = 3'h1 == deq_vec_1 ? buf_1_alu_code : buf_0_alu_code; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1394 = 3'h2 == deq_vec_1 ? buf_2_alu_code : _GEN_1393; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1395 = 3'h3 == deq_vec_1 ? buf_3_alu_code : _GEN_1394; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1396 = 3'h4 == deq_vec_1 ? buf_4_alu_code : _GEN_1395; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1397 = 3'h5 == deq_vec_1 ? buf_5_alu_code : _GEN_1396; // @[IssueUnit.scala 148:{15,15}]
  wire [3:0] _GEN_1398 = 3'h6 == deq_vec_1 ? buf_6_alu_code : _GEN_1397; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1401 = 3'h1 == deq_vec_1 ? buf_1_fu_code : buf_0_fu_code; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1402 = 3'h2 == deq_vec_1 ? buf_2_fu_code : _GEN_1401; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1403 = 3'h3 == deq_vec_1 ? buf_3_fu_code : _GEN_1402; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1404 = 3'h4 == deq_vec_1 ? buf_4_fu_code : _GEN_1403; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1405 = 3'h5 == deq_vec_1 ? buf_5_fu_code : _GEN_1404; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _GEN_1406 = 3'h6 == deq_vec_1 ? buf_6_fu_code : _GEN_1405; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1417 = 3'h1 == deq_vec_1 ? buf_1_npc : buf_0_npc; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1418 = 3'h2 == deq_vec_1 ? buf_2_npc : _GEN_1417; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1419 = 3'h3 == deq_vec_1 ? buf_3_npc : _GEN_1418; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1420 = 3'h4 == deq_vec_1 ? buf_4_npc : _GEN_1419; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1421 = 3'h5 == deq_vec_1 ? buf_5_npc : _GEN_1420; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1422 = 3'h6 == deq_vec_1 ? buf_6_npc : _GEN_1421; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1425 = 3'h1 == deq_vec_1 ? buf_1_pc : buf_0_pc; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1426 = 3'h2 == deq_vec_1 ? buf_2_pc : _GEN_1425; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1427 = 3'h3 == deq_vec_1 ? buf_3_pc : _GEN_1426; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1428 = 3'h4 == deq_vec_1 ? buf_4_pc : _GEN_1427; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1429 = 3'h5 == deq_vec_1 ? buf_5_pc : _GEN_1428; // @[IssueUnit.scala 148:{15,15}]
  wire [31:0] _GEN_1430 = 3'h6 == deq_vec_1 ? buf_6_pc : _GEN_1429; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1433 = 3'h1 == deq_vec_1 ? buf_1_valid : buf_0_valid; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1434 = 3'h2 == deq_vec_1 ? buf_2_valid : _GEN_1433; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1435 = 3'h3 == deq_vec_1 ? buf_3_valid : _GEN_1434; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1436 = 3'h4 == deq_vec_1 ? buf_4_valid : _GEN_1435; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1437 = 3'h5 == deq_vec_1 ? buf_5_valid : _GEN_1436; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1438 = 3'h6 == deq_vec_1 ? buf_6_valid : _GEN_1437; // @[IssueUnit.scala 148:{15,15}]
  wire  _GEN_1439 = 3'h7 == deq_vec_1 ? buf_7_valid : _GEN_1438; // @[IssueUnit.scala 148:{15,15}]
  wire [2:0] _T_121 = deq_vec_1 - 3'h1; // @[IssueUnit.scala 161:34]
  wire  up2_0 = 3'h0 >= _T_121 & deq_vec_valid_1; // @[IssueUnit.scala 161:41]
  wire  up1_0 = 3'h0 >= deq_vec_0 & deq_vec_valid_0 & ~up2_0; // @[IssueUnit.scala 158:55]
  wire  up2_1 = 3'h1 >= _T_121 & deq_vec_valid_1; // @[IssueUnit.scala 161:41]
  wire  up1_1 = 3'h1 >= deq_vec_0 & deq_vec_valid_0 & ~up2_1; // @[IssueUnit.scala 158:55]
  wire  up2_2 = 3'h2 >= _T_121 & deq_vec_valid_1; // @[IssueUnit.scala 161:41]
  wire  up1_2 = 3'h2 >= deq_vec_0 & deq_vec_valid_0 & ~up2_2; // @[IssueUnit.scala 158:55]
  wire  up2_3 = 3'h3 >= _T_121 & deq_vec_valid_1; // @[IssueUnit.scala 161:41]
  wire  up1_3 = 3'h3 >= deq_vec_0 & deq_vec_valid_0 & ~up2_3; // @[IssueUnit.scala 158:55]
  wire  up2_4 = 3'h4 >= _T_121 & deq_vec_valid_1; // @[IssueUnit.scala 161:41]
  wire  up1_4 = 3'h4 >= deq_vec_0 & deq_vec_valid_0 & ~up2_4; // @[IssueUnit.scala 158:55]
  wire  up2_5 = 3'h5 >= _T_121 & deq_vec_valid_1; // @[IssueUnit.scala 161:41]
  wire  up1_5 = 3'h5 >= deq_vec_0 & deq_vec_valid_0 & ~up2_5; // @[IssueUnit.scala 158:55]
  wire  up2_6 = 3'h6 >= _T_121 & deq_vec_valid_1; // @[IssueUnit.scala 161:41]
  wire  up1_6 = 3'h6 >= deq_vec_0 & deq_vec_valid_0 & ~up2_6; // @[IssueUnit.scala 158:55]
  wire  up1_7 = deq_vec_valid_0 & ~deq_vec_valid_1; // @[IssueUnit.scala 158:55]
  wire [3:0] _GEN_1440 = up1_0 ? buf_1_rob_addr : buf_0_rob_addr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1442 = up1_0 ? buf_1_rd_paddr : buf_0_rd_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1443 = up1_0 ? buf_1_rs2_paddr : buf_0_rs2_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1444 = up1_0 ? buf_1_rs1_paddr : buf_0_rs1_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1445 = up1_0 ? buf_1_pred_bpc : buf_0_pred_bpc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1446 = up1_0 ? buf_1_pred_br : buf_0_pred_br; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1447 = up1_0 ? buf_1_imm : buf_0_imm; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1448 = up1_0 ? buf_1_rd_en : buf_0_rd_en; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [1:0] _GEN_1452 = up1_0 ? buf_1_rs2_src : buf_0_rs2_src; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [1:0] _GEN_1453 = up1_0 ? buf_1_rs1_src : buf_0_rs1_src; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1454 = up1_0 ? buf_1_w_type : buf_0_w_type; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [2:0] _GEN_1455 = up1_0 ? buf_1_sys_code : buf_0_sys_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1458 = up1_0 ? buf_1_jmp_code : buf_0_jmp_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1459 = up1_0 ? buf_1_alu_code : buf_0_alu_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [2:0] _GEN_1460 = up1_0 ? buf_1_fu_code : buf_0_fu_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1461 = up1_0 ? buf_1_inst : buf_0_inst; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1462 = up1_0 ? buf_1_npc : buf_0_npc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1463 = up1_0 ? buf_1_pc : buf_0_pc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1464 = up1_0 ? buf_1_valid : buf_0_valid; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1465 = up2_0 ? buf_2_rob_addr : _GEN_1440; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1467 = up2_0 ? buf_2_rd_paddr : _GEN_1442; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1468 = up2_0 ? buf_2_rs2_paddr : _GEN_1443; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1469 = up2_0 ? buf_2_rs1_paddr : _GEN_1444; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1470 = up2_0 ? buf_2_pred_bpc : _GEN_1445; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1471 = up2_0 ? buf_2_pred_br : _GEN_1446; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1472 = up2_0 ? buf_2_imm : _GEN_1447; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1473 = up2_0 ? buf_2_rd_en : _GEN_1448; // @[IssueUnit.scala 171:19 173:18]
  wire [1:0] _GEN_1477 = up2_0 ? buf_2_rs2_src : _GEN_1452; // @[IssueUnit.scala 171:19 173:18]
  wire [1:0] _GEN_1478 = up2_0 ? buf_2_rs1_src : _GEN_1453; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1479 = up2_0 ? buf_2_w_type : _GEN_1454; // @[IssueUnit.scala 171:19 173:18]
  wire [2:0] _GEN_1480 = up2_0 ? buf_2_sys_code : _GEN_1455; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1483 = up2_0 ? buf_2_jmp_code : _GEN_1458; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1484 = up2_0 ? buf_2_alu_code : _GEN_1459; // @[IssueUnit.scala 171:19 173:18]
  wire [2:0] _GEN_1485 = up2_0 ? buf_2_fu_code : _GEN_1460; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1486 = up2_0 ? buf_2_inst : _GEN_1461; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1487 = up2_0 ? buf_2_npc : _GEN_1462; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1488 = up2_0 ? buf_2_pc : _GEN_1463; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1489 = up2_0 ? buf_2_valid : _GEN_1464; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1490 = up1_1 ? buf_2_rob_addr : buf_1_rob_addr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1492 = up1_1 ? buf_2_rd_paddr : buf_1_rd_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1493 = up1_1 ? buf_2_rs2_paddr : buf_1_rs2_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1494 = up1_1 ? buf_2_rs1_paddr : buf_1_rs1_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1495 = up1_1 ? buf_2_pred_bpc : buf_1_pred_bpc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1496 = up1_1 ? buf_2_pred_br : buf_1_pred_br; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1497 = up1_1 ? buf_2_imm : buf_1_imm; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1498 = up1_1 ? buf_2_rd_en : buf_1_rd_en; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [1:0] _GEN_1502 = up1_1 ? buf_2_rs2_src : buf_1_rs2_src; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [1:0] _GEN_1503 = up1_1 ? buf_2_rs1_src : buf_1_rs1_src; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1504 = up1_1 ? buf_2_w_type : buf_1_w_type; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [2:0] _GEN_1505 = up1_1 ? buf_2_sys_code : buf_1_sys_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1508 = up1_1 ? buf_2_jmp_code : buf_1_jmp_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1509 = up1_1 ? buf_2_alu_code : buf_1_alu_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [2:0] _GEN_1510 = up1_1 ? buf_2_fu_code : buf_1_fu_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1511 = up1_1 ? buf_2_inst : buf_1_inst; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1512 = up1_1 ? buf_2_npc : buf_1_npc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1513 = up1_1 ? buf_2_pc : buf_1_pc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1514 = up1_1 ? buf_2_valid : buf_1_valid; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1515 = up2_1 ? buf_3_rob_addr : _GEN_1490; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1517 = up2_1 ? buf_3_rd_paddr : _GEN_1492; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1518 = up2_1 ? buf_3_rs2_paddr : _GEN_1493; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1519 = up2_1 ? buf_3_rs1_paddr : _GEN_1494; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1520 = up2_1 ? buf_3_pred_bpc : _GEN_1495; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1521 = up2_1 ? buf_3_pred_br : _GEN_1496; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1522 = up2_1 ? buf_3_imm : _GEN_1497; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1523 = up2_1 ? buf_3_rd_en : _GEN_1498; // @[IssueUnit.scala 171:19 173:18]
  wire [1:0] _GEN_1527 = up2_1 ? buf_3_rs2_src : _GEN_1502; // @[IssueUnit.scala 171:19 173:18]
  wire [1:0] _GEN_1528 = up2_1 ? buf_3_rs1_src : _GEN_1503; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1529 = up2_1 ? buf_3_w_type : _GEN_1504; // @[IssueUnit.scala 171:19 173:18]
  wire [2:0] _GEN_1530 = up2_1 ? buf_3_sys_code : _GEN_1505; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1533 = up2_1 ? buf_3_jmp_code : _GEN_1508; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1534 = up2_1 ? buf_3_alu_code : _GEN_1509; // @[IssueUnit.scala 171:19 173:18]
  wire [2:0] _GEN_1535 = up2_1 ? buf_3_fu_code : _GEN_1510; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1536 = up2_1 ? buf_3_inst : _GEN_1511; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1537 = up2_1 ? buf_3_npc : _GEN_1512; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1538 = up2_1 ? buf_3_pc : _GEN_1513; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1539 = up2_1 ? buf_3_valid : _GEN_1514; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1540 = up1_2 ? buf_3_rob_addr : buf_2_rob_addr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1542 = up1_2 ? buf_3_rd_paddr : buf_2_rd_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1543 = up1_2 ? buf_3_rs2_paddr : buf_2_rs2_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1544 = up1_2 ? buf_3_rs1_paddr : buf_2_rs1_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1545 = up1_2 ? buf_3_pred_bpc : buf_2_pred_bpc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1546 = up1_2 ? buf_3_pred_br : buf_2_pred_br; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1547 = up1_2 ? buf_3_imm : buf_2_imm; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1548 = up1_2 ? buf_3_rd_en : buf_2_rd_en; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [1:0] _GEN_1552 = up1_2 ? buf_3_rs2_src : buf_2_rs2_src; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [1:0] _GEN_1553 = up1_2 ? buf_3_rs1_src : buf_2_rs1_src; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1554 = up1_2 ? buf_3_w_type : buf_2_w_type; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [2:0] _GEN_1555 = up1_2 ? buf_3_sys_code : buf_2_sys_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1558 = up1_2 ? buf_3_jmp_code : buf_2_jmp_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1559 = up1_2 ? buf_3_alu_code : buf_2_alu_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [2:0] _GEN_1560 = up1_2 ? buf_3_fu_code : buf_2_fu_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1561 = up1_2 ? buf_3_inst : buf_2_inst; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1562 = up1_2 ? buf_3_npc : buf_2_npc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1563 = up1_2 ? buf_3_pc : buf_2_pc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1564 = up1_2 ? buf_3_valid : buf_2_valid; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1565 = up2_2 ? buf_4_rob_addr : _GEN_1540; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1567 = up2_2 ? buf_4_rd_paddr : _GEN_1542; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1568 = up2_2 ? buf_4_rs2_paddr : _GEN_1543; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1569 = up2_2 ? buf_4_rs1_paddr : _GEN_1544; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1570 = up2_2 ? buf_4_pred_bpc : _GEN_1545; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1571 = up2_2 ? buf_4_pred_br : _GEN_1546; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1572 = up2_2 ? buf_4_imm : _GEN_1547; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1573 = up2_2 ? buf_4_rd_en : _GEN_1548; // @[IssueUnit.scala 171:19 173:18]
  wire [1:0] _GEN_1577 = up2_2 ? buf_4_rs2_src : _GEN_1552; // @[IssueUnit.scala 171:19 173:18]
  wire [1:0] _GEN_1578 = up2_2 ? buf_4_rs1_src : _GEN_1553; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1579 = up2_2 ? buf_4_w_type : _GEN_1554; // @[IssueUnit.scala 171:19 173:18]
  wire [2:0] _GEN_1580 = up2_2 ? buf_4_sys_code : _GEN_1555; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1583 = up2_2 ? buf_4_jmp_code : _GEN_1558; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1584 = up2_2 ? buf_4_alu_code : _GEN_1559; // @[IssueUnit.scala 171:19 173:18]
  wire [2:0] _GEN_1585 = up2_2 ? buf_4_fu_code : _GEN_1560; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1586 = up2_2 ? buf_4_inst : _GEN_1561; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1587 = up2_2 ? buf_4_npc : _GEN_1562; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1588 = up2_2 ? buf_4_pc : _GEN_1563; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1589 = up2_2 ? buf_4_valid : _GEN_1564; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1590 = up1_3 ? buf_4_rob_addr : buf_3_rob_addr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1592 = up1_3 ? buf_4_rd_paddr : buf_3_rd_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1593 = up1_3 ? buf_4_rs2_paddr : buf_3_rs2_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1594 = up1_3 ? buf_4_rs1_paddr : buf_3_rs1_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1595 = up1_3 ? buf_4_pred_bpc : buf_3_pred_bpc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1596 = up1_3 ? buf_4_pred_br : buf_3_pred_br; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1597 = up1_3 ? buf_4_imm : buf_3_imm; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1598 = up1_3 ? buf_4_rd_en : buf_3_rd_en; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [1:0] _GEN_1602 = up1_3 ? buf_4_rs2_src : buf_3_rs2_src; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [1:0] _GEN_1603 = up1_3 ? buf_4_rs1_src : buf_3_rs1_src; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1604 = up1_3 ? buf_4_w_type : buf_3_w_type; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [2:0] _GEN_1605 = up1_3 ? buf_4_sys_code : buf_3_sys_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1608 = up1_3 ? buf_4_jmp_code : buf_3_jmp_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1609 = up1_3 ? buf_4_alu_code : buf_3_alu_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [2:0] _GEN_1610 = up1_3 ? buf_4_fu_code : buf_3_fu_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1611 = up1_3 ? buf_4_inst : buf_3_inst; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1612 = up1_3 ? buf_4_npc : buf_3_npc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1613 = up1_3 ? buf_4_pc : buf_3_pc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1614 = up1_3 ? buf_4_valid : buf_3_valid; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1615 = up2_3 ? buf_5_rob_addr : _GEN_1590; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1617 = up2_3 ? buf_5_rd_paddr : _GEN_1592; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1618 = up2_3 ? buf_5_rs2_paddr : _GEN_1593; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1619 = up2_3 ? buf_5_rs1_paddr : _GEN_1594; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1620 = up2_3 ? buf_5_pred_bpc : _GEN_1595; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1621 = up2_3 ? buf_5_pred_br : _GEN_1596; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1622 = up2_3 ? buf_5_imm : _GEN_1597; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1623 = up2_3 ? buf_5_rd_en : _GEN_1598; // @[IssueUnit.scala 171:19 173:18]
  wire [1:0] _GEN_1627 = up2_3 ? buf_5_rs2_src : _GEN_1602; // @[IssueUnit.scala 171:19 173:18]
  wire [1:0] _GEN_1628 = up2_3 ? buf_5_rs1_src : _GEN_1603; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1629 = up2_3 ? buf_5_w_type : _GEN_1604; // @[IssueUnit.scala 171:19 173:18]
  wire [2:0] _GEN_1630 = up2_3 ? buf_5_sys_code : _GEN_1605; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1633 = up2_3 ? buf_5_jmp_code : _GEN_1608; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1634 = up2_3 ? buf_5_alu_code : _GEN_1609; // @[IssueUnit.scala 171:19 173:18]
  wire [2:0] _GEN_1635 = up2_3 ? buf_5_fu_code : _GEN_1610; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1636 = up2_3 ? buf_5_inst : _GEN_1611; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1637 = up2_3 ? buf_5_npc : _GEN_1612; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1638 = up2_3 ? buf_5_pc : _GEN_1613; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1639 = up2_3 ? buf_5_valid : _GEN_1614; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1640 = up1_4 ? buf_5_rob_addr : buf_4_rob_addr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1642 = up1_4 ? buf_5_rd_paddr : buf_4_rd_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1643 = up1_4 ? buf_5_rs2_paddr : buf_4_rs2_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1644 = up1_4 ? buf_5_rs1_paddr : buf_4_rs1_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1645 = up1_4 ? buf_5_pred_bpc : buf_4_pred_bpc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1646 = up1_4 ? buf_5_pred_br : buf_4_pred_br; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1647 = up1_4 ? buf_5_imm : buf_4_imm; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1648 = up1_4 ? buf_5_rd_en : buf_4_rd_en; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [1:0] _GEN_1652 = up1_4 ? buf_5_rs2_src : buf_4_rs2_src; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [1:0] _GEN_1653 = up1_4 ? buf_5_rs1_src : buf_4_rs1_src; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1654 = up1_4 ? buf_5_w_type : buf_4_w_type; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [2:0] _GEN_1655 = up1_4 ? buf_5_sys_code : buf_4_sys_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1658 = up1_4 ? buf_5_jmp_code : buf_4_jmp_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1659 = up1_4 ? buf_5_alu_code : buf_4_alu_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [2:0] _GEN_1660 = up1_4 ? buf_5_fu_code : buf_4_fu_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1661 = up1_4 ? buf_5_inst : buf_4_inst; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1662 = up1_4 ? buf_5_npc : buf_4_npc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1663 = up1_4 ? buf_5_pc : buf_4_pc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1664 = up1_4 ? buf_5_valid : buf_4_valid; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1665 = up2_4 ? buf_6_rob_addr : _GEN_1640; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1667 = up2_4 ? buf_6_rd_paddr : _GEN_1642; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1668 = up2_4 ? buf_6_rs2_paddr : _GEN_1643; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1669 = up2_4 ? buf_6_rs1_paddr : _GEN_1644; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1670 = up2_4 ? buf_6_pred_bpc : _GEN_1645; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1671 = up2_4 ? buf_6_pred_br : _GEN_1646; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1672 = up2_4 ? buf_6_imm : _GEN_1647; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1673 = up2_4 ? buf_6_rd_en : _GEN_1648; // @[IssueUnit.scala 171:19 173:18]
  wire [1:0] _GEN_1677 = up2_4 ? buf_6_rs2_src : _GEN_1652; // @[IssueUnit.scala 171:19 173:18]
  wire [1:0] _GEN_1678 = up2_4 ? buf_6_rs1_src : _GEN_1653; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1679 = up2_4 ? buf_6_w_type : _GEN_1654; // @[IssueUnit.scala 171:19 173:18]
  wire [2:0] _GEN_1680 = up2_4 ? buf_6_sys_code : _GEN_1655; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1683 = up2_4 ? buf_6_jmp_code : _GEN_1658; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1684 = up2_4 ? buf_6_alu_code : _GEN_1659; // @[IssueUnit.scala 171:19 173:18]
  wire [2:0] _GEN_1685 = up2_4 ? buf_6_fu_code : _GEN_1660; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1686 = up2_4 ? buf_6_inst : _GEN_1661; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1687 = up2_4 ? buf_6_npc : _GEN_1662; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1688 = up2_4 ? buf_6_pc : _GEN_1663; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1689 = up2_4 ? buf_6_valid : _GEN_1664; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1690 = up1_5 ? buf_6_rob_addr : buf_5_rob_addr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1692 = up1_5 ? buf_6_rd_paddr : buf_5_rd_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1693 = up1_5 ? buf_6_rs2_paddr : buf_5_rs2_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1694 = up1_5 ? buf_6_rs1_paddr : buf_5_rs1_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1695 = up1_5 ? buf_6_pred_bpc : buf_5_pred_bpc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1696 = up1_5 ? buf_6_pred_br : buf_5_pred_br; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1697 = up1_5 ? buf_6_imm : buf_5_imm; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1698 = up1_5 ? buf_6_rd_en : buf_5_rd_en; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [1:0] _GEN_1702 = up1_5 ? buf_6_rs2_src : buf_5_rs2_src; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [1:0] _GEN_1703 = up1_5 ? buf_6_rs1_src : buf_5_rs1_src; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1704 = up1_5 ? buf_6_w_type : buf_5_w_type; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [2:0] _GEN_1705 = up1_5 ? buf_6_sys_code : buf_5_sys_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1708 = up1_5 ? buf_6_jmp_code : buf_5_jmp_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1709 = up1_5 ? buf_6_alu_code : buf_5_alu_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [2:0] _GEN_1710 = up1_5 ? buf_6_fu_code : buf_5_fu_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1711 = up1_5 ? buf_6_inst : buf_5_inst; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1712 = up1_5 ? buf_6_npc : buf_5_npc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1713 = up1_5 ? buf_6_pc : buf_5_pc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1714 = up1_5 ? buf_6_valid : buf_5_valid; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1715 = up2_5 ? buf_7_rob_addr : _GEN_1690; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1717 = up2_5 ? buf_7_rd_paddr : _GEN_1692; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1718 = up2_5 ? buf_7_rs2_paddr : _GEN_1693; // @[IssueUnit.scala 171:19 173:18]
  wire [5:0] _GEN_1719 = up2_5 ? buf_7_rs1_paddr : _GEN_1694; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1720 = up2_5 ? buf_7_pred_bpc : _GEN_1695; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1721 = up2_5 ? buf_7_pred_br : _GEN_1696; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1722 = up2_5 ? buf_7_imm : _GEN_1697; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1723 = up2_5 ? buf_7_rd_en : _GEN_1698; // @[IssueUnit.scala 171:19 173:18]
  wire [1:0] _GEN_1727 = up2_5 ? buf_7_rs2_src : _GEN_1702; // @[IssueUnit.scala 171:19 173:18]
  wire [1:0] _GEN_1728 = up2_5 ? buf_7_rs1_src : _GEN_1703; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1729 = up2_5 ? buf_7_w_type : _GEN_1704; // @[IssueUnit.scala 171:19 173:18]
  wire [2:0] _GEN_1730 = up2_5 ? buf_7_sys_code : _GEN_1705; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1733 = up2_5 ? buf_7_jmp_code : _GEN_1708; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1734 = up2_5 ? buf_7_alu_code : _GEN_1709; // @[IssueUnit.scala 171:19 173:18]
  wire [2:0] _GEN_1735 = up2_5 ? buf_7_fu_code : _GEN_1710; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1736 = up2_5 ? buf_7_inst : _GEN_1711; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1737 = up2_5 ? buf_7_npc : _GEN_1712; // @[IssueUnit.scala 171:19 173:18]
  wire [31:0] _GEN_1738 = up2_5 ? buf_7_pc : _GEN_1713; // @[IssueUnit.scala 171:19 173:18]
  wire  _GEN_1739 = up2_5 ? buf_7_valid : _GEN_1714; // @[IssueUnit.scala 171:19 173:18]
  wire [3:0] _GEN_1740 = up1_6 ? buf_7_rob_addr : buf_6_rob_addr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1742 = up1_6 ? buf_7_rd_paddr : buf_6_rd_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1743 = up1_6 ? buf_7_rs2_paddr : buf_6_rs2_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [5:0] _GEN_1744 = up1_6 ? buf_7_rs1_paddr : buf_6_rs1_paddr; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1745 = up1_6 ? buf_7_pred_bpc : buf_6_pred_bpc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1746 = up1_6 ? buf_7_pred_br : buf_6_pred_br; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1747 = up1_6 ? buf_7_imm : buf_6_imm; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1748 = up1_6 ? buf_7_rd_en : buf_6_rd_en; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [1:0] _GEN_1752 = up1_6 ? buf_7_rs2_src : buf_6_rs2_src; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [1:0] _GEN_1753 = up1_6 ? buf_7_rs1_src : buf_6_rs1_src; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1754 = up1_6 ? buf_7_w_type : buf_6_w_type; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [2:0] _GEN_1755 = up1_6 ? buf_7_sys_code : buf_6_sys_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1758 = up1_6 ? buf_7_jmp_code : buf_6_jmp_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1759 = up1_6 ? buf_7_alu_code : buf_6_alu_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [2:0] _GEN_1760 = up1_6 ? buf_7_fu_code : buf_6_fu_code; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1761 = up1_6 ? buf_7_inst : buf_6_inst; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1762 = up1_6 ? buf_7_npc : buf_6_npc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [31:0] _GEN_1763 = up1_6 ? buf_7_pc : buf_6_pc; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire  _GEN_1764 = up1_6 ? buf_7_valid : buf_6_valid; // @[IssueUnit.scala 164:19 166:18 97:20]
  wire [3:0] _GEN_1765 = up2_6 ? 4'h0 : _GEN_1740; // @[IssueUnit.scala 171:19 175:18]
  wire [5:0] _GEN_1767 = up2_6 ? 6'h0 : _GEN_1742; // @[IssueUnit.scala 171:19 175:18]
  wire [5:0] _GEN_1768 = up2_6 ? 6'h0 : _GEN_1743; // @[IssueUnit.scala 171:19 175:18]
  wire [5:0] _GEN_1769 = up2_6 ? 6'h0 : _GEN_1744; // @[IssueUnit.scala 171:19 175:18]
  wire [31:0] _GEN_1770 = up2_6 ? 32'h0 : _GEN_1745; // @[IssueUnit.scala 171:19 175:18]
  wire  _GEN_1771 = up2_6 ? 1'h0 : _GEN_1746; // @[IssueUnit.scala 171:19 175:18]
  wire [31:0] _GEN_1772 = up2_6 ? 32'h0 : _GEN_1747; // @[IssueUnit.scala 171:19 175:18]
  wire  _GEN_1773 = up2_6 ? 1'h0 : _GEN_1748; // @[IssueUnit.scala 171:19 175:18]
  wire [1:0] _GEN_1777 = up2_6 ? 2'h0 : _GEN_1752; // @[IssueUnit.scala 171:19 175:18]
  wire [1:0] _GEN_1778 = up2_6 ? 2'h0 : _GEN_1753; // @[IssueUnit.scala 171:19 175:18]
  wire  _GEN_1779 = up2_6 ? 1'h0 : _GEN_1754; // @[IssueUnit.scala 171:19 175:18]
  wire [2:0] _GEN_1780 = up2_6 ? 3'h0 : _GEN_1755; // @[IssueUnit.scala 171:19 175:18]
  wire [3:0] _GEN_1783 = up2_6 ? 4'h0 : _GEN_1758; // @[IssueUnit.scala 171:19 175:18]
  wire [3:0] _GEN_1784 = up2_6 ? 4'h0 : _GEN_1759; // @[IssueUnit.scala 171:19 175:18]
  wire [2:0] _GEN_1785 = up2_6 ? 3'h0 : _GEN_1760; // @[IssueUnit.scala 171:19 175:18]
  wire [31:0] _GEN_1786 = up2_6 ? 32'h0 : _GEN_1761; // @[IssueUnit.scala 171:19 175:18]
  wire [31:0] _GEN_1787 = up2_6 ? 32'h0 : _GEN_1762; // @[IssueUnit.scala 171:19 175:18]
  wire [31:0] _GEN_1788 = up2_6 ? 32'h0 : _GEN_1763; // @[IssueUnit.scala 171:19 175:18]
  wire  _GEN_1789 = up2_6 ? 1'h0 : _GEN_1764; // @[IssueUnit.scala 171:19 175:18]
  wire [3:0] _GEN_1790 = up1_7 ? 4'h0 : buf_7_rob_addr; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [5:0] _GEN_1792 = up1_7 ? 6'h0 : buf_7_rd_paddr; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [5:0] _GEN_1793 = up1_7 ? 6'h0 : buf_7_rs2_paddr; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [5:0] _GEN_1794 = up1_7 ? 6'h0 : buf_7_rs1_paddr; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [31:0] _GEN_1795 = up1_7 ? 32'h0 : buf_7_pred_bpc; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire  _GEN_1796 = up1_7 ? 1'h0 : buf_7_pred_br; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [31:0] _GEN_1797 = up1_7 ? 32'h0 : buf_7_imm; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire  _GEN_1798 = up1_7 ? 1'h0 : buf_7_rd_en; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [1:0] _GEN_1802 = up1_7 ? 2'h0 : buf_7_rs2_src; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [1:0] _GEN_1803 = up1_7 ? 2'h0 : buf_7_rs1_src; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire  _GEN_1804 = up1_7 ? 1'h0 : buf_7_w_type; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [2:0] _GEN_1805 = up1_7 ? 3'h0 : buf_7_sys_code; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [3:0] _GEN_1808 = up1_7 ? 4'h0 : buf_7_jmp_code; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [3:0] _GEN_1809 = up1_7 ? 4'h0 : buf_7_alu_code; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [2:0] _GEN_1810 = up1_7 ? 3'h0 : buf_7_fu_code; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [31:0] _GEN_1811 = up1_7 ? 32'h0 : buf_7_inst; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [31:0] _GEN_1812 = up1_7 ? 32'h0 : buf_7_npc; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [31:0] _GEN_1813 = up1_7 ? 32'h0 : buf_7_pc; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire  _GEN_1814 = up1_7 ? 1'h0 : buf_7_valid; // @[IssueUnit.scala 164:19 168:18 97:20]
  wire [3:0] _GEN_1815 = deq_vec_valid_1 ? 4'h0 : _GEN_1790; // @[IssueUnit.scala 171:19 175:18]
  wire [5:0] _GEN_1817 = deq_vec_valid_1 ? 6'h0 : _GEN_1792; // @[IssueUnit.scala 171:19 175:18]
  wire [5:0] _GEN_1818 = deq_vec_valid_1 ? 6'h0 : _GEN_1793; // @[IssueUnit.scala 171:19 175:18]
  wire [5:0] _GEN_1819 = deq_vec_valid_1 ? 6'h0 : _GEN_1794; // @[IssueUnit.scala 171:19 175:18]
  wire [31:0] _GEN_1820 = deq_vec_valid_1 ? 32'h0 : _GEN_1795; // @[IssueUnit.scala 171:19 175:18]
  wire  _GEN_1821 = deq_vec_valid_1 ? 1'h0 : _GEN_1796; // @[IssueUnit.scala 171:19 175:18]
  wire [31:0] _GEN_1822 = deq_vec_valid_1 ? 32'h0 : _GEN_1797; // @[IssueUnit.scala 171:19 175:18]
  wire  _GEN_1823 = deq_vec_valid_1 ? 1'h0 : _GEN_1798; // @[IssueUnit.scala 171:19 175:18]
  wire [1:0] _GEN_1827 = deq_vec_valid_1 ? 2'h0 : _GEN_1802; // @[IssueUnit.scala 171:19 175:18]
  wire [1:0] _GEN_1828 = deq_vec_valid_1 ? 2'h0 : _GEN_1803; // @[IssueUnit.scala 171:19 175:18]
  wire  _GEN_1829 = deq_vec_valid_1 ? 1'h0 : _GEN_1804; // @[IssueUnit.scala 171:19 175:18]
  wire [2:0] _GEN_1830 = deq_vec_valid_1 ? 3'h0 : _GEN_1805; // @[IssueUnit.scala 171:19 175:18]
  wire [3:0] _GEN_1833 = deq_vec_valid_1 ? 4'h0 : _GEN_1808; // @[IssueUnit.scala 171:19 175:18]
  wire [3:0] _GEN_1834 = deq_vec_valid_1 ? 4'h0 : _GEN_1809; // @[IssueUnit.scala 171:19 175:18]
  wire [2:0] _GEN_1835 = deq_vec_valid_1 ? 3'h0 : _GEN_1810; // @[IssueUnit.scala 171:19 175:18]
  wire [31:0] _GEN_1836 = deq_vec_valid_1 ? 32'h0 : _GEN_1811; // @[IssueUnit.scala 171:19 175:18]
  wire [31:0] _GEN_1837 = deq_vec_valid_1 ? 32'h0 : _GEN_1812; // @[IssueUnit.scala 171:19 175:18]
  wire [31:0] _GEN_1838 = deq_vec_valid_1 ? 32'h0 : _GEN_1813; // @[IssueUnit.scala 171:19 175:18]
  wire  _GEN_1839 = deq_vec_valid_1 ? 1'h0 : _GEN_1814; // @[IssueUnit.scala 171:19 175:18]
  wire  _T_155 = ~io_flush; // @[IssueUnit.scala 197:40]
  wire [3:0] _GEN_1842 = 3'h0 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1465; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1843 = 3'h1 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1515; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1844 = 3'h2 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1565; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1845 = 3'h3 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1615; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1846 = 3'h4 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1665; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1847 = 3'h5 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1715; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1848 = 3'h6 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1765; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1849 = 3'h7 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1815; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1858 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1467; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1859 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1517; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1860 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1567; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1861 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1617; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1862 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1667; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1863 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1717; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1864 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1767; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1865 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1817; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1866 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1468; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1867 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1518; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1868 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1568; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1869 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1618; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1870 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1668; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1871 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1718; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1872 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1768; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1873 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1818; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1874 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1469; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1875 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1519; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1876 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1569; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1877 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1619; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1878 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1669; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1879 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1719; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1880 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1769; // @[IssueUnit.scala 198:{48,48}]
  wire [5:0] _GEN_1881 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1819; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1882 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_bpc : _GEN_1470; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1883 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_bpc : _GEN_1520; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1884 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_bpc : _GEN_1570; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1885 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_bpc : _GEN_1620; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1886 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_bpc : _GEN_1670; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1887 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_bpc : _GEN_1720; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1888 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_bpc : _GEN_1770; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1889 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_bpc : _GEN_1820; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1890 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_br : _GEN_1471; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1891 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_br : _GEN_1521; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1892 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_br : _GEN_1571; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1893 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_br : _GEN_1621; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1894 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_br : _GEN_1671; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1895 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_br : _GEN_1721; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1896 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_br : _GEN_1771; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1897 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pred_br : _GEN_1821; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1898 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1472; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1899 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1522; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1900 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1572; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1901 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1622; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1902 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1672; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1903 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1722; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1904 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1772; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_1905 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1822; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1906 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1473; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1907 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1523; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1908 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1573; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1909 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1623; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1910 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1673; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1911 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1723; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1912 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1773; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1913 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1823; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1938 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1477; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1939 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1527; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1940 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1577; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1941 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1627; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1942 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1677; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1943 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1727; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1944 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1777; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1945 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1827; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1946 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1478; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1947 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1528; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1948 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1578; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1949 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1628; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1950 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1678; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1951 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1728; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1952 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1778; // @[IssueUnit.scala 198:{48,48}]
  wire [1:0] _GEN_1953 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1828; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1954 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1479; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1955 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1529; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1956 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1579; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1957 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1629; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1958 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1679; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1959 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1729; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1960 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1779; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_1961 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1829; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_1962 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_sys_code : _GEN_1480; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_1963 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_sys_code : _GEN_1530; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_1964 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_sys_code : _GEN_1580; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_1965 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_sys_code : _GEN_1630; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_1966 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_sys_code : _GEN_1680; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_1967 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_sys_code : _GEN_1730; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_1968 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_sys_code : _GEN_1780; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_1969 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_sys_code : _GEN_1830; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1986 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_jmp_code : _GEN_1483; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1987 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_jmp_code : _GEN_1533; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1988 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_jmp_code : _GEN_1583; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1989 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_jmp_code : _GEN_1633; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1990 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_jmp_code : _GEN_1683; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1991 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_jmp_code : _GEN_1733; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1992 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_jmp_code : _GEN_1783; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1993 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_jmp_code : _GEN_1833; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1994 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1484; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1995 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1534; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1996 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1584; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1997 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1634; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1998 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1684; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_1999 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1734; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_2000 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1784; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_2001 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1834; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_2002 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1485; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_2003 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1535; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_2004 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1585; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_2005 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1635; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_2006 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1685; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_2007 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1735; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_2008 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1785; // @[IssueUnit.scala 198:{48,48}]
  wire [2:0] _GEN_2009 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1835; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2010 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_inst : _GEN_1486; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2011 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_inst : _GEN_1536; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2012 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_inst : _GEN_1586; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2013 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_inst : _GEN_1636; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2014 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_inst : _GEN_1686; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2015 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_inst : _GEN_1736; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2016 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_inst : _GEN_1786; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2017 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_inst : _GEN_1836; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2018 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_npc : _GEN_1487; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2019 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_npc : _GEN_1537; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2020 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_npc : _GEN_1587; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2021 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_npc : _GEN_1637; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2022 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_npc : _GEN_1687; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2023 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_npc : _GEN_1737; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2024 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_npc : _GEN_1787; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2025 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_npc : _GEN_1837; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2026 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1488; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2027 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1538; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2028 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1588; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2029 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1638; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2030 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1688; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2031 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1738; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2032 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1788; // @[IssueUnit.scala 198:{48,48}]
  wire [31:0] _GEN_2033 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1838; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_2034 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1489; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_2035 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1539; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_2036 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1589; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_2037 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1639; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_2038 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1689; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_2039 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1739; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_2040 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1789; // @[IssueUnit.scala 198:{48,48}]
  wire  _GEN_2041 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1839; // @[IssueUnit.scala 198:{48,48}]
  wire [3:0] _GEN_2042 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1842 : _GEN_1465; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2043 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1843 : _GEN_1515; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2044 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1844 : _GEN_1565; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2045 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1845 : _GEN_1615; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2046 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1846 : _GEN_1665; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2047 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1847 : _GEN_1715; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2048 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1848 : _GEN_1765; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2049 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1849 : _GEN_1815; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2058 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1858 : _GEN_1467; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2059 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1859 : _GEN_1517; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2060 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1860 : _GEN_1567; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2061 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1861 : _GEN_1617; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2062 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1862 : _GEN_1667; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2063 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1863 : _GEN_1717; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2064 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1864 : _GEN_1767; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2065 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1865 : _GEN_1817; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2066 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1866 : _GEN_1468; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2067 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1867 : _GEN_1518; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2068 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1868 : _GEN_1568; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2069 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1869 : _GEN_1618; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2070 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1870 : _GEN_1668; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2071 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1871 : _GEN_1718; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2072 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1872 : _GEN_1768; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2073 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1873 : _GEN_1818; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2074 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1874 : _GEN_1469; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2075 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1875 : _GEN_1519; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2076 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1876 : _GEN_1569; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2077 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1877 : _GEN_1619; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2078 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1878 : _GEN_1669; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2079 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1879 : _GEN_1719; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2080 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1880 : _GEN_1769; // @[IssueUnit.scala 197:51]
  wire [5:0] _GEN_2081 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1881 : _GEN_1819; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2082 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1882 : _GEN_1470; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2083 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1883 : _GEN_1520; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2084 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1884 : _GEN_1570; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2085 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1885 : _GEN_1620; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2086 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1886 : _GEN_1670; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2087 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1887 : _GEN_1720; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2088 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1888 : _GEN_1770; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2089 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1889 : _GEN_1820; // @[IssueUnit.scala 197:51]
  wire  _GEN_2090 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1890 : _GEN_1471; // @[IssueUnit.scala 197:51]
  wire  _GEN_2091 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1891 : _GEN_1521; // @[IssueUnit.scala 197:51]
  wire  _GEN_2092 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1892 : _GEN_1571; // @[IssueUnit.scala 197:51]
  wire  _GEN_2093 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1893 : _GEN_1621; // @[IssueUnit.scala 197:51]
  wire  _GEN_2094 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1894 : _GEN_1671; // @[IssueUnit.scala 197:51]
  wire  _GEN_2095 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1895 : _GEN_1721; // @[IssueUnit.scala 197:51]
  wire  _GEN_2096 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1896 : _GEN_1771; // @[IssueUnit.scala 197:51]
  wire  _GEN_2097 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1897 : _GEN_1821; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2098 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1898 : _GEN_1472; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2099 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1899 : _GEN_1522; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2100 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1900 : _GEN_1572; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2101 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1901 : _GEN_1622; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2102 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1902 : _GEN_1672; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2103 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1903 : _GEN_1722; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2104 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1904 : _GEN_1772; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2105 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1905 : _GEN_1822; // @[IssueUnit.scala 197:51]
  wire  _GEN_2106 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1906 : _GEN_1473; // @[IssueUnit.scala 197:51]
  wire  _GEN_2107 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1907 : _GEN_1523; // @[IssueUnit.scala 197:51]
  wire  _GEN_2108 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1908 : _GEN_1573; // @[IssueUnit.scala 197:51]
  wire  _GEN_2109 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1909 : _GEN_1623; // @[IssueUnit.scala 197:51]
  wire  _GEN_2110 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1910 : _GEN_1673; // @[IssueUnit.scala 197:51]
  wire  _GEN_2111 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1911 : _GEN_1723; // @[IssueUnit.scala 197:51]
  wire  _GEN_2112 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1912 : _GEN_1773; // @[IssueUnit.scala 197:51]
  wire  _GEN_2113 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1913 : _GEN_1823; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2138 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1938 : _GEN_1477; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2139 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1939 : _GEN_1527; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2140 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1940 : _GEN_1577; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2141 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1941 : _GEN_1627; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2142 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1942 : _GEN_1677; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2143 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1943 : _GEN_1727; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2144 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1944 : _GEN_1777; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2145 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1945 : _GEN_1827; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2146 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1946 : _GEN_1478; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2147 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1947 : _GEN_1528; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2148 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1948 : _GEN_1578; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2149 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1949 : _GEN_1628; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2150 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1950 : _GEN_1678; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2151 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1951 : _GEN_1728; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2152 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1952 : _GEN_1778; // @[IssueUnit.scala 197:51]
  wire [1:0] _GEN_2153 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1953 : _GEN_1828; // @[IssueUnit.scala 197:51]
  wire  _GEN_2154 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1954 : _GEN_1479; // @[IssueUnit.scala 197:51]
  wire  _GEN_2155 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1955 : _GEN_1529; // @[IssueUnit.scala 197:51]
  wire  _GEN_2156 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1956 : _GEN_1579; // @[IssueUnit.scala 197:51]
  wire  _GEN_2157 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1957 : _GEN_1629; // @[IssueUnit.scala 197:51]
  wire  _GEN_2158 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1958 : _GEN_1679; // @[IssueUnit.scala 197:51]
  wire  _GEN_2159 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1959 : _GEN_1729; // @[IssueUnit.scala 197:51]
  wire  _GEN_2160 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1960 : _GEN_1779; // @[IssueUnit.scala 197:51]
  wire  _GEN_2161 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1961 : _GEN_1829; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2162 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1962 : _GEN_1480; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2163 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1963 : _GEN_1530; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2164 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1964 : _GEN_1580; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2165 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1965 : _GEN_1630; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2166 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1966 : _GEN_1680; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2167 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1967 : _GEN_1730; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2168 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1968 : _GEN_1780; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2169 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1969 : _GEN_1830; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2186 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1986 : _GEN_1483; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2187 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1987 : _GEN_1533; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2188 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1988 : _GEN_1583; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2189 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1989 : _GEN_1633; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2190 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1990 : _GEN_1683; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2191 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1991 : _GEN_1733; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2192 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1992 : _GEN_1783; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2193 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1993 : _GEN_1833; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2194 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1994 : _GEN_1484; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2195 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1995 : _GEN_1534; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2196 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1996 : _GEN_1584; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2197 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1997 : _GEN_1634; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2198 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1998 : _GEN_1684; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2199 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1999 : _GEN_1734; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2200 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2000 : _GEN_1784; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2201 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2001 : _GEN_1834; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2202 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2002 : _GEN_1485; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2203 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2003 : _GEN_1535; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2204 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2004 : _GEN_1585; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2205 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2005 : _GEN_1635; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2206 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2006 : _GEN_1685; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2207 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2007 : _GEN_1735; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2208 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2008 : _GEN_1785; // @[IssueUnit.scala 197:51]
  wire [2:0] _GEN_2209 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2009 : _GEN_1835; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2210 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2010 : _GEN_1486; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2211 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2011 : _GEN_1536; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2212 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2012 : _GEN_1586; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2213 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2013 : _GEN_1636; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2214 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2014 : _GEN_1686; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2215 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2015 : _GEN_1736; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2216 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2016 : _GEN_1786; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2217 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2017 : _GEN_1836; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2218 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2018 : _GEN_1487; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2219 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2019 : _GEN_1537; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2220 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2020 : _GEN_1587; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2221 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2021 : _GEN_1637; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2222 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2022 : _GEN_1687; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2223 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2023 : _GEN_1737; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2224 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2024 : _GEN_1787; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2225 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2025 : _GEN_1837; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2226 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2026 : _GEN_1488; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2227 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2027 : _GEN_1538; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2228 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2028 : _GEN_1588; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2229 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2029 : _GEN_1638; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2230 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2030 : _GEN_1688; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2231 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2031 : _GEN_1738; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2232 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2032 : _GEN_1788; // @[IssueUnit.scala 197:51]
  wire [31:0] _GEN_2233 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2033 : _GEN_1838; // @[IssueUnit.scala 197:51]
  wire  _GEN_2234 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2034 : _GEN_1489; // @[IssueUnit.scala 197:51]
  wire  _GEN_2235 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2035 : _GEN_1539; // @[IssueUnit.scala 197:51]
  wire  _GEN_2236 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2036 : _GEN_1589; // @[IssueUnit.scala 197:51]
  wire  _GEN_2237 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2037 : _GEN_1639; // @[IssueUnit.scala 197:51]
  wire  _GEN_2238 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2038 : _GEN_1689; // @[IssueUnit.scala 197:51]
  wire  _GEN_2239 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2039 : _GEN_1739; // @[IssueUnit.scala 197:51]
  wire  _GEN_2240 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2040 : _GEN_1789; // @[IssueUnit.scala 197:51]
  wire  _GEN_2241 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_2041 : _GEN_1839; // @[IssueUnit.scala 197:51]
  wire [3:0] _GEN_2243 = io_in_bits_vec_0_valid ? enq_vec_real_1 : enq_vec_real_0; // @[IssueUnit.scala 95:{32,32}]
  wire [3:0] _GEN_2850 = {{2'd0}, num_enq}; // @[IssueUnit.scala 202:44]
  wire [3:0] _T_164 = enq_vec_0 + _GEN_2850; // @[IssueUnit.scala 202:44]
  wire [3:0] next_enq_vec_0 = _T_164 - _GEN_2848; // @[IssueUnit.scala 202:54]
  wire [3:0] _T_168 = enq_vec_1 + _GEN_2850; // @[IssueUnit.scala 202:44]
  wire [3:0] next_enq_vec_1 = _T_168 - _GEN_2848; // @[IssueUnit.scala 202:54]
  wire [1:0] _T_172 = {io_out_0_valid,io_out_1_valid}; // @[Cat.scala 30:58]
  assign io_in_ready = enq_ready & ~has_sys; // @[IssueUnit.scala 208:28]
  assign io_out_0_valid = _GEN_1239 & deq_vec_valid_0; // @[IssueUnit.scala 149:34]
  assign io_out_0_pc = 3'h7 == deq_vec_0 ? buf_7_pc : _GEN_1230; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_npc = 3'h7 == deq_vec_0 ? buf_7_npc : _GEN_1222; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_inst = 3'h7 == deq_vec_0 ? buf_7_inst : _GEN_1214; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_fu_code = 3'h7 == deq_vec_0 ? buf_7_fu_code : _GEN_1206; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_alu_code = 3'h7 == deq_vec_0 ? buf_7_alu_code : _GEN_1198; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_jmp_code = 3'h7 == deq_vec_0 ? buf_7_jmp_code : _GEN_1190; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_sys_code = 3'h7 == deq_vec_0 ? buf_7_sys_code : _GEN_1166; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_w_type = 3'h7 == deq_vec_0 ? buf_7_w_type : _GEN_1158; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_rs1_src = 3'h7 == deq_vec_0 ? buf_7_rs1_src : _GEN_1150; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_rs2_src = 3'h7 == deq_vec_0 ? buf_7_rs2_src : _GEN_1142; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_rd_en = 3'h7 == deq_vec_0 ? buf_7_rd_en : _GEN_1110; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_imm = 3'h7 == deq_vec_0 ? buf_7_imm : _GEN_1102; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_pred_br = 3'h7 == deq_vec_0 ? buf_7_pred_br : _GEN_1094; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_pred_bpc = 3'h7 == deq_vec_0 ? buf_7_pred_bpc : _GEN_1086; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_rs1_paddr = 3'h7 == deq_vec_0 ? buf_7_rs1_paddr : _GEN_1078; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_rs2_paddr = 3'h7 == deq_vec_0 ? buf_7_rs2_paddr : _GEN_1070; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_rd_paddr = 3'h7 == deq_vec_0 ? buf_7_rd_paddr : _GEN_1062; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_0_rob_addr = 3'h7 == deq_vec_0 ? buf_7_rob_addr : _GEN_1046; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_valid = _GEN_1439 & deq_vec_valid_1; // @[IssueUnit.scala 149:34]
  assign io_out_1_pc = 3'h7 == deq_vec_1 ? buf_7_pc : _GEN_1430; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_npc = 3'h7 == deq_vec_1 ? buf_7_npc : _GEN_1422; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_fu_code = 3'h7 == deq_vec_1 ? buf_7_fu_code : _GEN_1406; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_alu_code = 3'h7 == deq_vec_1 ? buf_7_alu_code : _GEN_1398; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_jmp_code = 3'h7 == deq_vec_1 ? buf_7_jmp_code : _GEN_1390; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_w_type = 3'h7 == deq_vec_1 ? buf_7_w_type : _GEN_1358; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_rs1_src = 3'h7 == deq_vec_1 ? buf_7_rs1_src : _GEN_1350; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_rs2_src = 3'h7 == deq_vec_1 ? buf_7_rs2_src : _GEN_1342; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_rd_en = 3'h7 == deq_vec_1 ? buf_7_rd_en : _GEN_1310; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_imm = 3'h7 == deq_vec_1 ? buf_7_imm : _GEN_1302; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_pred_br = 3'h7 == deq_vec_1 ? buf_7_pred_br : _GEN_1294; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_pred_bpc = 3'h7 == deq_vec_1 ? buf_7_pred_bpc : _GEN_1286; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_rs1_paddr = 3'h7 == deq_vec_1 ? buf_7_rs1_paddr : _GEN_1278; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_rs2_paddr = 3'h7 == deq_vec_1 ? buf_7_rs2_paddr : _GEN_1270; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_rd_paddr = 3'h7 == deq_vec_1 ? buf_7_rd_paddr : _GEN_1262; // @[IssueUnit.scala 148:{15,15}]
  assign io_out_1_rob_addr = 3'h7 == deq_vec_1 ? buf_7_rob_addr : _GEN_1246; // @[IssueUnit.scala 148:{15,15}]
  always @(posedge clock) begin
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_valid <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_valid <= _GEN_2234;
      end
    end else begin
      buf_0_valid <= _GEN_2234;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_pc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_pc <= _GEN_2226;
      end
    end else begin
      buf_0_pc <= _GEN_2226;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_npc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_npc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_npc <= io_in_bits_vec_1_npc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_npc <= _GEN_2218;
      end
    end else begin
      buf_0_npc <= _GEN_2218;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_inst <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_inst <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_inst <= io_in_bits_vec_1_inst; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_inst <= _GEN_2210;
      end
    end else begin
      buf_0_inst <= _GEN_2210;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_fu_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_fu_code <= _GEN_2202;
      end
    end else begin
      buf_0_fu_code <= _GEN_2202;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_alu_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_alu_code <= _GEN_2194;
      end
    end else begin
      buf_0_alu_code <= _GEN_2194;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_jmp_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_jmp_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_jmp_code <= io_in_bits_vec_1_jmp_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_jmp_code <= _GEN_2186;
      end
    end else begin
      buf_0_jmp_code <= _GEN_2186;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_sys_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_sys_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_sys_code <= io_in_bits_vec_1_sys_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_sys_code <= _GEN_2162;
      end
    end else begin
      buf_0_sys_code <= _GEN_2162;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_w_type <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_w_type <= _GEN_2154;
      end
    end else begin
      buf_0_w_type <= _GEN_2154;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_rs1_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_rs1_src <= _GEN_2146;
      end
    end else begin
      buf_0_rs1_src <= _GEN_2146;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_rs2_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_rs2_src <= _GEN_2138;
      end
    end else begin
      buf_0_rs2_src <= _GEN_2138;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_rd_en <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_rd_en <= _GEN_2106;
      end
    end else begin
      buf_0_rd_en <= _GEN_2106;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_imm <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_imm <= _GEN_2098;
      end
    end else begin
      buf_0_imm <= _GEN_2098;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_pred_br <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_pred_br <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_pred_br <= io_in_bits_vec_1_pred_br; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_pred_br <= _GEN_2090;
      end
    end else begin
      buf_0_pred_br <= _GEN_2090;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_pred_bpc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_pred_bpc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_pred_bpc <= io_in_bits_vec_1_pred_bpc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_pred_bpc <= _GEN_2082;
      end
    end else begin
      buf_0_pred_bpc <= _GEN_2082;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_rs1_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_rs1_paddr <= _GEN_2074;
      end
    end else begin
      buf_0_rs1_paddr <= _GEN_2074;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_rs2_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_rs2_paddr <= _GEN_2066;
      end
    end else begin
      buf_0_rs2_paddr <= _GEN_2066;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_rd_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_rd_paddr <= _GEN_2058;
      end
    end else begin
      buf_0_rd_paddr <= _GEN_2058;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_0_rob_addr <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h0 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_0_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 198:48]
      end else begin
        buf_0_rob_addr <= _GEN_2042;
      end
    end else begin
      buf_0_rob_addr <= _GEN_2042;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_valid <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_valid <= _GEN_2235;
      end
    end else begin
      buf_1_valid <= _GEN_2235;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_pc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_pc <= _GEN_2227;
      end
    end else begin
      buf_1_pc <= _GEN_2227;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_npc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_npc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_npc <= io_in_bits_vec_1_npc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_npc <= _GEN_2219;
      end
    end else begin
      buf_1_npc <= _GEN_2219;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_inst <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_inst <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_inst <= io_in_bits_vec_1_inst; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_inst <= _GEN_2211;
      end
    end else begin
      buf_1_inst <= _GEN_2211;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_fu_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_fu_code <= _GEN_2203;
      end
    end else begin
      buf_1_fu_code <= _GEN_2203;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_alu_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_alu_code <= _GEN_2195;
      end
    end else begin
      buf_1_alu_code <= _GEN_2195;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_jmp_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_jmp_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_jmp_code <= io_in_bits_vec_1_jmp_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_jmp_code <= _GEN_2187;
      end
    end else begin
      buf_1_jmp_code <= _GEN_2187;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_sys_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_sys_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_sys_code <= io_in_bits_vec_1_sys_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_sys_code <= _GEN_2163;
      end
    end else begin
      buf_1_sys_code <= _GEN_2163;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_w_type <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_w_type <= _GEN_2155;
      end
    end else begin
      buf_1_w_type <= _GEN_2155;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_rs1_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_rs1_src <= _GEN_2147;
      end
    end else begin
      buf_1_rs1_src <= _GEN_2147;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_rs2_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_rs2_src <= _GEN_2139;
      end
    end else begin
      buf_1_rs2_src <= _GEN_2139;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_rd_en <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_rd_en <= _GEN_2107;
      end
    end else begin
      buf_1_rd_en <= _GEN_2107;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_imm <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_imm <= _GEN_2099;
      end
    end else begin
      buf_1_imm <= _GEN_2099;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_pred_br <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_pred_br <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_pred_br <= io_in_bits_vec_1_pred_br; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_pred_br <= _GEN_2091;
      end
    end else begin
      buf_1_pred_br <= _GEN_2091;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_pred_bpc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_pred_bpc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_pred_bpc <= io_in_bits_vec_1_pred_bpc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_pred_bpc <= _GEN_2083;
      end
    end else begin
      buf_1_pred_bpc <= _GEN_2083;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_rs1_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_rs1_paddr <= _GEN_2075;
      end
    end else begin
      buf_1_rs1_paddr <= _GEN_2075;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_rs2_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_rs2_paddr <= _GEN_2067;
      end
    end else begin
      buf_1_rs2_paddr <= _GEN_2067;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_rd_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_rd_paddr <= _GEN_2059;
      end
    end else begin
      buf_1_rd_paddr <= _GEN_2059;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_1_rob_addr <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h1 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_1_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 198:48]
      end else begin
        buf_1_rob_addr <= _GEN_2043;
      end
    end else begin
      buf_1_rob_addr <= _GEN_2043;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_valid <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_valid <= _GEN_2236;
      end
    end else begin
      buf_2_valid <= _GEN_2236;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_pc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_pc <= _GEN_2228;
      end
    end else begin
      buf_2_pc <= _GEN_2228;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_npc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_npc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_npc <= io_in_bits_vec_1_npc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_npc <= _GEN_2220;
      end
    end else begin
      buf_2_npc <= _GEN_2220;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_inst <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_inst <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_inst <= io_in_bits_vec_1_inst; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_inst <= _GEN_2212;
      end
    end else begin
      buf_2_inst <= _GEN_2212;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_fu_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_fu_code <= _GEN_2204;
      end
    end else begin
      buf_2_fu_code <= _GEN_2204;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_alu_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_alu_code <= _GEN_2196;
      end
    end else begin
      buf_2_alu_code <= _GEN_2196;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_jmp_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_jmp_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_jmp_code <= io_in_bits_vec_1_jmp_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_jmp_code <= _GEN_2188;
      end
    end else begin
      buf_2_jmp_code <= _GEN_2188;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_sys_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_sys_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_sys_code <= io_in_bits_vec_1_sys_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_sys_code <= _GEN_2164;
      end
    end else begin
      buf_2_sys_code <= _GEN_2164;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_w_type <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_w_type <= _GEN_2156;
      end
    end else begin
      buf_2_w_type <= _GEN_2156;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_rs1_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_rs1_src <= _GEN_2148;
      end
    end else begin
      buf_2_rs1_src <= _GEN_2148;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_rs2_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_rs2_src <= _GEN_2140;
      end
    end else begin
      buf_2_rs2_src <= _GEN_2140;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_rd_en <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_rd_en <= _GEN_2108;
      end
    end else begin
      buf_2_rd_en <= _GEN_2108;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_imm <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_imm <= _GEN_2100;
      end
    end else begin
      buf_2_imm <= _GEN_2100;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_pred_br <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_pred_br <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_pred_br <= io_in_bits_vec_1_pred_br; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_pred_br <= _GEN_2092;
      end
    end else begin
      buf_2_pred_br <= _GEN_2092;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_pred_bpc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_pred_bpc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_pred_bpc <= io_in_bits_vec_1_pred_bpc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_pred_bpc <= _GEN_2084;
      end
    end else begin
      buf_2_pred_bpc <= _GEN_2084;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_rs1_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_rs1_paddr <= _GEN_2076;
      end
    end else begin
      buf_2_rs1_paddr <= _GEN_2076;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_rs2_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_rs2_paddr <= _GEN_2068;
      end
    end else begin
      buf_2_rs2_paddr <= _GEN_2068;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_rd_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_rd_paddr <= _GEN_2060;
      end
    end else begin
      buf_2_rd_paddr <= _GEN_2060;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_2_rob_addr <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h2 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_2_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 198:48]
      end else begin
        buf_2_rob_addr <= _GEN_2044;
      end
    end else begin
      buf_2_rob_addr <= _GEN_2044;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_valid <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_valid <= _GEN_2237;
      end
    end else begin
      buf_3_valid <= _GEN_2237;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_pc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_pc <= _GEN_2229;
      end
    end else begin
      buf_3_pc <= _GEN_2229;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_npc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_npc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_npc <= io_in_bits_vec_1_npc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_npc <= _GEN_2221;
      end
    end else begin
      buf_3_npc <= _GEN_2221;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_inst <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_inst <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_inst <= io_in_bits_vec_1_inst; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_inst <= _GEN_2213;
      end
    end else begin
      buf_3_inst <= _GEN_2213;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_fu_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_fu_code <= _GEN_2205;
      end
    end else begin
      buf_3_fu_code <= _GEN_2205;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_alu_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_alu_code <= _GEN_2197;
      end
    end else begin
      buf_3_alu_code <= _GEN_2197;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_jmp_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_jmp_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_jmp_code <= io_in_bits_vec_1_jmp_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_jmp_code <= _GEN_2189;
      end
    end else begin
      buf_3_jmp_code <= _GEN_2189;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_sys_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_sys_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_sys_code <= io_in_bits_vec_1_sys_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_sys_code <= _GEN_2165;
      end
    end else begin
      buf_3_sys_code <= _GEN_2165;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_w_type <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_w_type <= _GEN_2157;
      end
    end else begin
      buf_3_w_type <= _GEN_2157;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_rs1_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_rs1_src <= _GEN_2149;
      end
    end else begin
      buf_3_rs1_src <= _GEN_2149;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_rs2_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_rs2_src <= _GEN_2141;
      end
    end else begin
      buf_3_rs2_src <= _GEN_2141;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_rd_en <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_rd_en <= _GEN_2109;
      end
    end else begin
      buf_3_rd_en <= _GEN_2109;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_imm <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_imm <= _GEN_2101;
      end
    end else begin
      buf_3_imm <= _GEN_2101;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_pred_br <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_pred_br <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_pred_br <= io_in_bits_vec_1_pred_br; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_pred_br <= _GEN_2093;
      end
    end else begin
      buf_3_pred_br <= _GEN_2093;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_pred_bpc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_pred_bpc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_pred_bpc <= io_in_bits_vec_1_pred_bpc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_pred_bpc <= _GEN_2085;
      end
    end else begin
      buf_3_pred_bpc <= _GEN_2085;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_rs1_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_rs1_paddr <= _GEN_2077;
      end
    end else begin
      buf_3_rs1_paddr <= _GEN_2077;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_rs2_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_rs2_paddr <= _GEN_2069;
      end
    end else begin
      buf_3_rs2_paddr <= _GEN_2069;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_rd_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_rd_paddr <= _GEN_2061;
      end
    end else begin
      buf_3_rd_paddr <= _GEN_2061;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_3_rob_addr <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h3 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_3_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 198:48]
      end else begin
        buf_3_rob_addr <= _GEN_2045;
      end
    end else begin
      buf_3_rob_addr <= _GEN_2045;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_valid <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_valid <= _GEN_2238;
      end
    end else begin
      buf_4_valid <= _GEN_2238;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_pc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_pc <= _GEN_2230;
      end
    end else begin
      buf_4_pc <= _GEN_2230;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_npc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_npc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_npc <= io_in_bits_vec_1_npc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_npc <= _GEN_2222;
      end
    end else begin
      buf_4_npc <= _GEN_2222;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_inst <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_inst <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_inst <= io_in_bits_vec_1_inst; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_inst <= _GEN_2214;
      end
    end else begin
      buf_4_inst <= _GEN_2214;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_fu_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_fu_code <= _GEN_2206;
      end
    end else begin
      buf_4_fu_code <= _GEN_2206;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_alu_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_alu_code <= _GEN_2198;
      end
    end else begin
      buf_4_alu_code <= _GEN_2198;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_jmp_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_jmp_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_jmp_code <= io_in_bits_vec_1_jmp_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_jmp_code <= _GEN_2190;
      end
    end else begin
      buf_4_jmp_code <= _GEN_2190;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_sys_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_sys_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_sys_code <= io_in_bits_vec_1_sys_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_sys_code <= _GEN_2166;
      end
    end else begin
      buf_4_sys_code <= _GEN_2166;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_w_type <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_w_type <= _GEN_2158;
      end
    end else begin
      buf_4_w_type <= _GEN_2158;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_rs1_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_rs1_src <= _GEN_2150;
      end
    end else begin
      buf_4_rs1_src <= _GEN_2150;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_rs2_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_rs2_src <= _GEN_2142;
      end
    end else begin
      buf_4_rs2_src <= _GEN_2142;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_rd_en <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_rd_en <= _GEN_2110;
      end
    end else begin
      buf_4_rd_en <= _GEN_2110;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_imm <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_imm <= _GEN_2102;
      end
    end else begin
      buf_4_imm <= _GEN_2102;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_pred_br <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_pred_br <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_pred_br <= io_in_bits_vec_1_pred_br; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_pred_br <= _GEN_2094;
      end
    end else begin
      buf_4_pred_br <= _GEN_2094;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_pred_bpc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_pred_bpc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_pred_bpc <= io_in_bits_vec_1_pred_bpc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_pred_bpc <= _GEN_2086;
      end
    end else begin
      buf_4_pred_bpc <= _GEN_2086;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_rs1_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_rs1_paddr <= _GEN_2078;
      end
    end else begin
      buf_4_rs1_paddr <= _GEN_2078;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_rs2_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_rs2_paddr <= _GEN_2070;
      end
    end else begin
      buf_4_rs2_paddr <= _GEN_2070;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_rd_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_rd_paddr <= _GEN_2062;
      end
    end else begin
      buf_4_rd_paddr <= _GEN_2062;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_4_rob_addr <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h4 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_4_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 198:48]
      end else begin
        buf_4_rob_addr <= _GEN_2046;
      end
    end else begin
      buf_4_rob_addr <= _GEN_2046;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_valid <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_valid <= _GEN_2239;
      end
    end else begin
      buf_5_valid <= _GEN_2239;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_pc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_pc <= _GEN_2231;
      end
    end else begin
      buf_5_pc <= _GEN_2231;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_npc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_npc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_npc <= io_in_bits_vec_1_npc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_npc <= _GEN_2223;
      end
    end else begin
      buf_5_npc <= _GEN_2223;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_inst <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_inst <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_inst <= io_in_bits_vec_1_inst; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_inst <= _GEN_2215;
      end
    end else begin
      buf_5_inst <= _GEN_2215;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_fu_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_fu_code <= _GEN_2207;
      end
    end else begin
      buf_5_fu_code <= _GEN_2207;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_alu_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_alu_code <= _GEN_2199;
      end
    end else begin
      buf_5_alu_code <= _GEN_2199;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_jmp_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_jmp_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_jmp_code <= io_in_bits_vec_1_jmp_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_jmp_code <= _GEN_2191;
      end
    end else begin
      buf_5_jmp_code <= _GEN_2191;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_sys_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_sys_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_sys_code <= io_in_bits_vec_1_sys_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_sys_code <= _GEN_2167;
      end
    end else begin
      buf_5_sys_code <= _GEN_2167;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_w_type <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_w_type <= _GEN_2159;
      end
    end else begin
      buf_5_w_type <= _GEN_2159;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_rs1_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_rs1_src <= _GEN_2151;
      end
    end else begin
      buf_5_rs1_src <= _GEN_2151;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_rs2_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_rs2_src <= _GEN_2143;
      end
    end else begin
      buf_5_rs2_src <= _GEN_2143;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_rd_en <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_rd_en <= _GEN_2111;
      end
    end else begin
      buf_5_rd_en <= _GEN_2111;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_imm <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_imm <= _GEN_2103;
      end
    end else begin
      buf_5_imm <= _GEN_2103;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_pred_br <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_pred_br <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_pred_br <= io_in_bits_vec_1_pred_br; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_pred_br <= _GEN_2095;
      end
    end else begin
      buf_5_pred_br <= _GEN_2095;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_pred_bpc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_pred_bpc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_pred_bpc <= io_in_bits_vec_1_pred_bpc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_pred_bpc <= _GEN_2087;
      end
    end else begin
      buf_5_pred_bpc <= _GEN_2087;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_rs1_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_rs1_paddr <= _GEN_2079;
      end
    end else begin
      buf_5_rs1_paddr <= _GEN_2079;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_rs2_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_rs2_paddr <= _GEN_2071;
      end
    end else begin
      buf_5_rs2_paddr <= _GEN_2071;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_rd_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_rd_paddr <= _GEN_2063;
      end
    end else begin
      buf_5_rd_paddr <= _GEN_2063;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_5_rob_addr <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h5 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_5_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 198:48]
      end else begin
        buf_5_rob_addr <= _GEN_2047;
      end
    end else begin
      buf_5_rob_addr <= _GEN_2047;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_valid <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_valid <= _GEN_2240;
      end
    end else begin
      buf_6_valid <= _GEN_2240;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_pc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_pc <= _GEN_2232;
      end
    end else begin
      buf_6_pc <= _GEN_2232;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_npc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_npc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_npc <= io_in_bits_vec_1_npc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_npc <= _GEN_2224;
      end
    end else begin
      buf_6_npc <= _GEN_2224;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_inst <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_inst <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_inst <= io_in_bits_vec_1_inst; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_inst <= _GEN_2216;
      end
    end else begin
      buf_6_inst <= _GEN_2216;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_fu_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_fu_code <= _GEN_2208;
      end
    end else begin
      buf_6_fu_code <= _GEN_2208;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_alu_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_alu_code <= _GEN_2200;
      end
    end else begin
      buf_6_alu_code <= _GEN_2200;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_jmp_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_jmp_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_jmp_code <= io_in_bits_vec_1_jmp_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_jmp_code <= _GEN_2192;
      end
    end else begin
      buf_6_jmp_code <= _GEN_2192;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_sys_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_sys_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_sys_code <= io_in_bits_vec_1_sys_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_sys_code <= _GEN_2168;
      end
    end else begin
      buf_6_sys_code <= _GEN_2168;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_w_type <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_w_type <= _GEN_2160;
      end
    end else begin
      buf_6_w_type <= _GEN_2160;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_rs1_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_rs1_src <= _GEN_2152;
      end
    end else begin
      buf_6_rs1_src <= _GEN_2152;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_rs2_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_rs2_src <= _GEN_2144;
      end
    end else begin
      buf_6_rs2_src <= _GEN_2144;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_rd_en <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_rd_en <= _GEN_2112;
      end
    end else begin
      buf_6_rd_en <= _GEN_2112;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_imm <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_imm <= _GEN_2104;
      end
    end else begin
      buf_6_imm <= _GEN_2104;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_pred_br <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_pred_br <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_pred_br <= io_in_bits_vec_1_pred_br; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_pred_br <= _GEN_2096;
      end
    end else begin
      buf_6_pred_br <= _GEN_2096;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_pred_bpc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_pred_bpc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_pred_bpc <= io_in_bits_vec_1_pred_bpc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_pred_bpc <= _GEN_2088;
      end
    end else begin
      buf_6_pred_bpc <= _GEN_2088;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_rs1_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_rs1_paddr <= _GEN_2080;
      end
    end else begin
      buf_6_rs1_paddr <= _GEN_2080;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_rs2_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_rs2_paddr <= _GEN_2072;
      end
    end else begin
      buf_6_rs2_paddr <= _GEN_2072;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_rd_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_rd_paddr <= _GEN_2064;
      end
    end else begin
      buf_6_rd_paddr <= _GEN_2064;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_6_rob_addr <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h6 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_6_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 198:48]
      end else begin
        buf_6_rob_addr <= _GEN_2048;
      end
    end else begin
      buf_6_rob_addr <= _GEN_2048;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_valid <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_valid <= _GEN_2241;
      end
    end else begin
      buf_7_valid <= _GEN_2241;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_pc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_pc <= _GEN_2233;
      end
    end else begin
      buf_7_pc <= _GEN_2233;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_npc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_npc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_npc <= io_in_bits_vec_1_npc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_npc <= _GEN_2225;
      end
    end else begin
      buf_7_npc <= _GEN_2225;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_inst <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_inst <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_inst <= io_in_bits_vec_1_inst; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_inst <= _GEN_2217;
      end
    end else begin
      buf_7_inst <= _GEN_2217;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_fu_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_fu_code <= _GEN_2209;
      end
    end else begin
      buf_7_fu_code <= _GEN_2209;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_alu_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_alu_code <= _GEN_2201;
      end
    end else begin
      buf_7_alu_code <= _GEN_2201;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_jmp_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_jmp_code <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_jmp_code <= io_in_bits_vec_1_jmp_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_jmp_code <= _GEN_2193;
      end
    end else begin
      buf_7_jmp_code <= _GEN_2193;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_sys_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_sys_code <= 3'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_sys_code <= io_in_bits_vec_1_sys_code; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_sys_code <= _GEN_2169;
      end
    end else begin
      buf_7_sys_code <= _GEN_2169;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_w_type <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_w_type <= _GEN_2161;
      end
    end else begin
      buf_7_w_type <= _GEN_2161;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_rs1_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_rs1_src <= _GEN_2153;
      end
    end else begin
      buf_7_rs1_src <= _GEN_2153;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_rs2_src <= 2'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_rs2_src <= _GEN_2145;
      end
    end else begin
      buf_7_rs2_src <= _GEN_2145;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_rd_en <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_rd_en <= _GEN_2113;
      end
    end else begin
      buf_7_rd_en <= _GEN_2113;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_imm <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_imm <= _GEN_2105;
      end
    end else begin
      buf_7_imm <= _GEN_2105;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_pred_br <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_pred_br <= 1'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_pred_br <= io_in_bits_vec_1_pred_br; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_pred_br <= _GEN_2097;
      end
    end else begin
      buf_7_pred_br <= _GEN_2097;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_pred_bpc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_pred_bpc <= 32'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_pred_bpc <= io_in_bits_vec_1_pred_bpc; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_pred_bpc <= _GEN_2089;
      end
    end else begin
      buf_7_pred_bpc <= _GEN_2089;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_rs1_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_rs1_paddr <= _GEN_2081;
      end
    end else begin
      buf_7_rs1_paddr <= _GEN_2081;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_rs2_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_rs2_paddr <= _GEN_2073;
      end
    end else begin
      buf_7_rs2_paddr <= _GEN_2073;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_rd_paddr <= 6'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_rd_paddr <= _GEN_2065;
      end
    end else begin
      buf_7_rd_paddr <= _GEN_2065;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      buf_7_rob_addr <= 4'h0; // @[IssueUnit.scala 214:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 197:51]
      if (3'h7 == _GEN_2243[2:0]) begin // @[IssueUnit.scala 198:48]
        buf_7_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 198:48]
      end else begin
        buf_7_rob_addr <= _GEN_2049;
      end
    end else begin
      buf_7_rob_addr <= _GEN_2049;
    end
    if (reset) begin // @[IssueUnit.scala 102:24]
      enq_vec_0 <= 4'h0; // @[IssueUnit.scala 102:24]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      enq_vec_0 <= 4'h0; // @[IssueUnit.scala 216:13]
    end else if ((_T | (|_T_172)) & _T_155) begin // @[IssueUnit.scala 204:70]
      enq_vec_0 <= next_enq_vec_0; // @[IssueUnit.scala 205:13]
    end
    if (reset) begin // @[IssueUnit.scala 102:24]
      enq_vec_1 <= 4'h1; // @[IssueUnit.scala 102:24]
    end else if (io_flush) begin // @[IssueUnit.scala 212:19]
      enq_vec_1 <= 4'h1; // @[IssueUnit.scala 216:13]
    end else if ((_T | (|_T_172)) & _T_155) begin // @[IssueUnit.scala 204:70]
      enq_vec_1 <= next_enq_vec_1; // @[IssueUnit.scala 205:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  buf_0_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  buf_0_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  buf_0_npc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  buf_0_inst = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  buf_0_fu_code = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  buf_0_alu_code = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  buf_0_jmp_code = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  buf_0_sys_code = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  buf_0_w_type = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  buf_0_rs1_src = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  buf_0_rs2_src = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  buf_0_rd_en = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  buf_0_imm = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  buf_0_pred_br = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  buf_0_pred_bpc = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  buf_0_rs1_paddr = _RAND_15[5:0];
  _RAND_16 = {1{`RANDOM}};
  buf_0_rs2_paddr = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  buf_0_rd_paddr = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  buf_0_rob_addr = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  buf_1_valid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  buf_1_pc = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  buf_1_npc = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  buf_1_inst = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  buf_1_fu_code = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  buf_1_alu_code = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  buf_1_jmp_code = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  buf_1_sys_code = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  buf_1_w_type = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  buf_1_rs1_src = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  buf_1_rs2_src = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  buf_1_rd_en = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  buf_1_imm = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  buf_1_pred_br = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  buf_1_pred_bpc = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  buf_1_rs1_paddr = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  buf_1_rs2_paddr = _RAND_35[5:0];
  _RAND_36 = {1{`RANDOM}};
  buf_1_rd_paddr = _RAND_36[5:0];
  _RAND_37 = {1{`RANDOM}};
  buf_1_rob_addr = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  buf_2_valid = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  buf_2_pc = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  buf_2_npc = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  buf_2_inst = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  buf_2_fu_code = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  buf_2_alu_code = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  buf_2_jmp_code = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  buf_2_sys_code = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  buf_2_w_type = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  buf_2_rs1_src = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  buf_2_rs2_src = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  buf_2_rd_en = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  buf_2_imm = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  buf_2_pred_br = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  buf_2_pred_bpc = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  buf_2_rs1_paddr = _RAND_53[5:0];
  _RAND_54 = {1{`RANDOM}};
  buf_2_rs2_paddr = _RAND_54[5:0];
  _RAND_55 = {1{`RANDOM}};
  buf_2_rd_paddr = _RAND_55[5:0];
  _RAND_56 = {1{`RANDOM}};
  buf_2_rob_addr = _RAND_56[3:0];
  _RAND_57 = {1{`RANDOM}};
  buf_3_valid = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  buf_3_pc = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  buf_3_npc = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  buf_3_inst = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  buf_3_fu_code = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  buf_3_alu_code = _RAND_62[3:0];
  _RAND_63 = {1{`RANDOM}};
  buf_3_jmp_code = _RAND_63[3:0];
  _RAND_64 = {1{`RANDOM}};
  buf_3_sys_code = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  buf_3_w_type = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  buf_3_rs1_src = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  buf_3_rs2_src = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  buf_3_rd_en = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  buf_3_imm = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  buf_3_pred_br = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  buf_3_pred_bpc = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  buf_3_rs1_paddr = _RAND_72[5:0];
  _RAND_73 = {1{`RANDOM}};
  buf_3_rs2_paddr = _RAND_73[5:0];
  _RAND_74 = {1{`RANDOM}};
  buf_3_rd_paddr = _RAND_74[5:0];
  _RAND_75 = {1{`RANDOM}};
  buf_3_rob_addr = _RAND_75[3:0];
  _RAND_76 = {1{`RANDOM}};
  buf_4_valid = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  buf_4_pc = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  buf_4_npc = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  buf_4_inst = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  buf_4_fu_code = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  buf_4_alu_code = _RAND_81[3:0];
  _RAND_82 = {1{`RANDOM}};
  buf_4_jmp_code = _RAND_82[3:0];
  _RAND_83 = {1{`RANDOM}};
  buf_4_sys_code = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  buf_4_w_type = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  buf_4_rs1_src = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  buf_4_rs2_src = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  buf_4_rd_en = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  buf_4_imm = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  buf_4_pred_br = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  buf_4_pred_bpc = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  buf_4_rs1_paddr = _RAND_91[5:0];
  _RAND_92 = {1{`RANDOM}};
  buf_4_rs2_paddr = _RAND_92[5:0];
  _RAND_93 = {1{`RANDOM}};
  buf_4_rd_paddr = _RAND_93[5:0];
  _RAND_94 = {1{`RANDOM}};
  buf_4_rob_addr = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  buf_5_valid = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  buf_5_pc = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  buf_5_npc = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  buf_5_inst = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  buf_5_fu_code = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  buf_5_alu_code = _RAND_100[3:0];
  _RAND_101 = {1{`RANDOM}};
  buf_5_jmp_code = _RAND_101[3:0];
  _RAND_102 = {1{`RANDOM}};
  buf_5_sys_code = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  buf_5_w_type = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  buf_5_rs1_src = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  buf_5_rs2_src = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  buf_5_rd_en = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  buf_5_imm = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  buf_5_pred_br = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  buf_5_pred_bpc = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  buf_5_rs1_paddr = _RAND_110[5:0];
  _RAND_111 = {1{`RANDOM}};
  buf_5_rs2_paddr = _RAND_111[5:0];
  _RAND_112 = {1{`RANDOM}};
  buf_5_rd_paddr = _RAND_112[5:0];
  _RAND_113 = {1{`RANDOM}};
  buf_5_rob_addr = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  buf_6_valid = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  buf_6_pc = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  buf_6_npc = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  buf_6_inst = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  buf_6_fu_code = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  buf_6_alu_code = _RAND_119[3:0];
  _RAND_120 = {1{`RANDOM}};
  buf_6_jmp_code = _RAND_120[3:0];
  _RAND_121 = {1{`RANDOM}};
  buf_6_sys_code = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  buf_6_w_type = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  buf_6_rs1_src = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  buf_6_rs2_src = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  buf_6_rd_en = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  buf_6_imm = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  buf_6_pred_br = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  buf_6_pred_bpc = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  buf_6_rs1_paddr = _RAND_129[5:0];
  _RAND_130 = {1{`RANDOM}};
  buf_6_rs2_paddr = _RAND_130[5:0];
  _RAND_131 = {1{`RANDOM}};
  buf_6_rd_paddr = _RAND_131[5:0];
  _RAND_132 = {1{`RANDOM}};
  buf_6_rob_addr = _RAND_132[3:0];
  _RAND_133 = {1{`RANDOM}};
  buf_7_valid = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  buf_7_pc = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  buf_7_npc = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  buf_7_inst = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  buf_7_fu_code = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  buf_7_alu_code = _RAND_138[3:0];
  _RAND_139 = {1{`RANDOM}};
  buf_7_jmp_code = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  buf_7_sys_code = _RAND_140[2:0];
  _RAND_141 = {1{`RANDOM}};
  buf_7_w_type = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  buf_7_rs1_src = _RAND_142[1:0];
  _RAND_143 = {1{`RANDOM}};
  buf_7_rs2_src = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  buf_7_rd_en = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  buf_7_imm = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  buf_7_pred_br = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  buf_7_pred_bpc = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  buf_7_rs1_paddr = _RAND_148[5:0];
  _RAND_149 = {1{`RANDOM}};
  buf_7_rs2_paddr = _RAND_149[5:0];
  _RAND_150 = {1{`RANDOM}};
  buf_7_rd_paddr = _RAND_150[5:0];
  _RAND_151 = {1{`RANDOM}};
  buf_7_rob_addr = _RAND_151[3:0];
  _RAND_152 = {1{`RANDOM}};
  enq_vec_0 = _RAND_152[3:0];
  _RAND_153 = {1{`RANDOM}};
  enq_vec_1 = _RAND_153[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_MemIssueQueueOutOfOrder(
  input         clock,
  input         reset,
  input         io_flush,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_vec_0_valid,
  input  [31:0] io_in_bits_vec_0_pc,
  input  [2:0]  io_in_bits_vec_0_fu_code,
  input  [3:0]  io_in_bits_vec_0_alu_code,
  input  [1:0]  io_in_bits_vec_0_mem_code,
  input  [1:0]  io_in_bits_vec_0_mem_size,
  input         io_in_bits_vec_0_w_type,
  input  [1:0]  io_in_bits_vec_0_rs1_src,
  input  [1:0]  io_in_bits_vec_0_rs2_src,
  input         io_in_bits_vec_0_rd_en,
  input  [31:0] io_in_bits_vec_0_imm,
  input  [5:0]  io_in_bits_vec_0_rs1_paddr,
  input  [5:0]  io_in_bits_vec_0_rs2_paddr,
  input  [5:0]  io_in_bits_vec_0_rd_paddr,
  input         io_in_bits_vec_1_valid,
  input  [31:0] io_in_bits_vec_1_pc,
  input  [2:0]  io_in_bits_vec_1_fu_code,
  input  [3:0]  io_in_bits_vec_1_alu_code,
  input  [1:0]  io_in_bits_vec_1_mem_code,
  input  [1:0]  io_in_bits_vec_1_mem_size,
  input         io_in_bits_vec_1_w_type,
  input  [1:0]  io_in_bits_vec_1_rs1_src,
  input  [1:0]  io_in_bits_vec_1_rs2_src,
  input         io_in_bits_vec_1_rd_en,
  input  [31:0] io_in_bits_vec_1_imm,
  input  [5:0]  io_in_bits_vec_1_rs1_paddr,
  input  [5:0]  io_in_bits_vec_1_rs2_paddr,
  input  [5:0]  io_in_bits_vec_1_rd_paddr,
  input  [3:0]  io_rob_addr_0,
  input  [3:0]  io_rob_addr_1,
  output        io_out_0_valid,
  output [31:0] io_out_0_pc,
  output [2:0]  io_out_0_fu_code,
  output [3:0]  io_out_0_alu_code,
  output [1:0]  io_out_0_mem_code,
  output [1:0]  io_out_0_mem_size,
  output        io_out_0_w_type,
  output [1:0]  io_out_0_rs1_src,
  output [1:0]  io_out_0_rs2_src,
  output        io_out_0_rd_en,
  output [31:0] io_out_0_imm,
  output [5:0]  io_out_0_rs1_paddr,
  output [5:0]  io_out_0_rs2_paddr,
  output [5:0]  io_out_0_rd_paddr,
  output [3:0]  io_out_0_rob_addr,
  input         io_avail_list_0,
  input         io_avail_list_1,
  input         io_avail_list_2,
  input         io_avail_list_3,
  input         io_avail_list_4,
  input         io_avail_list_5,
  input         io_avail_list_6,
  input         io_avail_list_7,
  input         io_avail_list_8,
  input         io_avail_list_9,
  input         io_avail_list_10,
  input         io_avail_list_11,
  input         io_avail_list_12,
  input         io_avail_list_13,
  input         io_avail_list_14,
  input         io_avail_list_15,
  input         io_avail_list_16,
  input         io_avail_list_17,
  input         io_avail_list_18,
  input         io_avail_list_19,
  input         io_avail_list_20,
  input         io_avail_list_21,
  input         io_avail_list_22,
  input         io_avail_list_23,
  input         io_avail_list_24,
  input         io_avail_list_25,
  input         io_avail_list_26,
  input         io_avail_list_27,
  input         io_avail_list_28,
  input         io_avail_list_29,
  input         io_avail_list_30,
  input         io_avail_list_31,
  input         io_avail_list_32,
  input         io_avail_list_33,
  input         io_avail_list_34,
  input         io_avail_list_35,
  input         io_avail_list_36,
  input         io_avail_list_37,
  input         io_avail_list_38,
  input         io_avail_list_39,
  input         io_avail_list_40,
  input         io_avail_list_41,
  input         io_avail_list_42,
  input         io_avail_list_43,
  input         io_avail_list_44,
  input         io_avail_list_45,
  input         io_avail_list_46,
  input         io_avail_list_47,
  input         io_avail_list_48,
  input         io_avail_list_49,
  input         io_avail_list_50,
  input         io_avail_list_51,
  input         io_avail_list_52,
  input         io_avail_list_53,
  input         io_avail_list_54,
  input         io_avail_list_55,
  input         io_avail_list_56,
  input         io_avail_list_57,
  input         io_avail_list_58,
  input         io_avail_list_59,
  input         io_avail_list_60,
  input         io_avail_list_61,
  input         io_avail_list_62,
  input         io_avail_list_63,
  input         io_fu_ready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
`endif // RANDOMIZE_REG_INIT
  reg  buf_0_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_0_pc; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_0_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_0_alu_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_0_mem_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_0_mem_size; // @[IssueUnit.scala 97:20]
  reg  buf_0_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_0_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_0_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_0_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_0_imm; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_0_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_0_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_0_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_0_rob_addr; // @[IssueUnit.scala 97:20]
  reg  buf_1_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_1_pc; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_1_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_1_alu_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_1_mem_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_1_mem_size; // @[IssueUnit.scala 97:20]
  reg  buf_1_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_1_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_1_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_1_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_1_imm; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_1_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_1_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_1_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_1_rob_addr; // @[IssueUnit.scala 97:20]
  reg  buf_2_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_2_pc; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_2_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_2_alu_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_2_mem_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_2_mem_size; // @[IssueUnit.scala 97:20]
  reg  buf_2_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_2_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_2_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_2_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_2_imm; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_2_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_2_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_2_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_2_rob_addr; // @[IssueUnit.scala 97:20]
  reg  buf_3_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_3_pc; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_3_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_3_alu_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_3_mem_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_3_mem_size; // @[IssueUnit.scala 97:20]
  reg  buf_3_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_3_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_3_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_3_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_3_imm; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_3_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_3_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_3_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_3_rob_addr; // @[IssueUnit.scala 97:20]
  reg  buf_4_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_4_pc; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_4_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_4_alu_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_4_mem_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_4_mem_size; // @[IssueUnit.scala 97:20]
  reg  buf_4_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_4_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_4_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_4_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_4_imm; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_4_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_4_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_4_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_4_rob_addr; // @[IssueUnit.scala 97:20]
  reg  buf_5_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_5_pc; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_5_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_5_alu_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_5_mem_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_5_mem_size; // @[IssueUnit.scala 97:20]
  reg  buf_5_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_5_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_5_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_5_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_5_imm; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_5_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_5_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_5_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_5_rob_addr; // @[IssueUnit.scala 97:20]
  reg  buf_6_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_6_pc; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_6_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_6_alu_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_6_mem_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_6_mem_size; // @[IssueUnit.scala 97:20]
  reg  buf_6_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_6_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_6_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_6_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_6_imm; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_6_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_6_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_6_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_6_rob_addr; // @[IssueUnit.scala 97:20]
  reg  buf_7_valid; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_7_pc; // @[IssueUnit.scala 97:20]
  reg [2:0] buf_7_fu_code; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_7_alu_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_7_mem_code; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_7_mem_size; // @[IssueUnit.scala 97:20]
  reg  buf_7_w_type; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_7_rs1_src; // @[IssueUnit.scala 97:20]
  reg [1:0] buf_7_rs2_src; // @[IssueUnit.scala 97:20]
  reg  buf_7_rd_en; // @[IssueUnit.scala 97:20]
  reg [31:0] buf_7_imm; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_7_rs1_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_7_rs2_paddr; // @[IssueUnit.scala 97:20]
  reg [5:0] buf_7_rd_paddr; // @[IssueUnit.scala 97:20]
  reg [3:0] buf_7_rob_addr; // @[IssueUnit.scala 97:20]
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_1 = io_in_bits_vec_0_valid + io_in_bits_vec_1_valid; // @[Bitwise.scala 47:55]
  wire [1:0] num_enq = _T ? _T_1 : 2'h0; // @[IssueUnit.scala 99:20]
  reg [3:0] enq_vec_0; // @[IssueUnit.scala 102:24]
  reg [3:0] enq_vec_1; // @[IssueUnit.scala 102:24]
  wire [3:0] _GEN_2440 = {{3'd0}, io_out_0_valid}; // @[IssueUnit.scala 103:44]
  wire [3:0] enq_vec_real_0 = enq_vec_0 - _GEN_2440; // @[IssueUnit.scala 103:44]
  wire [3:0] enq_vec_real_1 = enq_vec_1 - _GEN_2440; // @[IssueUnit.scala 103:44]
  wire  is_store_0 = buf_0_mem_code == 2'h3; // @[IssueUnit.scala 243:37]
  wire  is_store_1 = buf_1_mem_code == 2'h3; // @[IssueUnit.scala 243:37]
  wire  is_store_2 = buf_2_mem_code == 2'h3; // @[IssueUnit.scala 243:37]
  wire  is_store_3 = buf_3_mem_code == 2'h3; // @[IssueUnit.scala 243:37]
  wire  is_store_4 = buf_4_mem_code == 2'h3; // @[IssueUnit.scala 243:37]
  wire  is_store_5 = buf_5_mem_code == 2'h3; // @[IssueUnit.scala 243:37]
  wire  is_store_6 = buf_6_mem_code == 2'h3; // @[IssueUnit.scala 243:37]
  wire  is_store_7 = buf_7_mem_code == 2'h3; // @[IssueUnit.scala 243:37]
  wire [1:0] _T_17 = {is_store_0,is_store_1}; // @[Cat.scala 30:58]
  wire  store_mask_1 = ~(|_T_17); // @[IssueUnit.scala 248:22]
  wire [2:0] _T_20 = {is_store_0,is_store_1,is_store_2}; // @[Cat.scala 30:58]
  wire  store_mask_2 = ~(|_T_20); // @[IssueUnit.scala 248:22]
  wire [3:0] _T_23 = {is_store_0,is_store_1,is_store_2,is_store_3}; // @[Cat.scala 30:58]
  wire  store_mask_3 = ~(|_T_23); // @[IssueUnit.scala 248:22]
  wire [4:0] _T_26 = {is_store_0,is_store_1,is_store_2,is_store_3,is_store_4}; // @[Cat.scala 30:58]
  wire  store_mask_4 = ~(|_T_26); // @[IssueUnit.scala 248:22]
  wire [5:0] _T_29 = {is_store_0,is_store_1,is_store_2,is_store_3,is_store_4,is_store_5}; // @[Cat.scala 30:58]
  wire  store_mask_5 = ~(|_T_29); // @[IssueUnit.scala 248:22]
  wire [6:0] _T_32 = {is_store_0,is_store_1,is_store_2,is_store_3,is_store_4,is_store_5,is_store_6}; // @[Cat.scala 30:58]
  wire  store_mask_6 = ~(|_T_32); // @[IssueUnit.scala 248:22]
  wire [7:0] _T_35 = {is_store_0,is_store_1,is_store_2,is_store_3,is_store_4,is_store_5,is_store_6,is_store_7}; // @[Cat.scala 30:58]
  wire  store_mask_7 = ~(|_T_35); // @[IssueUnit.scala 248:22]
  wire  _GEN_1 = 6'h1 == buf_0_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_2 = 6'h2 == buf_0_rs1_paddr ? io_avail_list_2 : _GEN_1; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_3 = 6'h3 == buf_0_rs1_paddr ? io_avail_list_3 : _GEN_2; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_4 = 6'h4 == buf_0_rs1_paddr ? io_avail_list_4 : _GEN_3; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_5 = 6'h5 == buf_0_rs1_paddr ? io_avail_list_5 : _GEN_4; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_6 = 6'h6 == buf_0_rs1_paddr ? io_avail_list_6 : _GEN_5; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_7 = 6'h7 == buf_0_rs1_paddr ? io_avail_list_7 : _GEN_6; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_8 = 6'h8 == buf_0_rs1_paddr ? io_avail_list_8 : _GEN_7; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_9 = 6'h9 == buf_0_rs1_paddr ? io_avail_list_9 : _GEN_8; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_10 = 6'ha == buf_0_rs1_paddr ? io_avail_list_10 : _GEN_9; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_11 = 6'hb == buf_0_rs1_paddr ? io_avail_list_11 : _GEN_10; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_12 = 6'hc == buf_0_rs1_paddr ? io_avail_list_12 : _GEN_11; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_13 = 6'hd == buf_0_rs1_paddr ? io_avail_list_13 : _GEN_12; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_14 = 6'he == buf_0_rs1_paddr ? io_avail_list_14 : _GEN_13; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_15 = 6'hf == buf_0_rs1_paddr ? io_avail_list_15 : _GEN_14; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_16 = 6'h10 == buf_0_rs1_paddr ? io_avail_list_16 : _GEN_15; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_17 = 6'h11 == buf_0_rs1_paddr ? io_avail_list_17 : _GEN_16; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_18 = 6'h12 == buf_0_rs1_paddr ? io_avail_list_18 : _GEN_17; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_19 = 6'h13 == buf_0_rs1_paddr ? io_avail_list_19 : _GEN_18; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_20 = 6'h14 == buf_0_rs1_paddr ? io_avail_list_20 : _GEN_19; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_21 = 6'h15 == buf_0_rs1_paddr ? io_avail_list_21 : _GEN_20; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_22 = 6'h16 == buf_0_rs1_paddr ? io_avail_list_22 : _GEN_21; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_23 = 6'h17 == buf_0_rs1_paddr ? io_avail_list_23 : _GEN_22; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_24 = 6'h18 == buf_0_rs1_paddr ? io_avail_list_24 : _GEN_23; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_25 = 6'h19 == buf_0_rs1_paddr ? io_avail_list_25 : _GEN_24; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_26 = 6'h1a == buf_0_rs1_paddr ? io_avail_list_26 : _GEN_25; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_27 = 6'h1b == buf_0_rs1_paddr ? io_avail_list_27 : _GEN_26; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_28 = 6'h1c == buf_0_rs1_paddr ? io_avail_list_28 : _GEN_27; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_29 = 6'h1d == buf_0_rs1_paddr ? io_avail_list_29 : _GEN_28; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_30 = 6'h1e == buf_0_rs1_paddr ? io_avail_list_30 : _GEN_29; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_31 = 6'h1f == buf_0_rs1_paddr ? io_avail_list_31 : _GEN_30; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_32 = 6'h20 == buf_0_rs1_paddr ? io_avail_list_32 : _GEN_31; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_33 = 6'h21 == buf_0_rs1_paddr ? io_avail_list_33 : _GEN_32; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_34 = 6'h22 == buf_0_rs1_paddr ? io_avail_list_34 : _GEN_33; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_35 = 6'h23 == buf_0_rs1_paddr ? io_avail_list_35 : _GEN_34; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_36 = 6'h24 == buf_0_rs1_paddr ? io_avail_list_36 : _GEN_35; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_37 = 6'h25 == buf_0_rs1_paddr ? io_avail_list_37 : _GEN_36; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_38 = 6'h26 == buf_0_rs1_paddr ? io_avail_list_38 : _GEN_37; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_39 = 6'h27 == buf_0_rs1_paddr ? io_avail_list_39 : _GEN_38; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_40 = 6'h28 == buf_0_rs1_paddr ? io_avail_list_40 : _GEN_39; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_41 = 6'h29 == buf_0_rs1_paddr ? io_avail_list_41 : _GEN_40; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_42 = 6'h2a == buf_0_rs1_paddr ? io_avail_list_42 : _GEN_41; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_43 = 6'h2b == buf_0_rs1_paddr ? io_avail_list_43 : _GEN_42; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_44 = 6'h2c == buf_0_rs1_paddr ? io_avail_list_44 : _GEN_43; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_45 = 6'h2d == buf_0_rs1_paddr ? io_avail_list_45 : _GEN_44; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_46 = 6'h2e == buf_0_rs1_paddr ? io_avail_list_46 : _GEN_45; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_47 = 6'h2f == buf_0_rs1_paddr ? io_avail_list_47 : _GEN_46; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_48 = 6'h30 == buf_0_rs1_paddr ? io_avail_list_48 : _GEN_47; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_49 = 6'h31 == buf_0_rs1_paddr ? io_avail_list_49 : _GEN_48; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_50 = 6'h32 == buf_0_rs1_paddr ? io_avail_list_50 : _GEN_49; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_51 = 6'h33 == buf_0_rs1_paddr ? io_avail_list_51 : _GEN_50; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_52 = 6'h34 == buf_0_rs1_paddr ? io_avail_list_52 : _GEN_51; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_53 = 6'h35 == buf_0_rs1_paddr ? io_avail_list_53 : _GEN_52; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_54 = 6'h36 == buf_0_rs1_paddr ? io_avail_list_54 : _GEN_53; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_55 = 6'h37 == buf_0_rs1_paddr ? io_avail_list_55 : _GEN_54; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_56 = 6'h38 == buf_0_rs1_paddr ? io_avail_list_56 : _GEN_55; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_57 = 6'h39 == buf_0_rs1_paddr ? io_avail_list_57 : _GEN_56; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_58 = 6'h3a == buf_0_rs1_paddr ? io_avail_list_58 : _GEN_57; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_59 = 6'h3b == buf_0_rs1_paddr ? io_avail_list_59 : _GEN_58; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_60 = 6'h3c == buf_0_rs1_paddr ? io_avail_list_60 : _GEN_59; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_61 = 6'h3d == buf_0_rs1_paddr ? io_avail_list_61 : _GEN_60; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_62 = 6'h3e == buf_0_rs1_paddr ? io_avail_list_62 : _GEN_61; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_63 = 6'h3f == buf_0_rs1_paddr ? io_avail_list_63 : _GEN_62; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_65 = 6'h1 == buf_0_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_66 = 6'h2 == buf_0_rs2_paddr ? io_avail_list_2 : _GEN_65; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_67 = 6'h3 == buf_0_rs2_paddr ? io_avail_list_3 : _GEN_66; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_68 = 6'h4 == buf_0_rs2_paddr ? io_avail_list_4 : _GEN_67; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_69 = 6'h5 == buf_0_rs2_paddr ? io_avail_list_5 : _GEN_68; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_70 = 6'h6 == buf_0_rs2_paddr ? io_avail_list_6 : _GEN_69; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_71 = 6'h7 == buf_0_rs2_paddr ? io_avail_list_7 : _GEN_70; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_72 = 6'h8 == buf_0_rs2_paddr ? io_avail_list_8 : _GEN_71; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_73 = 6'h9 == buf_0_rs2_paddr ? io_avail_list_9 : _GEN_72; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_74 = 6'ha == buf_0_rs2_paddr ? io_avail_list_10 : _GEN_73; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_75 = 6'hb == buf_0_rs2_paddr ? io_avail_list_11 : _GEN_74; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_76 = 6'hc == buf_0_rs2_paddr ? io_avail_list_12 : _GEN_75; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_77 = 6'hd == buf_0_rs2_paddr ? io_avail_list_13 : _GEN_76; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_78 = 6'he == buf_0_rs2_paddr ? io_avail_list_14 : _GEN_77; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_79 = 6'hf == buf_0_rs2_paddr ? io_avail_list_15 : _GEN_78; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_80 = 6'h10 == buf_0_rs2_paddr ? io_avail_list_16 : _GEN_79; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_81 = 6'h11 == buf_0_rs2_paddr ? io_avail_list_17 : _GEN_80; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_82 = 6'h12 == buf_0_rs2_paddr ? io_avail_list_18 : _GEN_81; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_83 = 6'h13 == buf_0_rs2_paddr ? io_avail_list_19 : _GEN_82; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_84 = 6'h14 == buf_0_rs2_paddr ? io_avail_list_20 : _GEN_83; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_85 = 6'h15 == buf_0_rs2_paddr ? io_avail_list_21 : _GEN_84; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_86 = 6'h16 == buf_0_rs2_paddr ? io_avail_list_22 : _GEN_85; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_87 = 6'h17 == buf_0_rs2_paddr ? io_avail_list_23 : _GEN_86; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_88 = 6'h18 == buf_0_rs2_paddr ? io_avail_list_24 : _GEN_87; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_89 = 6'h19 == buf_0_rs2_paddr ? io_avail_list_25 : _GEN_88; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_90 = 6'h1a == buf_0_rs2_paddr ? io_avail_list_26 : _GEN_89; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_91 = 6'h1b == buf_0_rs2_paddr ? io_avail_list_27 : _GEN_90; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_92 = 6'h1c == buf_0_rs2_paddr ? io_avail_list_28 : _GEN_91; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_93 = 6'h1d == buf_0_rs2_paddr ? io_avail_list_29 : _GEN_92; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_94 = 6'h1e == buf_0_rs2_paddr ? io_avail_list_30 : _GEN_93; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_95 = 6'h1f == buf_0_rs2_paddr ? io_avail_list_31 : _GEN_94; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_96 = 6'h20 == buf_0_rs2_paddr ? io_avail_list_32 : _GEN_95; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_97 = 6'h21 == buf_0_rs2_paddr ? io_avail_list_33 : _GEN_96; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_98 = 6'h22 == buf_0_rs2_paddr ? io_avail_list_34 : _GEN_97; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_99 = 6'h23 == buf_0_rs2_paddr ? io_avail_list_35 : _GEN_98; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_100 = 6'h24 == buf_0_rs2_paddr ? io_avail_list_36 : _GEN_99; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_101 = 6'h25 == buf_0_rs2_paddr ? io_avail_list_37 : _GEN_100; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_102 = 6'h26 == buf_0_rs2_paddr ? io_avail_list_38 : _GEN_101; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_103 = 6'h27 == buf_0_rs2_paddr ? io_avail_list_39 : _GEN_102; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_104 = 6'h28 == buf_0_rs2_paddr ? io_avail_list_40 : _GEN_103; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_105 = 6'h29 == buf_0_rs2_paddr ? io_avail_list_41 : _GEN_104; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_106 = 6'h2a == buf_0_rs2_paddr ? io_avail_list_42 : _GEN_105; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_107 = 6'h2b == buf_0_rs2_paddr ? io_avail_list_43 : _GEN_106; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_108 = 6'h2c == buf_0_rs2_paddr ? io_avail_list_44 : _GEN_107; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_109 = 6'h2d == buf_0_rs2_paddr ? io_avail_list_45 : _GEN_108; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_110 = 6'h2e == buf_0_rs2_paddr ? io_avail_list_46 : _GEN_109; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_111 = 6'h2f == buf_0_rs2_paddr ? io_avail_list_47 : _GEN_110; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_112 = 6'h30 == buf_0_rs2_paddr ? io_avail_list_48 : _GEN_111; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_113 = 6'h31 == buf_0_rs2_paddr ? io_avail_list_49 : _GEN_112; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_114 = 6'h32 == buf_0_rs2_paddr ? io_avail_list_50 : _GEN_113; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_115 = 6'h33 == buf_0_rs2_paddr ? io_avail_list_51 : _GEN_114; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_116 = 6'h34 == buf_0_rs2_paddr ? io_avail_list_52 : _GEN_115; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_117 = 6'h35 == buf_0_rs2_paddr ? io_avail_list_53 : _GEN_116; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_118 = 6'h36 == buf_0_rs2_paddr ? io_avail_list_54 : _GEN_117; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_119 = 6'h37 == buf_0_rs2_paddr ? io_avail_list_55 : _GEN_118; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_120 = 6'h38 == buf_0_rs2_paddr ? io_avail_list_56 : _GEN_119; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_121 = 6'h39 == buf_0_rs2_paddr ? io_avail_list_57 : _GEN_120; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_122 = 6'h3a == buf_0_rs2_paddr ? io_avail_list_58 : _GEN_121; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_123 = 6'h3b == buf_0_rs2_paddr ? io_avail_list_59 : _GEN_122; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_124 = 6'h3c == buf_0_rs2_paddr ? io_avail_list_60 : _GEN_123; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_125 = 6'h3d == buf_0_rs2_paddr ? io_avail_list_61 : _GEN_124; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_126 = 6'h3e == buf_0_rs2_paddr ? io_avail_list_62 : _GEN_125; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_127 = 6'h3f == buf_0_rs2_paddr ? io_avail_list_63 : _GEN_126; // @[IssueUnit.scala 268:{32,32}]
  wire  ready_list_0 = _GEN_63 & _GEN_127 & io_fu_ready; // @[IssueUnit.scala 268:45]
  wire  _GEN_129 = 6'h1 == buf_1_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_130 = 6'h2 == buf_1_rs1_paddr ? io_avail_list_2 : _GEN_129; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_131 = 6'h3 == buf_1_rs1_paddr ? io_avail_list_3 : _GEN_130; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_132 = 6'h4 == buf_1_rs1_paddr ? io_avail_list_4 : _GEN_131; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_133 = 6'h5 == buf_1_rs1_paddr ? io_avail_list_5 : _GEN_132; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_134 = 6'h6 == buf_1_rs1_paddr ? io_avail_list_6 : _GEN_133; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_135 = 6'h7 == buf_1_rs1_paddr ? io_avail_list_7 : _GEN_134; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_136 = 6'h8 == buf_1_rs1_paddr ? io_avail_list_8 : _GEN_135; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_137 = 6'h9 == buf_1_rs1_paddr ? io_avail_list_9 : _GEN_136; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_138 = 6'ha == buf_1_rs1_paddr ? io_avail_list_10 : _GEN_137; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_139 = 6'hb == buf_1_rs1_paddr ? io_avail_list_11 : _GEN_138; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_140 = 6'hc == buf_1_rs1_paddr ? io_avail_list_12 : _GEN_139; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_141 = 6'hd == buf_1_rs1_paddr ? io_avail_list_13 : _GEN_140; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_142 = 6'he == buf_1_rs1_paddr ? io_avail_list_14 : _GEN_141; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_143 = 6'hf == buf_1_rs1_paddr ? io_avail_list_15 : _GEN_142; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_144 = 6'h10 == buf_1_rs1_paddr ? io_avail_list_16 : _GEN_143; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_145 = 6'h11 == buf_1_rs1_paddr ? io_avail_list_17 : _GEN_144; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_146 = 6'h12 == buf_1_rs1_paddr ? io_avail_list_18 : _GEN_145; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_147 = 6'h13 == buf_1_rs1_paddr ? io_avail_list_19 : _GEN_146; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_148 = 6'h14 == buf_1_rs1_paddr ? io_avail_list_20 : _GEN_147; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_149 = 6'h15 == buf_1_rs1_paddr ? io_avail_list_21 : _GEN_148; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_150 = 6'h16 == buf_1_rs1_paddr ? io_avail_list_22 : _GEN_149; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_151 = 6'h17 == buf_1_rs1_paddr ? io_avail_list_23 : _GEN_150; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_152 = 6'h18 == buf_1_rs1_paddr ? io_avail_list_24 : _GEN_151; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_153 = 6'h19 == buf_1_rs1_paddr ? io_avail_list_25 : _GEN_152; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_154 = 6'h1a == buf_1_rs1_paddr ? io_avail_list_26 : _GEN_153; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_155 = 6'h1b == buf_1_rs1_paddr ? io_avail_list_27 : _GEN_154; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_156 = 6'h1c == buf_1_rs1_paddr ? io_avail_list_28 : _GEN_155; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_157 = 6'h1d == buf_1_rs1_paddr ? io_avail_list_29 : _GEN_156; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_158 = 6'h1e == buf_1_rs1_paddr ? io_avail_list_30 : _GEN_157; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_159 = 6'h1f == buf_1_rs1_paddr ? io_avail_list_31 : _GEN_158; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_160 = 6'h20 == buf_1_rs1_paddr ? io_avail_list_32 : _GEN_159; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_161 = 6'h21 == buf_1_rs1_paddr ? io_avail_list_33 : _GEN_160; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_162 = 6'h22 == buf_1_rs1_paddr ? io_avail_list_34 : _GEN_161; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_163 = 6'h23 == buf_1_rs1_paddr ? io_avail_list_35 : _GEN_162; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_164 = 6'h24 == buf_1_rs1_paddr ? io_avail_list_36 : _GEN_163; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_165 = 6'h25 == buf_1_rs1_paddr ? io_avail_list_37 : _GEN_164; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_166 = 6'h26 == buf_1_rs1_paddr ? io_avail_list_38 : _GEN_165; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_167 = 6'h27 == buf_1_rs1_paddr ? io_avail_list_39 : _GEN_166; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_168 = 6'h28 == buf_1_rs1_paddr ? io_avail_list_40 : _GEN_167; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_169 = 6'h29 == buf_1_rs1_paddr ? io_avail_list_41 : _GEN_168; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_170 = 6'h2a == buf_1_rs1_paddr ? io_avail_list_42 : _GEN_169; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_171 = 6'h2b == buf_1_rs1_paddr ? io_avail_list_43 : _GEN_170; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_172 = 6'h2c == buf_1_rs1_paddr ? io_avail_list_44 : _GEN_171; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_173 = 6'h2d == buf_1_rs1_paddr ? io_avail_list_45 : _GEN_172; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_174 = 6'h2e == buf_1_rs1_paddr ? io_avail_list_46 : _GEN_173; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_175 = 6'h2f == buf_1_rs1_paddr ? io_avail_list_47 : _GEN_174; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_176 = 6'h30 == buf_1_rs1_paddr ? io_avail_list_48 : _GEN_175; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_177 = 6'h31 == buf_1_rs1_paddr ? io_avail_list_49 : _GEN_176; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_178 = 6'h32 == buf_1_rs1_paddr ? io_avail_list_50 : _GEN_177; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_179 = 6'h33 == buf_1_rs1_paddr ? io_avail_list_51 : _GEN_178; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_180 = 6'h34 == buf_1_rs1_paddr ? io_avail_list_52 : _GEN_179; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_181 = 6'h35 == buf_1_rs1_paddr ? io_avail_list_53 : _GEN_180; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_182 = 6'h36 == buf_1_rs1_paddr ? io_avail_list_54 : _GEN_181; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_183 = 6'h37 == buf_1_rs1_paddr ? io_avail_list_55 : _GEN_182; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_184 = 6'h38 == buf_1_rs1_paddr ? io_avail_list_56 : _GEN_183; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_185 = 6'h39 == buf_1_rs1_paddr ? io_avail_list_57 : _GEN_184; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_186 = 6'h3a == buf_1_rs1_paddr ? io_avail_list_58 : _GEN_185; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_187 = 6'h3b == buf_1_rs1_paddr ? io_avail_list_59 : _GEN_186; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_188 = 6'h3c == buf_1_rs1_paddr ? io_avail_list_60 : _GEN_187; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_189 = 6'h3d == buf_1_rs1_paddr ? io_avail_list_61 : _GEN_188; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_190 = 6'h3e == buf_1_rs1_paddr ? io_avail_list_62 : _GEN_189; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_191 = 6'h3f == buf_1_rs1_paddr ? io_avail_list_63 : _GEN_190; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_193 = 6'h1 == buf_1_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_194 = 6'h2 == buf_1_rs2_paddr ? io_avail_list_2 : _GEN_193; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_195 = 6'h3 == buf_1_rs2_paddr ? io_avail_list_3 : _GEN_194; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_196 = 6'h4 == buf_1_rs2_paddr ? io_avail_list_4 : _GEN_195; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_197 = 6'h5 == buf_1_rs2_paddr ? io_avail_list_5 : _GEN_196; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_198 = 6'h6 == buf_1_rs2_paddr ? io_avail_list_6 : _GEN_197; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_199 = 6'h7 == buf_1_rs2_paddr ? io_avail_list_7 : _GEN_198; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_200 = 6'h8 == buf_1_rs2_paddr ? io_avail_list_8 : _GEN_199; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_201 = 6'h9 == buf_1_rs2_paddr ? io_avail_list_9 : _GEN_200; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_202 = 6'ha == buf_1_rs2_paddr ? io_avail_list_10 : _GEN_201; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_203 = 6'hb == buf_1_rs2_paddr ? io_avail_list_11 : _GEN_202; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_204 = 6'hc == buf_1_rs2_paddr ? io_avail_list_12 : _GEN_203; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_205 = 6'hd == buf_1_rs2_paddr ? io_avail_list_13 : _GEN_204; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_206 = 6'he == buf_1_rs2_paddr ? io_avail_list_14 : _GEN_205; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_207 = 6'hf == buf_1_rs2_paddr ? io_avail_list_15 : _GEN_206; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_208 = 6'h10 == buf_1_rs2_paddr ? io_avail_list_16 : _GEN_207; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_209 = 6'h11 == buf_1_rs2_paddr ? io_avail_list_17 : _GEN_208; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_210 = 6'h12 == buf_1_rs2_paddr ? io_avail_list_18 : _GEN_209; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_211 = 6'h13 == buf_1_rs2_paddr ? io_avail_list_19 : _GEN_210; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_212 = 6'h14 == buf_1_rs2_paddr ? io_avail_list_20 : _GEN_211; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_213 = 6'h15 == buf_1_rs2_paddr ? io_avail_list_21 : _GEN_212; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_214 = 6'h16 == buf_1_rs2_paddr ? io_avail_list_22 : _GEN_213; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_215 = 6'h17 == buf_1_rs2_paddr ? io_avail_list_23 : _GEN_214; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_216 = 6'h18 == buf_1_rs2_paddr ? io_avail_list_24 : _GEN_215; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_217 = 6'h19 == buf_1_rs2_paddr ? io_avail_list_25 : _GEN_216; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_218 = 6'h1a == buf_1_rs2_paddr ? io_avail_list_26 : _GEN_217; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_219 = 6'h1b == buf_1_rs2_paddr ? io_avail_list_27 : _GEN_218; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_220 = 6'h1c == buf_1_rs2_paddr ? io_avail_list_28 : _GEN_219; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_221 = 6'h1d == buf_1_rs2_paddr ? io_avail_list_29 : _GEN_220; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_222 = 6'h1e == buf_1_rs2_paddr ? io_avail_list_30 : _GEN_221; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_223 = 6'h1f == buf_1_rs2_paddr ? io_avail_list_31 : _GEN_222; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_224 = 6'h20 == buf_1_rs2_paddr ? io_avail_list_32 : _GEN_223; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_225 = 6'h21 == buf_1_rs2_paddr ? io_avail_list_33 : _GEN_224; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_226 = 6'h22 == buf_1_rs2_paddr ? io_avail_list_34 : _GEN_225; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_227 = 6'h23 == buf_1_rs2_paddr ? io_avail_list_35 : _GEN_226; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_228 = 6'h24 == buf_1_rs2_paddr ? io_avail_list_36 : _GEN_227; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_229 = 6'h25 == buf_1_rs2_paddr ? io_avail_list_37 : _GEN_228; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_230 = 6'h26 == buf_1_rs2_paddr ? io_avail_list_38 : _GEN_229; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_231 = 6'h27 == buf_1_rs2_paddr ? io_avail_list_39 : _GEN_230; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_232 = 6'h28 == buf_1_rs2_paddr ? io_avail_list_40 : _GEN_231; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_233 = 6'h29 == buf_1_rs2_paddr ? io_avail_list_41 : _GEN_232; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_234 = 6'h2a == buf_1_rs2_paddr ? io_avail_list_42 : _GEN_233; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_235 = 6'h2b == buf_1_rs2_paddr ? io_avail_list_43 : _GEN_234; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_236 = 6'h2c == buf_1_rs2_paddr ? io_avail_list_44 : _GEN_235; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_237 = 6'h2d == buf_1_rs2_paddr ? io_avail_list_45 : _GEN_236; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_238 = 6'h2e == buf_1_rs2_paddr ? io_avail_list_46 : _GEN_237; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_239 = 6'h2f == buf_1_rs2_paddr ? io_avail_list_47 : _GEN_238; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_240 = 6'h30 == buf_1_rs2_paddr ? io_avail_list_48 : _GEN_239; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_241 = 6'h31 == buf_1_rs2_paddr ? io_avail_list_49 : _GEN_240; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_242 = 6'h32 == buf_1_rs2_paddr ? io_avail_list_50 : _GEN_241; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_243 = 6'h33 == buf_1_rs2_paddr ? io_avail_list_51 : _GEN_242; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_244 = 6'h34 == buf_1_rs2_paddr ? io_avail_list_52 : _GEN_243; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_245 = 6'h35 == buf_1_rs2_paddr ? io_avail_list_53 : _GEN_244; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_246 = 6'h36 == buf_1_rs2_paddr ? io_avail_list_54 : _GEN_245; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_247 = 6'h37 == buf_1_rs2_paddr ? io_avail_list_55 : _GEN_246; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_248 = 6'h38 == buf_1_rs2_paddr ? io_avail_list_56 : _GEN_247; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_249 = 6'h39 == buf_1_rs2_paddr ? io_avail_list_57 : _GEN_248; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_250 = 6'h3a == buf_1_rs2_paddr ? io_avail_list_58 : _GEN_249; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_251 = 6'h3b == buf_1_rs2_paddr ? io_avail_list_59 : _GEN_250; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_252 = 6'h3c == buf_1_rs2_paddr ? io_avail_list_60 : _GEN_251; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_253 = 6'h3d == buf_1_rs2_paddr ? io_avail_list_61 : _GEN_252; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_254 = 6'h3e == buf_1_rs2_paddr ? io_avail_list_62 : _GEN_253; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_255 = 6'h3f == buf_1_rs2_paddr ? io_avail_list_63 : _GEN_254; // @[IssueUnit.scala 268:{32,32}]
  wire  ready_list_1 = _GEN_191 & _GEN_255 & io_fu_ready & store_mask_1; // @[IssueUnit.scala 268:57]
  wire  _GEN_257 = 6'h1 == buf_2_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_258 = 6'h2 == buf_2_rs1_paddr ? io_avail_list_2 : _GEN_257; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_259 = 6'h3 == buf_2_rs1_paddr ? io_avail_list_3 : _GEN_258; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_260 = 6'h4 == buf_2_rs1_paddr ? io_avail_list_4 : _GEN_259; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_261 = 6'h5 == buf_2_rs1_paddr ? io_avail_list_5 : _GEN_260; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_262 = 6'h6 == buf_2_rs1_paddr ? io_avail_list_6 : _GEN_261; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_263 = 6'h7 == buf_2_rs1_paddr ? io_avail_list_7 : _GEN_262; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_264 = 6'h8 == buf_2_rs1_paddr ? io_avail_list_8 : _GEN_263; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_265 = 6'h9 == buf_2_rs1_paddr ? io_avail_list_9 : _GEN_264; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_266 = 6'ha == buf_2_rs1_paddr ? io_avail_list_10 : _GEN_265; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_267 = 6'hb == buf_2_rs1_paddr ? io_avail_list_11 : _GEN_266; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_268 = 6'hc == buf_2_rs1_paddr ? io_avail_list_12 : _GEN_267; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_269 = 6'hd == buf_2_rs1_paddr ? io_avail_list_13 : _GEN_268; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_270 = 6'he == buf_2_rs1_paddr ? io_avail_list_14 : _GEN_269; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_271 = 6'hf == buf_2_rs1_paddr ? io_avail_list_15 : _GEN_270; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_272 = 6'h10 == buf_2_rs1_paddr ? io_avail_list_16 : _GEN_271; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_273 = 6'h11 == buf_2_rs1_paddr ? io_avail_list_17 : _GEN_272; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_274 = 6'h12 == buf_2_rs1_paddr ? io_avail_list_18 : _GEN_273; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_275 = 6'h13 == buf_2_rs1_paddr ? io_avail_list_19 : _GEN_274; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_276 = 6'h14 == buf_2_rs1_paddr ? io_avail_list_20 : _GEN_275; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_277 = 6'h15 == buf_2_rs1_paddr ? io_avail_list_21 : _GEN_276; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_278 = 6'h16 == buf_2_rs1_paddr ? io_avail_list_22 : _GEN_277; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_279 = 6'h17 == buf_2_rs1_paddr ? io_avail_list_23 : _GEN_278; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_280 = 6'h18 == buf_2_rs1_paddr ? io_avail_list_24 : _GEN_279; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_281 = 6'h19 == buf_2_rs1_paddr ? io_avail_list_25 : _GEN_280; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_282 = 6'h1a == buf_2_rs1_paddr ? io_avail_list_26 : _GEN_281; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_283 = 6'h1b == buf_2_rs1_paddr ? io_avail_list_27 : _GEN_282; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_284 = 6'h1c == buf_2_rs1_paddr ? io_avail_list_28 : _GEN_283; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_285 = 6'h1d == buf_2_rs1_paddr ? io_avail_list_29 : _GEN_284; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_286 = 6'h1e == buf_2_rs1_paddr ? io_avail_list_30 : _GEN_285; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_287 = 6'h1f == buf_2_rs1_paddr ? io_avail_list_31 : _GEN_286; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_288 = 6'h20 == buf_2_rs1_paddr ? io_avail_list_32 : _GEN_287; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_289 = 6'h21 == buf_2_rs1_paddr ? io_avail_list_33 : _GEN_288; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_290 = 6'h22 == buf_2_rs1_paddr ? io_avail_list_34 : _GEN_289; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_291 = 6'h23 == buf_2_rs1_paddr ? io_avail_list_35 : _GEN_290; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_292 = 6'h24 == buf_2_rs1_paddr ? io_avail_list_36 : _GEN_291; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_293 = 6'h25 == buf_2_rs1_paddr ? io_avail_list_37 : _GEN_292; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_294 = 6'h26 == buf_2_rs1_paddr ? io_avail_list_38 : _GEN_293; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_295 = 6'h27 == buf_2_rs1_paddr ? io_avail_list_39 : _GEN_294; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_296 = 6'h28 == buf_2_rs1_paddr ? io_avail_list_40 : _GEN_295; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_297 = 6'h29 == buf_2_rs1_paddr ? io_avail_list_41 : _GEN_296; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_298 = 6'h2a == buf_2_rs1_paddr ? io_avail_list_42 : _GEN_297; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_299 = 6'h2b == buf_2_rs1_paddr ? io_avail_list_43 : _GEN_298; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_300 = 6'h2c == buf_2_rs1_paddr ? io_avail_list_44 : _GEN_299; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_301 = 6'h2d == buf_2_rs1_paddr ? io_avail_list_45 : _GEN_300; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_302 = 6'h2e == buf_2_rs1_paddr ? io_avail_list_46 : _GEN_301; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_303 = 6'h2f == buf_2_rs1_paddr ? io_avail_list_47 : _GEN_302; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_304 = 6'h30 == buf_2_rs1_paddr ? io_avail_list_48 : _GEN_303; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_305 = 6'h31 == buf_2_rs1_paddr ? io_avail_list_49 : _GEN_304; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_306 = 6'h32 == buf_2_rs1_paddr ? io_avail_list_50 : _GEN_305; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_307 = 6'h33 == buf_2_rs1_paddr ? io_avail_list_51 : _GEN_306; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_308 = 6'h34 == buf_2_rs1_paddr ? io_avail_list_52 : _GEN_307; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_309 = 6'h35 == buf_2_rs1_paddr ? io_avail_list_53 : _GEN_308; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_310 = 6'h36 == buf_2_rs1_paddr ? io_avail_list_54 : _GEN_309; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_311 = 6'h37 == buf_2_rs1_paddr ? io_avail_list_55 : _GEN_310; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_312 = 6'h38 == buf_2_rs1_paddr ? io_avail_list_56 : _GEN_311; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_313 = 6'h39 == buf_2_rs1_paddr ? io_avail_list_57 : _GEN_312; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_314 = 6'h3a == buf_2_rs1_paddr ? io_avail_list_58 : _GEN_313; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_315 = 6'h3b == buf_2_rs1_paddr ? io_avail_list_59 : _GEN_314; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_316 = 6'h3c == buf_2_rs1_paddr ? io_avail_list_60 : _GEN_315; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_317 = 6'h3d == buf_2_rs1_paddr ? io_avail_list_61 : _GEN_316; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_318 = 6'h3e == buf_2_rs1_paddr ? io_avail_list_62 : _GEN_317; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_319 = 6'h3f == buf_2_rs1_paddr ? io_avail_list_63 : _GEN_318; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_321 = 6'h1 == buf_2_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_322 = 6'h2 == buf_2_rs2_paddr ? io_avail_list_2 : _GEN_321; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_323 = 6'h3 == buf_2_rs2_paddr ? io_avail_list_3 : _GEN_322; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_324 = 6'h4 == buf_2_rs2_paddr ? io_avail_list_4 : _GEN_323; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_325 = 6'h5 == buf_2_rs2_paddr ? io_avail_list_5 : _GEN_324; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_326 = 6'h6 == buf_2_rs2_paddr ? io_avail_list_6 : _GEN_325; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_327 = 6'h7 == buf_2_rs2_paddr ? io_avail_list_7 : _GEN_326; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_328 = 6'h8 == buf_2_rs2_paddr ? io_avail_list_8 : _GEN_327; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_329 = 6'h9 == buf_2_rs2_paddr ? io_avail_list_9 : _GEN_328; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_330 = 6'ha == buf_2_rs2_paddr ? io_avail_list_10 : _GEN_329; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_331 = 6'hb == buf_2_rs2_paddr ? io_avail_list_11 : _GEN_330; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_332 = 6'hc == buf_2_rs2_paddr ? io_avail_list_12 : _GEN_331; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_333 = 6'hd == buf_2_rs2_paddr ? io_avail_list_13 : _GEN_332; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_334 = 6'he == buf_2_rs2_paddr ? io_avail_list_14 : _GEN_333; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_335 = 6'hf == buf_2_rs2_paddr ? io_avail_list_15 : _GEN_334; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_336 = 6'h10 == buf_2_rs2_paddr ? io_avail_list_16 : _GEN_335; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_337 = 6'h11 == buf_2_rs2_paddr ? io_avail_list_17 : _GEN_336; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_338 = 6'h12 == buf_2_rs2_paddr ? io_avail_list_18 : _GEN_337; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_339 = 6'h13 == buf_2_rs2_paddr ? io_avail_list_19 : _GEN_338; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_340 = 6'h14 == buf_2_rs2_paddr ? io_avail_list_20 : _GEN_339; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_341 = 6'h15 == buf_2_rs2_paddr ? io_avail_list_21 : _GEN_340; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_342 = 6'h16 == buf_2_rs2_paddr ? io_avail_list_22 : _GEN_341; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_343 = 6'h17 == buf_2_rs2_paddr ? io_avail_list_23 : _GEN_342; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_344 = 6'h18 == buf_2_rs2_paddr ? io_avail_list_24 : _GEN_343; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_345 = 6'h19 == buf_2_rs2_paddr ? io_avail_list_25 : _GEN_344; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_346 = 6'h1a == buf_2_rs2_paddr ? io_avail_list_26 : _GEN_345; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_347 = 6'h1b == buf_2_rs2_paddr ? io_avail_list_27 : _GEN_346; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_348 = 6'h1c == buf_2_rs2_paddr ? io_avail_list_28 : _GEN_347; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_349 = 6'h1d == buf_2_rs2_paddr ? io_avail_list_29 : _GEN_348; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_350 = 6'h1e == buf_2_rs2_paddr ? io_avail_list_30 : _GEN_349; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_351 = 6'h1f == buf_2_rs2_paddr ? io_avail_list_31 : _GEN_350; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_352 = 6'h20 == buf_2_rs2_paddr ? io_avail_list_32 : _GEN_351; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_353 = 6'h21 == buf_2_rs2_paddr ? io_avail_list_33 : _GEN_352; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_354 = 6'h22 == buf_2_rs2_paddr ? io_avail_list_34 : _GEN_353; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_355 = 6'h23 == buf_2_rs2_paddr ? io_avail_list_35 : _GEN_354; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_356 = 6'h24 == buf_2_rs2_paddr ? io_avail_list_36 : _GEN_355; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_357 = 6'h25 == buf_2_rs2_paddr ? io_avail_list_37 : _GEN_356; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_358 = 6'h26 == buf_2_rs2_paddr ? io_avail_list_38 : _GEN_357; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_359 = 6'h27 == buf_2_rs2_paddr ? io_avail_list_39 : _GEN_358; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_360 = 6'h28 == buf_2_rs2_paddr ? io_avail_list_40 : _GEN_359; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_361 = 6'h29 == buf_2_rs2_paddr ? io_avail_list_41 : _GEN_360; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_362 = 6'h2a == buf_2_rs2_paddr ? io_avail_list_42 : _GEN_361; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_363 = 6'h2b == buf_2_rs2_paddr ? io_avail_list_43 : _GEN_362; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_364 = 6'h2c == buf_2_rs2_paddr ? io_avail_list_44 : _GEN_363; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_365 = 6'h2d == buf_2_rs2_paddr ? io_avail_list_45 : _GEN_364; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_366 = 6'h2e == buf_2_rs2_paddr ? io_avail_list_46 : _GEN_365; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_367 = 6'h2f == buf_2_rs2_paddr ? io_avail_list_47 : _GEN_366; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_368 = 6'h30 == buf_2_rs2_paddr ? io_avail_list_48 : _GEN_367; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_369 = 6'h31 == buf_2_rs2_paddr ? io_avail_list_49 : _GEN_368; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_370 = 6'h32 == buf_2_rs2_paddr ? io_avail_list_50 : _GEN_369; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_371 = 6'h33 == buf_2_rs2_paddr ? io_avail_list_51 : _GEN_370; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_372 = 6'h34 == buf_2_rs2_paddr ? io_avail_list_52 : _GEN_371; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_373 = 6'h35 == buf_2_rs2_paddr ? io_avail_list_53 : _GEN_372; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_374 = 6'h36 == buf_2_rs2_paddr ? io_avail_list_54 : _GEN_373; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_375 = 6'h37 == buf_2_rs2_paddr ? io_avail_list_55 : _GEN_374; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_376 = 6'h38 == buf_2_rs2_paddr ? io_avail_list_56 : _GEN_375; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_377 = 6'h39 == buf_2_rs2_paddr ? io_avail_list_57 : _GEN_376; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_378 = 6'h3a == buf_2_rs2_paddr ? io_avail_list_58 : _GEN_377; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_379 = 6'h3b == buf_2_rs2_paddr ? io_avail_list_59 : _GEN_378; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_380 = 6'h3c == buf_2_rs2_paddr ? io_avail_list_60 : _GEN_379; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_381 = 6'h3d == buf_2_rs2_paddr ? io_avail_list_61 : _GEN_380; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_382 = 6'h3e == buf_2_rs2_paddr ? io_avail_list_62 : _GEN_381; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_383 = 6'h3f == buf_2_rs2_paddr ? io_avail_list_63 : _GEN_382; // @[IssueUnit.scala 268:{32,32}]
  wire  ready_list_2 = _GEN_319 & _GEN_383 & io_fu_ready & store_mask_2; // @[IssueUnit.scala 268:57]
  wire  _GEN_385 = 6'h1 == buf_3_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_386 = 6'h2 == buf_3_rs1_paddr ? io_avail_list_2 : _GEN_385; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_387 = 6'h3 == buf_3_rs1_paddr ? io_avail_list_3 : _GEN_386; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_388 = 6'h4 == buf_3_rs1_paddr ? io_avail_list_4 : _GEN_387; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_389 = 6'h5 == buf_3_rs1_paddr ? io_avail_list_5 : _GEN_388; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_390 = 6'h6 == buf_3_rs1_paddr ? io_avail_list_6 : _GEN_389; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_391 = 6'h7 == buf_3_rs1_paddr ? io_avail_list_7 : _GEN_390; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_392 = 6'h8 == buf_3_rs1_paddr ? io_avail_list_8 : _GEN_391; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_393 = 6'h9 == buf_3_rs1_paddr ? io_avail_list_9 : _GEN_392; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_394 = 6'ha == buf_3_rs1_paddr ? io_avail_list_10 : _GEN_393; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_395 = 6'hb == buf_3_rs1_paddr ? io_avail_list_11 : _GEN_394; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_396 = 6'hc == buf_3_rs1_paddr ? io_avail_list_12 : _GEN_395; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_397 = 6'hd == buf_3_rs1_paddr ? io_avail_list_13 : _GEN_396; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_398 = 6'he == buf_3_rs1_paddr ? io_avail_list_14 : _GEN_397; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_399 = 6'hf == buf_3_rs1_paddr ? io_avail_list_15 : _GEN_398; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_400 = 6'h10 == buf_3_rs1_paddr ? io_avail_list_16 : _GEN_399; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_401 = 6'h11 == buf_3_rs1_paddr ? io_avail_list_17 : _GEN_400; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_402 = 6'h12 == buf_3_rs1_paddr ? io_avail_list_18 : _GEN_401; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_403 = 6'h13 == buf_3_rs1_paddr ? io_avail_list_19 : _GEN_402; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_404 = 6'h14 == buf_3_rs1_paddr ? io_avail_list_20 : _GEN_403; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_405 = 6'h15 == buf_3_rs1_paddr ? io_avail_list_21 : _GEN_404; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_406 = 6'h16 == buf_3_rs1_paddr ? io_avail_list_22 : _GEN_405; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_407 = 6'h17 == buf_3_rs1_paddr ? io_avail_list_23 : _GEN_406; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_408 = 6'h18 == buf_3_rs1_paddr ? io_avail_list_24 : _GEN_407; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_409 = 6'h19 == buf_3_rs1_paddr ? io_avail_list_25 : _GEN_408; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_410 = 6'h1a == buf_3_rs1_paddr ? io_avail_list_26 : _GEN_409; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_411 = 6'h1b == buf_3_rs1_paddr ? io_avail_list_27 : _GEN_410; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_412 = 6'h1c == buf_3_rs1_paddr ? io_avail_list_28 : _GEN_411; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_413 = 6'h1d == buf_3_rs1_paddr ? io_avail_list_29 : _GEN_412; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_414 = 6'h1e == buf_3_rs1_paddr ? io_avail_list_30 : _GEN_413; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_415 = 6'h1f == buf_3_rs1_paddr ? io_avail_list_31 : _GEN_414; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_416 = 6'h20 == buf_3_rs1_paddr ? io_avail_list_32 : _GEN_415; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_417 = 6'h21 == buf_3_rs1_paddr ? io_avail_list_33 : _GEN_416; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_418 = 6'h22 == buf_3_rs1_paddr ? io_avail_list_34 : _GEN_417; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_419 = 6'h23 == buf_3_rs1_paddr ? io_avail_list_35 : _GEN_418; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_420 = 6'h24 == buf_3_rs1_paddr ? io_avail_list_36 : _GEN_419; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_421 = 6'h25 == buf_3_rs1_paddr ? io_avail_list_37 : _GEN_420; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_422 = 6'h26 == buf_3_rs1_paddr ? io_avail_list_38 : _GEN_421; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_423 = 6'h27 == buf_3_rs1_paddr ? io_avail_list_39 : _GEN_422; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_424 = 6'h28 == buf_3_rs1_paddr ? io_avail_list_40 : _GEN_423; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_425 = 6'h29 == buf_3_rs1_paddr ? io_avail_list_41 : _GEN_424; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_426 = 6'h2a == buf_3_rs1_paddr ? io_avail_list_42 : _GEN_425; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_427 = 6'h2b == buf_3_rs1_paddr ? io_avail_list_43 : _GEN_426; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_428 = 6'h2c == buf_3_rs1_paddr ? io_avail_list_44 : _GEN_427; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_429 = 6'h2d == buf_3_rs1_paddr ? io_avail_list_45 : _GEN_428; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_430 = 6'h2e == buf_3_rs1_paddr ? io_avail_list_46 : _GEN_429; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_431 = 6'h2f == buf_3_rs1_paddr ? io_avail_list_47 : _GEN_430; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_432 = 6'h30 == buf_3_rs1_paddr ? io_avail_list_48 : _GEN_431; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_433 = 6'h31 == buf_3_rs1_paddr ? io_avail_list_49 : _GEN_432; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_434 = 6'h32 == buf_3_rs1_paddr ? io_avail_list_50 : _GEN_433; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_435 = 6'h33 == buf_3_rs1_paddr ? io_avail_list_51 : _GEN_434; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_436 = 6'h34 == buf_3_rs1_paddr ? io_avail_list_52 : _GEN_435; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_437 = 6'h35 == buf_3_rs1_paddr ? io_avail_list_53 : _GEN_436; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_438 = 6'h36 == buf_3_rs1_paddr ? io_avail_list_54 : _GEN_437; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_439 = 6'h37 == buf_3_rs1_paddr ? io_avail_list_55 : _GEN_438; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_440 = 6'h38 == buf_3_rs1_paddr ? io_avail_list_56 : _GEN_439; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_441 = 6'h39 == buf_3_rs1_paddr ? io_avail_list_57 : _GEN_440; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_442 = 6'h3a == buf_3_rs1_paddr ? io_avail_list_58 : _GEN_441; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_443 = 6'h3b == buf_3_rs1_paddr ? io_avail_list_59 : _GEN_442; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_444 = 6'h3c == buf_3_rs1_paddr ? io_avail_list_60 : _GEN_443; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_445 = 6'h3d == buf_3_rs1_paddr ? io_avail_list_61 : _GEN_444; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_446 = 6'h3e == buf_3_rs1_paddr ? io_avail_list_62 : _GEN_445; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_447 = 6'h3f == buf_3_rs1_paddr ? io_avail_list_63 : _GEN_446; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_449 = 6'h1 == buf_3_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_450 = 6'h2 == buf_3_rs2_paddr ? io_avail_list_2 : _GEN_449; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_451 = 6'h3 == buf_3_rs2_paddr ? io_avail_list_3 : _GEN_450; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_452 = 6'h4 == buf_3_rs2_paddr ? io_avail_list_4 : _GEN_451; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_453 = 6'h5 == buf_3_rs2_paddr ? io_avail_list_5 : _GEN_452; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_454 = 6'h6 == buf_3_rs2_paddr ? io_avail_list_6 : _GEN_453; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_455 = 6'h7 == buf_3_rs2_paddr ? io_avail_list_7 : _GEN_454; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_456 = 6'h8 == buf_3_rs2_paddr ? io_avail_list_8 : _GEN_455; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_457 = 6'h9 == buf_3_rs2_paddr ? io_avail_list_9 : _GEN_456; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_458 = 6'ha == buf_3_rs2_paddr ? io_avail_list_10 : _GEN_457; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_459 = 6'hb == buf_3_rs2_paddr ? io_avail_list_11 : _GEN_458; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_460 = 6'hc == buf_3_rs2_paddr ? io_avail_list_12 : _GEN_459; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_461 = 6'hd == buf_3_rs2_paddr ? io_avail_list_13 : _GEN_460; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_462 = 6'he == buf_3_rs2_paddr ? io_avail_list_14 : _GEN_461; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_463 = 6'hf == buf_3_rs2_paddr ? io_avail_list_15 : _GEN_462; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_464 = 6'h10 == buf_3_rs2_paddr ? io_avail_list_16 : _GEN_463; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_465 = 6'h11 == buf_3_rs2_paddr ? io_avail_list_17 : _GEN_464; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_466 = 6'h12 == buf_3_rs2_paddr ? io_avail_list_18 : _GEN_465; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_467 = 6'h13 == buf_3_rs2_paddr ? io_avail_list_19 : _GEN_466; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_468 = 6'h14 == buf_3_rs2_paddr ? io_avail_list_20 : _GEN_467; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_469 = 6'h15 == buf_3_rs2_paddr ? io_avail_list_21 : _GEN_468; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_470 = 6'h16 == buf_3_rs2_paddr ? io_avail_list_22 : _GEN_469; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_471 = 6'h17 == buf_3_rs2_paddr ? io_avail_list_23 : _GEN_470; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_472 = 6'h18 == buf_3_rs2_paddr ? io_avail_list_24 : _GEN_471; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_473 = 6'h19 == buf_3_rs2_paddr ? io_avail_list_25 : _GEN_472; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_474 = 6'h1a == buf_3_rs2_paddr ? io_avail_list_26 : _GEN_473; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_475 = 6'h1b == buf_3_rs2_paddr ? io_avail_list_27 : _GEN_474; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_476 = 6'h1c == buf_3_rs2_paddr ? io_avail_list_28 : _GEN_475; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_477 = 6'h1d == buf_3_rs2_paddr ? io_avail_list_29 : _GEN_476; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_478 = 6'h1e == buf_3_rs2_paddr ? io_avail_list_30 : _GEN_477; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_479 = 6'h1f == buf_3_rs2_paddr ? io_avail_list_31 : _GEN_478; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_480 = 6'h20 == buf_3_rs2_paddr ? io_avail_list_32 : _GEN_479; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_481 = 6'h21 == buf_3_rs2_paddr ? io_avail_list_33 : _GEN_480; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_482 = 6'h22 == buf_3_rs2_paddr ? io_avail_list_34 : _GEN_481; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_483 = 6'h23 == buf_3_rs2_paddr ? io_avail_list_35 : _GEN_482; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_484 = 6'h24 == buf_3_rs2_paddr ? io_avail_list_36 : _GEN_483; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_485 = 6'h25 == buf_3_rs2_paddr ? io_avail_list_37 : _GEN_484; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_486 = 6'h26 == buf_3_rs2_paddr ? io_avail_list_38 : _GEN_485; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_487 = 6'h27 == buf_3_rs2_paddr ? io_avail_list_39 : _GEN_486; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_488 = 6'h28 == buf_3_rs2_paddr ? io_avail_list_40 : _GEN_487; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_489 = 6'h29 == buf_3_rs2_paddr ? io_avail_list_41 : _GEN_488; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_490 = 6'h2a == buf_3_rs2_paddr ? io_avail_list_42 : _GEN_489; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_491 = 6'h2b == buf_3_rs2_paddr ? io_avail_list_43 : _GEN_490; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_492 = 6'h2c == buf_3_rs2_paddr ? io_avail_list_44 : _GEN_491; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_493 = 6'h2d == buf_3_rs2_paddr ? io_avail_list_45 : _GEN_492; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_494 = 6'h2e == buf_3_rs2_paddr ? io_avail_list_46 : _GEN_493; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_495 = 6'h2f == buf_3_rs2_paddr ? io_avail_list_47 : _GEN_494; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_496 = 6'h30 == buf_3_rs2_paddr ? io_avail_list_48 : _GEN_495; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_497 = 6'h31 == buf_3_rs2_paddr ? io_avail_list_49 : _GEN_496; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_498 = 6'h32 == buf_3_rs2_paddr ? io_avail_list_50 : _GEN_497; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_499 = 6'h33 == buf_3_rs2_paddr ? io_avail_list_51 : _GEN_498; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_500 = 6'h34 == buf_3_rs2_paddr ? io_avail_list_52 : _GEN_499; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_501 = 6'h35 == buf_3_rs2_paddr ? io_avail_list_53 : _GEN_500; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_502 = 6'h36 == buf_3_rs2_paddr ? io_avail_list_54 : _GEN_501; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_503 = 6'h37 == buf_3_rs2_paddr ? io_avail_list_55 : _GEN_502; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_504 = 6'h38 == buf_3_rs2_paddr ? io_avail_list_56 : _GEN_503; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_505 = 6'h39 == buf_3_rs2_paddr ? io_avail_list_57 : _GEN_504; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_506 = 6'h3a == buf_3_rs2_paddr ? io_avail_list_58 : _GEN_505; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_507 = 6'h3b == buf_3_rs2_paddr ? io_avail_list_59 : _GEN_506; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_508 = 6'h3c == buf_3_rs2_paddr ? io_avail_list_60 : _GEN_507; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_509 = 6'h3d == buf_3_rs2_paddr ? io_avail_list_61 : _GEN_508; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_510 = 6'h3e == buf_3_rs2_paddr ? io_avail_list_62 : _GEN_509; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_511 = 6'h3f == buf_3_rs2_paddr ? io_avail_list_63 : _GEN_510; // @[IssueUnit.scala 268:{32,32}]
  wire  ready_list_3 = _GEN_447 & _GEN_511 & io_fu_ready & store_mask_3; // @[IssueUnit.scala 268:57]
  wire  _GEN_513 = 6'h1 == buf_4_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_514 = 6'h2 == buf_4_rs1_paddr ? io_avail_list_2 : _GEN_513; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_515 = 6'h3 == buf_4_rs1_paddr ? io_avail_list_3 : _GEN_514; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_516 = 6'h4 == buf_4_rs1_paddr ? io_avail_list_4 : _GEN_515; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_517 = 6'h5 == buf_4_rs1_paddr ? io_avail_list_5 : _GEN_516; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_518 = 6'h6 == buf_4_rs1_paddr ? io_avail_list_6 : _GEN_517; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_519 = 6'h7 == buf_4_rs1_paddr ? io_avail_list_7 : _GEN_518; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_520 = 6'h8 == buf_4_rs1_paddr ? io_avail_list_8 : _GEN_519; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_521 = 6'h9 == buf_4_rs1_paddr ? io_avail_list_9 : _GEN_520; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_522 = 6'ha == buf_4_rs1_paddr ? io_avail_list_10 : _GEN_521; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_523 = 6'hb == buf_4_rs1_paddr ? io_avail_list_11 : _GEN_522; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_524 = 6'hc == buf_4_rs1_paddr ? io_avail_list_12 : _GEN_523; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_525 = 6'hd == buf_4_rs1_paddr ? io_avail_list_13 : _GEN_524; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_526 = 6'he == buf_4_rs1_paddr ? io_avail_list_14 : _GEN_525; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_527 = 6'hf == buf_4_rs1_paddr ? io_avail_list_15 : _GEN_526; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_528 = 6'h10 == buf_4_rs1_paddr ? io_avail_list_16 : _GEN_527; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_529 = 6'h11 == buf_4_rs1_paddr ? io_avail_list_17 : _GEN_528; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_530 = 6'h12 == buf_4_rs1_paddr ? io_avail_list_18 : _GEN_529; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_531 = 6'h13 == buf_4_rs1_paddr ? io_avail_list_19 : _GEN_530; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_532 = 6'h14 == buf_4_rs1_paddr ? io_avail_list_20 : _GEN_531; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_533 = 6'h15 == buf_4_rs1_paddr ? io_avail_list_21 : _GEN_532; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_534 = 6'h16 == buf_4_rs1_paddr ? io_avail_list_22 : _GEN_533; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_535 = 6'h17 == buf_4_rs1_paddr ? io_avail_list_23 : _GEN_534; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_536 = 6'h18 == buf_4_rs1_paddr ? io_avail_list_24 : _GEN_535; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_537 = 6'h19 == buf_4_rs1_paddr ? io_avail_list_25 : _GEN_536; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_538 = 6'h1a == buf_4_rs1_paddr ? io_avail_list_26 : _GEN_537; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_539 = 6'h1b == buf_4_rs1_paddr ? io_avail_list_27 : _GEN_538; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_540 = 6'h1c == buf_4_rs1_paddr ? io_avail_list_28 : _GEN_539; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_541 = 6'h1d == buf_4_rs1_paddr ? io_avail_list_29 : _GEN_540; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_542 = 6'h1e == buf_4_rs1_paddr ? io_avail_list_30 : _GEN_541; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_543 = 6'h1f == buf_4_rs1_paddr ? io_avail_list_31 : _GEN_542; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_544 = 6'h20 == buf_4_rs1_paddr ? io_avail_list_32 : _GEN_543; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_545 = 6'h21 == buf_4_rs1_paddr ? io_avail_list_33 : _GEN_544; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_546 = 6'h22 == buf_4_rs1_paddr ? io_avail_list_34 : _GEN_545; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_547 = 6'h23 == buf_4_rs1_paddr ? io_avail_list_35 : _GEN_546; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_548 = 6'h24 == buf_4_rs1_paddr ? io_avail_list_36 : _GEN_547; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_549 = 6'h25 == buf_4_rs1_paddr ? io_avail_list_37 : _GEN_548; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_550 = 6'h26 == buf_4_rs1_paddr ? io_avail_list_38 : _GEN_549; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_551 = 6'h27 == buf_4_rs1_paddr ? io_avail_list_39 : _GEN_550; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_552 = 6'h28 == buf_4_rs1_paddr ? io_avail_list_40 : _GEN_551; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_553 = 6'h29 == buf_4_rs1_paddr ? io_avail_list_41 : _GEN_552; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_554 = 6'h2a == buf_4_rs1_paddr ? io_avail_list_42 : _GEN_553; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_555 = 6'h2b == buf_4_rs1_paddr ? io_avail_list_43 : _GEN_554; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_556 = 6'h2c == buf_4_rs1_paddr ? io_avail_list_44 : _GEN_555; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_557 = 6'h2d == buf_4_rs1_paddr ? io_avail_list_45 : _GEN_556; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_558 = 6'h2e == buf_4_rs1_paddr ? io_avail_list_46 : _GEN_557; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_559 = 6'h2f == buf_4_rs1_paddr ? io_avail_list_47 : _GEN_558; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_560 = 6'h30 == buf_4_rs1_paddr ? io_avail_list_48 : _GEN_559; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_561 = 6'h31 == buf_4_rs1_paddr ? io_avail_list_49 : _GEN_560; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_562 = 6'h32 == buf_4_rs1_paddr ? io_avail_list_50 : _GEN_561; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_563 = 6'h33 == buf_4_rs1_paddr ? io_avail_list_51 : _GEN_562; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_564 = 6'h34 == buf_4_rs1_paddr ? io_avail_list_52 : _GEN_563; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_565 = 6'h35 == buf_4_rs1_paddr ? io_avail_list_53 : _GEN_564; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_566 = 6'h36 == buf_4_rs1_paddr ? io_avail_list_54 : _GEN_565; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_567 = 6'h37 == buf_4_rs1_paddr ? io_avail_list_55 : _GEN_566; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_568 = 6'h38 == buf_4_rs1_paddr ? io_avail_list_56 : _GEN_567; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_569 = 6'h39 == buf_4_rs1_paddr ? io_avail_list_57 : _GEN_568; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_570 = 6'h3a == buf_4_rs1_paddr ? io_avail_list_58 : _GEN_569; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_571 = 6'h3b == buf_4_rs1_paddr ? io_avail_list_59 : _GEN_570; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_572 = 6'h3c == buf_4_rs1_paddr ? io_avail_list_60 : _GEN_571; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_573 = 6'h3d == buf_4_rs1_paddr ? io_avail_list_61 : _GEN_572; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_574 = 6'h3e == buf_4_rs1_paddr ? io_avail_list_62 : _GEN_573; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_575 = 6'h3f == buf_4_rs1_paddr ? io_avail_list_63 : _GEN_574; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_577 = 6'h1 == buf_4_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_578 = 6'h2 == buf_4_rs2_paddr ? io_avail_list_2 : _GEN_577; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_579 = 6'h3 == buf_4_rs2_paddr ? io_avail_list_3 : _GEN_578; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_580 = 6'h4 == buf_4_rs2_paddr ? io_avail_list_4 : _GEN_579; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_581 = 6'h5 == buf_4_rs2_paddr ? io_avail_list_5 : _GEN_580; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_582 = 6'h6 == buf_4_rs2_paddr ? io_avail_list_6 : _GEN_581; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_583 = 6'h7 == buf_4_rs2_paddr ? io_avail_list_7 : _GEN_582; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_584 = 6'h8 == buf_4_rs2_paddr ? io_avail_list_8 : _GEN_583; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_585 = 6'h9 == buf_4_rs2_paddr ? io_avail_list_9 : _GEN_584; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_586 = 6'ha == buf_4_rs2_paddr ? io_avail_list_10 : _GEN_585; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_587 = 6'hb == buf_4_rs2_paddr ? io_avail_list_11 : _GEN_586; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_588 = 6'hc == buf_4_rs2_paddr ? io_avail_list_12 : _GEN_587; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_589 = 6'hd == buf_4_rs2_paddr ? io_avail_list_13 : _GEN_588; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_590 = 6'he == buf_4_rs2_paddr ? io_avail_list_14 : _GEN_589; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_591 = 6'hf == buf_4_rs2_paddr ? io_avail_list_15 : _GEN_590; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_592 = 6'h10 == buf_4_rs2_paddr ? io_avail_list_16 : _GEN_591; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_593 = 6'h11 == buf_4_rs2_paddr ? io_avail_list_17 : _GEN_592; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_594 = 6'h12 == buf_4_rs2_paddr ? io_avail_list_18 : _GEN_593; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_595 = 6'h13 == buf_4_rs2_paddr ? io_avail_list_19 : _GEN_594; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_596 = 6'h14 == buf_4_rs2_paddr ? io_avail_list_20 : _GEN_595; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_597 = 6'h15 == buf_4_rs2_paddr ? io_avail_list_21 : _GEN_596; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_598 = 6'h16 == buf_4_rs2_paddr ? io_avail_list_22 : _GEN_597; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_599 = 6'h17 == buf_4_rs2_paddr ? io_avail_list_23 : _GEN_598; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_600 = 6'h18 == buf_4_rs2_paddr ? io_avail_list_24 : _GEN_599; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_601 = 6'h19 == buf_4_rs2_paddr ? io_avail_list_25 : _GEN_600; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_602 = 6'h1a == buf_4_rs2_paddr ? io_avail_list_26 : _GEN_601; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_603 = 6'h1b == buf_4_rs2_paddr ? io_avail_list_27 : _GEN_602; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_604 = 6'h1c == buf_4_rs2_paddr ? io_avail_list_28 : _GEN_603; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_605 = 6'h1d == buf_4_rs2_paddr ? io_avail_list_29 : _GEN_604; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_606 = 6'h1e == buf_4_rs2_paddr ? io_avail_list_30 : _GEN_605; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_607 = 6'h1f == buf_4_rs2_paddr ? io_avail_list_31 : _GEN_606; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_608 = 6'h20 == buf_4_rs2_paddr ? io_avail_list_32 : _GEN_607; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_609 = 6'h21 == buf_4_rs2_paddr ? io_avail_list_33 : _GEN_608; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_610 = 6'h22 == buf_4_rs2_paddr ? io_avail_list_34 : _GEN_609; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_611 = 6'h23 == buf_4_rs2_paddr ? io_avail_list_35 : _GEN_610; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_612 = 6'h24 == buf_4_rs2_paddr ? io_avail_list_36 : _GEN_611; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_613 = 6'h25 == buf_4_rs2_paddr ? io_avail_list_37 : _GEN_612; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_614 = 6'h26 == buf_4_rs2_paddr ? io_avail_list_38 : _GEN_613; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_615 = 6'h27 == buf_4_rs2_paddr ? io_avail_list_39 : _GEN_614; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_616 = 6'h28 == buf_4_rs2_paddr ? io_avail_list_40 : _GEN_615; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_617 = 6'h29 == buf_4_rs2_paddr ? io_avail_list_41 : _GEN_616; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_618 = 6'h2a == buf_4_rs2_paddr ? io_avail_list_42 : _GEN_617; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_619 = 6'h2b == buf_4_rs2_paddr ? io_avail_list_43 : _GEN_618; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_620 = 6'h2c == buf_4_rs2_paddr ? io_avail_list_44 : _GEN_619; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_621 = 6'h2d == buf_4_rs2_paddr ? io_avail_list_45 : _GEN_620; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_622 = 6'h2e == buf_4_rs2_paddr ? io_avail_list_46 : _GEN_621; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_623 = 6'h2f == buf_4_rs2_paddr ? io_avail_list_47 : _GEN_622; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_624 = 6'h30 == buf_4_rs2_paddr ? io_avail_list_48 : _GEN_623; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_625 = 6'h31 == buf_4_rs2_paddr ? io_avail_list_49 : _GEN_624; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_626 = 6'h32 == buf_4_rs2_paddr ? io_avail_list_50 : _GEN_625; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_627 = 6'h33 == buf_4_rs2_paddr ? io_avail_list_51 : _GEN_626; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_628 = 6'h34 == buf_4_rs2_paddr ? io_avail_list_52 : _GEN_627; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_629 = 6'h35 == buf_4_rs2_paddr ? io_avail_list_53 : _GEN_628; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_630 = 6'h36 == buf_4_rs2_paddr ? io_avail_list_54 : _GEN_629; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_631 = 6'h37 == buf_4_rs2_paddr ? io_avail_list_55 : _GEN_630; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_632 = 6'h38 == buf_4_rs2_paddr ? io_avail_list_56 : _GEN_631; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_633 = 6'h39 == buf_4_rs2_paddr ? io_avail_list_57 : _GEN_632; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_634 = 6'h3a == buf_4_rs2_paddr ? io_avail_list_58 : _GEN_633; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_635 = 6'h3b == buf_4_rs2_paddr ? io_avail_list_59 : _GEN_634; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_636 = 6'h3c == buf_4_rs2_paddr ? io_avail_list_60 : _GEN_635; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_637 = 6'h3d == buf_4_rs2_paddr ? io_avail_list_61 : _GEN_636; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_638 = 6'h3e == buf_4_rs2_paddr ? io_avail_list_62 : _GEN_637; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_639 = 6'h3f == buf_4_rs2_paddr ? io_avail_list_63 : _GEN_638; // @[IssueUnit.scala 268:{32,32}]
  wire  ready_list_4 = _GEN_575 & _GEN_639 & io_fu_ready & store_mask_4; // @[IssueUnit.scala 268:57]
  wire  _GEN_641 = 6'h1 == buf_5_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_642 = 6'h2 == buf_5_rs1_paddr ? io_avail_list_2 : _GEN_641; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_643 = 6'h3 == buf_5_rs1_paddr ? io_avail_list_3 : _GEN_642; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_644 = 6'h4 == buf_5_rs1_paddr ? io_avail_list_4 : _GEN_643; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_645 = 6'h5 == buf_5_rs1_paddr ? io_avail_list_5 : _GEN_644; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_646 = 6'h6 == buf_5_rs1_paddr ? io_avail_list_6 : _GEN_645; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_647 = 6'h7 == buf_5_rs1_paddr ? io_avail_list_7 : _GEN_646; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_648 = 6'h8 == buf_5_rs1_paddr ? io_avail_list_8 : _GEN_647; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_649 = 6'h9 == buf_5_rs1_paddr ? io_avail_list_9 : _GEN_648; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_650 = 6'ha == buf_5_rs1_paddr ? io_avail_list_10 : _GEN_649; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_651 = 6'hb == buf_5_rs1_paddr ? io_avail_list_11 : _GEN_650; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_652 = 6'hc == buf_5_rs1_paddr ? io_avail_list_12 : _GEN_651; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_653 = 6'hd == buf_5_rs1_paddr ? io_avail_list_13 : _GEN_652; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_654 = 6'he == buf_5_rs1_paddr ? io_avail_list_14 : _GEN_653; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_655 = 6'hf == buf_5_rs1_paddr ? io_avail_list_15 : _GEN_654; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_656 = 6'h10 == buf_5_rs1_paddr ? io_avail_list_16 : _GEN_655; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_657 = 6'h11 == buf_5_rs1_paddr ? io_avail_list_17 : _GEN_656; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_658 = 6'h12 == buf_5_rs1_paddr ? io_avail_list_18 : _GEN_657; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_659 = 6'h13 == buf_5_rs1_paddr ? io_avail_list_19 : _GEN_658; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_660 = 6'h14 == buf_5_rs1_paddr ? io_avail_list_20 : _GEN_659; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_661 = 6'h15 == buf_5_rs1_paddr ? io_avail_list_21 : _GEN_660; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_662 = 6'h16 == buf_5_rs1_paddr ? io_avail_list_22 : _GEN_661; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_663 = 6'h17 == buf_5_rs1_paddr ? io_avail_list_23 : _GEN_662; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_664 = 6'h18 == buf_5_rs1_paddr ? io_avail_list_24 : _GEN_663; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_665 = 6'h19 == buf_5_rs1_paddr ? io_avail_list_25 : _GEN_664; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_666 = 6'h1a == buf_5_rs1_paddr ? io_avail_list_26 : _GEN_665; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_667 = 6'h1b == buf_5_rs1_paddr ? io_avail_list_27 : _GEN_666; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_668 = 6'h1c == buf_5_rs1_paddr ? io_avail_list_28 : _GEN_667; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_669 = 6'h1d == buf_5_rs1_paddr ? io_avail_list_29 : _GEN_668; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_670 = 6'h1e == buf_5_rs1_paddr ? io_avail_list_30 : _GEN_669; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_671 = 6'h1f == buf_5_rs1_paddr ? io_avail_list_31 : _GEN_670; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_672 = 6'h20 == buf_5_rs1_paddr ? io_avail_list_32 : _GEN_671; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_673 = 6'h21 == buf_5_rs1_paddr ? io_avail_list_33 : _GEN_672; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_674 = 6'h22 == buf_5_rs1_paddr ? io_avail_list_34 : _GEN_673; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_675 = 6'h23 == buf_5_rs1_paddr ? io_avail_list_35 : _GEN_674; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_676 = 6'h24 == buf_5_rs1_paddr ? io_avail_list_36 : _GEN_675; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_677 = 6'h25 == buf_5_rs1_paddr ? io_avail_list_37 : _GEN_676; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_678 = 6'h26 == buf_5_rs1_paddr ? io_avail_list_38 : _GEN_677; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_679 = 6'h27 == buf_5_rs1_paddr ? io_avail_list_39 : _GEN_678; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_680 = 6'h28 == buf_5_rs1_paddr ? io_avail_list_40 : _GEN_679; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_681 = 6'h29 == buf_5_rs1_paddr ? io_avail_list_41 : _GEN_680; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_682 = 6'h2a == buf_5_rs1_paddr ? io_avail_list_42 : _GEN_681; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_683 = 6'h2b == buf_5_rs1_paddr ? io_avail_list_43 : _GEN_682; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_684 = 6'h2c == buf_5_rs1_paddr ? io_avail_list_44 : _GEN_683; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_685 = 6'h2d == buf_5_rs1_paddr ? io_avail_list_45 : _GEN_684; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_686 = 6'h2e == buf_5_rs1_paddr ? io_avail_list_46 : _GEN_685; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_687 = 6'h2f == buf_5_rs1_paddr ? io_avail_list_47 : _GEN_686; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_688 = 6'h30 == buf_5_rs1_paddr ? io_avail_list_48 : _GEN_687; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_689 = 6'h31 == buf_5_rs1_paddr ? io_avail_list_49 : _GEN_688; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_690 = 6'h32 == buf_5_rs1_paddr ? io_avail_list_50 : _GEN_689; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_691 = 6'h33 == buf_5_rs1_paddr ? io_avail_list_51 : _GEN_690; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_692 = 6'h34 == buf_5_rs1_paddr ? io_avail_list_52 : _GEN_691; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_693 = 6'h35 == buf_5_rs1_paddr ? io_avail_list_53 : _GEN_692; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_694 = 6'h36 == buf_5_rs1_paddr ? io_avail_list_54 : _GEN_693; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_695 = 6'h37 == buf_5_rs1_paddr ? io_avail_list_55 : _GEN_694; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_696 = 6'h38 == buf_5_rs1_paddr ? io_avail_list_56 : _GEN_695; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_697 = 6'h39 == buf_5_rs1_paddr ? io_avail_list_57 : _GEN_696; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_698 = 6'h3a == buf_5_rs1_paddr ? io_avail_list_58 : _GEN_697; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_699 = 6'h3b == buf_5_rs1_paddr ? io_avail_list_59 : _GEN_698; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_700 = 6'h3c == buf_5_rs1_paddr ? io_avail_list_60 : _GEN_699; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_701 = 6'h3d == buf_5_rs1_paddr ? io_avail_list_61 : _GEN_700; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_702 = 6'h3e == buf_5_rs1_paddr ? io_avail_list_62 : _GEN_701; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_703 = 6'h3f == buf_5_rs1_paddr ? io_avail_list_63 : _GEN_702; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_705 = 6'h1 == buf_5_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_706 = 6'h2 == buf_5_rs2_paddr ? io_avail_list_2 : _GEN_705; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_707 = 6'h3 == buf_5_rs2_paddr ? io_avail_list_3 : _GEN_706; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_708 = 6'h4 == buf_5_rs2_paddr ? io_avail_list_4 : _GEN_707; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_709 = 6'h5 == buf_5_rs2_paddr ? io_avail_list_5 : _GEN_708; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_710 = 6'h6 == buf_5_rs2_paddr ? io_avail_list_6 : _GEN_709; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_711 = 6'h7 == buf_5_rs2_paddr ? io_avail_list_7 : _GEN_710; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_712 = 6'h8 == buf_5_rs2_paddr ? io_avail_list_8 : _GEN_711; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_713 = 6'h9 == buf_5_rs2_paddr ? io_avail_list_9 : _GEN_712; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_714 = 6'ha == buf_5_rs2_paddr ? io_avail_list_10 : _GEN_713; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_715 = 6'hb == buf_5_rs2_paddr ? io_avail_list_11 : _GEN_714; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_716 = 6'hc == buf_5_rs2_paddr ? io_avail_list_12 : _GEN_715; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_717 = 6'hd == buf_5_rs2_paddr ? io_avail_list_13 : _GEN_716; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_718 = 6'he == buf_5_rs2_paddr ? io_avail_list_14 : _GEN_717; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_719 = 6'hf == buf_5_rs2_paddr ? io_avail_list_15 : _GEN_718; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_720 = 6'h10 == buf_5_rs2_paddr ? io_avail_list_16 : _GEN_719; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_721 = 6'h11 == buf_5_rs2_paddr ? io_avail_list_17 : _GEN_720; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_722 = 6'h12 == buf_5_rs2_paddr ? io_avail_list_18 : _GEN_721; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_723 = 6'h13 == buf_5_rs2_paddr ? io_avail_list_19 : _GEN_722; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_724 = 6'h14 == buf_5_rs2_paddr ? io_avail_list_20 : _GEN_723; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_725 = 6'h15 == buf_5_rs2_paddr ? io_avail_list_21 : _GEN_724; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_726 = 6'h16 == buf_5_rs2_paddr ? io_avail_list_22 : _GEN_725; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_727 = 6'h17 == buf_5_rs2_paddr ? io_avail_list_23 : _GEN_726; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_728 = 6'h18 == buf_5_rs2_paddr ? io_avail_list_24 : _GEN_727; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_729 = 6'h19 == buf_5_rs2_paddr ? io_avail_list_25 : _GEN_728; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_730 = 6'h1a == buf_5_rs2_paddr ? io_avail_list_26 : _GEN_729; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_731 = 6'h1b == buf_5_rs2_paddr ? io_avail_list_27 : _GEN_730; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_732 = 6'h1c == buf_5_rs2_paddr ? io_avail_list_28 : _GEN_731; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_733 = 6'h1d == buf_5_rs2_paddr ? io_avail_list_29 : _GEN_732; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_734 = 6'h1e == buf_5_rs2_paddr ? io_avail_list_30 : _GEN_733; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_735 = 6'h1f == buf_5_rs2_paddr ? io_avail_list_31 : _GEN_734; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_736 = 6'h20 == buf_5_rs2_paddr ? io_avail_list_32 : _GEN_735; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_737 = 6'h21 == buf_5_rs2_paddr ? io_avail_list_33 : _GEN_736; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_738 = 6'h22 == buf_5_rs2_paddr ? io_avail_list_34 : _GEN_737; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_739 = 6'h23 == buf_5_rs2_paddr ? io_avail_list_35 : _GEN_738; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_740 = 6'h24 == buf_5_rs2_paddr ? io_avail_list_36 : _GEN_739; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_741 = 6'h25 == buf_5_rs2_paddr ? io_avail_list_37 : _GEN_740; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_742 = 6'h26 == buf_5_rs2_paddr ? io_avail_list_38 : _GEN_741; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_743 = 6'h27 == buf_5_rs2_paddr ? io_avail_list_39 : _GEN_742; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_744 = 6'h28 == buf_5_rs2_paddr ? io_avail_list_40 : _GEN_743; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_745 = 6'h29 == buf_5_rs2_paddr ? io_avail_list_41 : _GEN_744; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_746 = 6'h2a == buf_5_rs2_paddr ? io_avail_list_42 : _GEN_745; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_747 = 6'h2b == buf_5_rs2_paddr ? io_avail_list_43 : _GEN_746; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_748 = 6'h2c == buf_5_rs2_paddr ? io_avail_list_44 : _GEN_747; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_749 = 6'h2d == buf_5_rs2_paddr ? io_avail_list_45 : _GEN_748; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_750 = 6'h2e == buf_5_rs2_paddr ? io_avail_list_46 : _GEN_749; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_751 = 6'h2f == buf_5_rs2_paddr ? io_avail_list_47 : _GEN_750; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_752 = 6'h30 == buf_5_rs2_paddr ? io_avail_list_48 : _GEN_751; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_753 = 6'h31 == buf_5_rs2_paddr ? io_avail_list_49 : _GEN_752; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_754 = 6'h32 == buf_5_rs2_paddr ? io_avail_list_50 : _GEN_753; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_755 = 6'h33 == buf_5_rs2_paddr ? io_avail_list_51 : _GEN_754; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_756 = 6'h34 == buf_5_rs2_paddr ? io_avail_list_52 : _GEN_755; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_757 = 6'h35 == buf_5_rs2_paddr ? io_avail_list_53 : _GEN_756; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_758 = 6'h36 == buf_5_rs2_paddr ? io_avail_list_54 : _GEN_757; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_759 = 6'h37 == buf_5_rs2_paddr ? io_avail_list_55 : _GEN_758; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_760 = 6'h38 == buf_5_rs2_paddr ? io_avail_list_56 : _GEN_759; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_761 = 6'h39 == buf_5_rs2_paddr ? io_avail_list_57 : _GEN_760; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_762 = 6'h3a == buf_5_rs2_paddr ? io_avail_list_58 : _GEN_761; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_763 = 6'h3b == buf_5_rs2_paddr ? io_avail_list_59 : _GEN_762; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_764 = 6'h3c == buf_5_rs2_paddr ? io_avail_list_60 : _GEN_763; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_765 = 6'h3d == buf_5_rs2_paddr ? io_avail_list_61 : _GEN_764; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_766 = 6'h3e == buf_5_rs2_paddr ? io_avail_list_62 : _GEN_765; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_767 = 6'h3f == buf_5_rs2_paddr ? io_avail_list_63 : _GEN_766; // @[IssueUnit.scala 268:{32,32}]
  wire  ready_list_5 = _GEN_703 & _GEN_767 & io_fu_ready & store_mask_5; // @[IssueUnit.scala 268:57]
  wire  _GEN_769 = 6'h1 == buf_6_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_770 = 6'h2 == buf_6_rs1_paddr ? io_avail_list_2 : _GEN_769; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_771 = 6'h3 == buf_6_rs1_paddr ? io_avail_list_3 : _GEN_770; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_772 = 6'h4 == buf_6_rs1_paddr ? io_avail_list_4 : _GEN_771; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_773 = 6'h5 == buf_6_rs1_paddr ? io_avail_list_5 : _GEN_772; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_774 = 6'h6 == buf_6_rs1_paddr ? io_avail_list_6 : _GEN_773; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_775 = 6'h7 == buf_6_rs1_paddr ? io_avail_list_7 : _GEN_774; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_776 = 6'h8 == buf_6_rs1_paddr ? io_avail_list_8 : _GEN_775; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_777 = 6'h9 == buf_6_rs1_paddr ? io_avail_list_9 : _GEN_776; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_778 = 6'ha == buf_6_rs1_paddr ? io_avail_list_10 : _GEN_777; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_779 = 6'hb == buf_6_rs1_paddr ? io_avail_list_11 : _GEN_778; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_780 = 6'hc == buf_6_rs1_paddr ? io_avail_list_12 : _GEN_779; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_781 = 6'hd == buf_6_rs1_paddr ? io_avail_list_13 : _GEN_780; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_782 = 6'he == buf_6_rs1_paddr ? io_avail_list_14 : _GEN_781; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_783 = 6'hf == buf_6_rs1_paddr ? io_avail_list_15 : _GEN_782; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_784 = 6'h10 == buf_6_rs1_paddr ? io_avail_list_16 : _GEN_783; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_785 = 6'h11 == buf_6_rs1_paddr ? io_avail_list_17 : _GEN_784; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_786 = 6'h12 == buf_6_rs1_paddr ? io_avail_list_18 : _GEN_785; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_787 = 6'h13 == buf_6_rs1_paddr ? io_avail_list_19 : _GEN_786; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_788 = 6'h14 == buf_6_rs1_paddr ? io_avail_list_20 : _GEN_787; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_789 = 6'h15 == buf_6_rs1_paddr ? io_avail_list_21 : _GEN_788; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_790 = 6'h16 == buf_6_rs1_paddr ? io_avail_list_22 : _GEN_789; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_791 = 6'h17 == buf_6_rs1_paddr ? io_avail_list_23 : _GEN_790; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_792 = 6'h18 == buf_6_rs1_paddr ? io_avail_list_24 : _GEN_791; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_793 = 6'h19 == buf_6_rs1_paddr ? io_avail_list_25 : _GEN_792; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_794 = 6'h1a == buf_6_rs1_paddr ? io_avail_list_26 : _GEN_793; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_795 = 6'h1b == buf_6_rs1_paddr ? io_avail_list_27 : _GEN_794; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_796 = 6'h1c == buf_6_rs1_paddr ? io_avail_list_28 : _GEN_795; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_797 = 6'h1d == buf_6_rs1_paddr ? io_avail_list_29 : _GEN_796; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_798 = 6'h1e == buf_6_rs1_paddr ? io_avail_list_30 : _GEN_797; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_799 = 6'h1f == buf_6_rs1_paddr ? io_avail_list_31 : _GEN_798; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_800 = 6'h20 == buf_6_rs1_paddr ? io_avail_list_32 : _GEN_799; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_801 = 6'h21 == buf_6_rs1_paddr ? io_avail_list_33 : _GEN_800; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_802 = 6'h22 == buf_6_rs1_paddr ? io_avail_list_34 : _GEN_801; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_803 = 6'h23 == buf_6_rs1_paddr ? io_avail_list_35 : _GEN_802; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_804 = 6'h24 == buf_6_rs1_paddr ? io_avail_list_36 : _GEN_803; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_805 = 6'h25 == buf_6_rs1_paddr ? io_avail_list_37 : _GEN_804; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_806 = 6'h26 == buf_6_rs1_paddr ? io_avail_list_38 : _GEN_805; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_807 = 6'h27 == buf_6_rs1_paddr ? io_avail_list_39 : _GEN_806; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_808 = 6'h28 == buf_6_rs1_paddr ? io_avail_list_40 : _GEN_807; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_809 = 6'h29 == buf_6_rs1_paddr ? io_avail_list_41 : _GEN_808; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_810 = 6'h2a == buf_6_rs1_paddr ? io_avail_list_42 : _GEN_809; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_811 = 6'h2b == buf_6_rs1_paddr ? io_avail_list_43 : _GEN_810; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_812 = 6'h2c == buf_6_rs1_paddr ? io_avail_list_44 : _GEN_811; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_813 = 6'h2d == buf_6_rs1_paddr ? io_avail_list_45 : _GEN_812; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_814 = 6'h2e == buf_6_rs1_paddr ? io_avail_list_46 : _GEN_813; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_815 = 6'h2f == buf_6_rs1_paddr ? io_avail_list_47 : _GEN_814; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_816 = 6'h30 == buf_6_rs1_paddr ? io_avail_list_48 : _GEN_815; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_817 = 6'h31 == buf_6_rs1_paddr ? io_avail_list_49 : _GEN_816; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_818 = 6'h32 == buf_6_rs1_paddr ? io_avail_list_50 : _GEN_817; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_819 = 6'h33 == buf_6_rs1_paddr ? io_avail_list_51 : _GEN_818; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_820 = 6'h34 == buf_6_rs1_paddr ? io_avail_list_52 : _GEN_819; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_821 = 6'h35 == buf_6_rs1_paddr ? io_avail_list_53 : _GEN_820; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_822 = 6'h36 == buf_6_rs1_paddr ? io_avail_list_54 : _GEN_821; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_823 = 6'h37 == buf_6_rs1_paddr ? io_avail_list_55 : _GEN_822; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_824 = 6'h38 == buf_6_rs1_paddr ? io_avail_list_56 : _GEN_823; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_825 = 6'h39 == buf_6_rs1_paddr ? io_avail_list_57 : _GEN_824; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_826 = 6'h3a == buf_6_rs1_paddr ? io_avail_list_58 : _GEN_825; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_827 = 6'h3b == buf_6_rs1_paddr ? io_avail_list_59 : _GEN_826; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_828 = 6'h3c == buf_6_rs1_paddr ? io_avail_list_60 : _GEN_827; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_829 = 6'h3d == buf_6_rs1_paddr ? io_avail_list_61 : _GEN_828; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_830 = 6'h3e == buf_6_rs1_paddr ? io_avail_list_62 : _GEN_829; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_831 = 6'h3f == buf_6_rs1_paddr ? io_avail_list_63 : _GEN_830; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_833 = 6'h1 == buf_6_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_834 = 6'h2 == buf_6_rs2_paddr ? io_avail_list_2 : _GEN_833; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_835 = 6'h3 == buf_6_rs2_paddr ? io_avail_list_3 : _GEN_834; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_836 = 6'h4 == buf_6_rs2_paddr ? io_avail_list_4 : _GEN_835; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_837 = 6'h5 == buf_6_rs2_paddr ? io_avail_list_5 : _GEN_836; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_838 = 6'h6 == buf_6_rs2_paddr ? io_avail_list_6 : _GEN_837; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_839 = 6'h7 == buf_6_rs2_paddr ? io_avail_list_7 : _GEN_838; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_840 = 6'h8 == buf_6_rs2_paddr ? io_avail_list_8 : _GEN_839; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_841 = 6'h9 == buf_6_rs2_paddr ? io_avail_list_9 : _GEN_840; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_842 = 6'ha == buf_6_rs2_paddr ? io_avail_list_10 : _GEN_841; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_843 = 6'hb == buf_6_rs2_paddr ? io_avail_list_11 : _GEN_842; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_844 = 6'hc == buf_6_rs2_paddr ? io_avail_list_12 : _GEN_843; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_845 = 6'hd == buf_6_rs2_paddr ? io_avail_list_13 : _GEN_844; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_846 = 6'he == buf_6_rs2_paddr ? io_avail_list_14 : _GEN_845; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_847 = 6'hf == buf_6_rs2_paddr ? io_avail_list_15 : _GEN_846; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_848 = 6'h10 == buf_6_rs2_paddr ? io_avail_list_16 : _GEN_847; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_849 = 6'h11 == buf_6_rs2_paddr ? io_avail_list_17 : _GEN_848; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_850 = 6'h12 == buf_6_rs2_paddr ? io_avail_list_18 : _GEN_849; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_851 = 6'h13 == buf_6_rs2_paddr ? io_avail_list_19 : _GEN_850; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_852 = 6'h14 == buf_6_rs2_paddr ? io_avail_list_20 : _GEN_851; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_853 = 6'h15 == buf_6_rs2_paddr ? io_avail_list_21 : _GEN_852; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_854 = 6'h16 == buf_6_rs2_paddr ? io_avail_list_22 : _GEN_853; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_855 = 6'h17 == buf_6_rs2_paddr ? io_avail_list_23 : _GEN_854; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_856 = 6'h18 == buf_6_rs2_paddr ? io_avail_list_24 : _GEN_855; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_857 = 6'h19 == buf_6_rs2_paddr ? io_avail_list_25 : _GEN_856; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_858 = 6'h1a == buf_6_rs2_paddr ? io_avail_list_26 : _GEN_857; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_859 = 6'h1b == buf_6_rs2_paddr ? io_avail_list_27 : _GEN_858; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_860 = 6'h1c == buf_6_rs2_paddr ? io_avail_list_28 : _GEN_859; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_861 = 6'h1d == buf_6_rs2_paddr ? io_avail_list_29 : _GEN_860; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_862 = 6'h1e == buf_6_rs2_paddr ? io_avail_list_30 : _GEN_861; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_863 = 6'h1f == buf_6_rs2_paddr ? io_avail_list_31 : _GEN_862; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_864 = 6'h20 == buf_6_rs2_paddr ? io_avail_list_32 : _GEN_863; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_865 = 6'h21 == buf_6_rs2_paddr ? io_avail_list_33 : _GEN_864; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_866 = 6'h22 == buf_6_rs2_paddr ? io_avail_list_34 : _GEN_865; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_867 = 6'h23 == buf_6_rs2_paddr ? io_avail_list_35 : _GEN_866; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_868 = 6'h24 == buf_6_rs2_paddr ? io_avail_list_36 : _GEN_867; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_869 = 6'h25 == buf_6_rs2_paddr ? io_avail_list_37 : _GEN_868; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_870 = 6'h26 == buf_6_rs2_paddr ? io_avail_list_38 : _GEN_869; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_871 = 6'h27 == buf_6_rs2_paddr ? io_avail_list_39 : _GEN_870; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_872 = 6'h28 == buf_6_rs2_paddr ? io_avail_list_40 : _GEN_871; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_873 = 6'h29 == buf_6_rs2_paddr ? io_avail_list_41 : _GEN_872; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_874 = 6'h2a == buf_6_rs2_paddr ? io_avail_list_42 : _GEN_873; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_875 = 6'h2b == buf_6_rs2_paddr ? io_avail_list_43 : _GEN_874; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_876 = 6'h2c == buf_6_rs2_paddr ? io_avail_list_44 : _GEN_875; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_877 = 6'h2d == buf_6_rs2_paddr ? io_avail_list_45 : _GEN_876; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_878 = 6'h2e == buf_6_rs2_paddr ? io_avail_list_46 : _GEN_877; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_879 = 6'h2f == buf_6_rs2_paddr ? io_avail_list_47 : _GEN_878; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_880 = 6'h30 == buf_6_rs2_paddr ? io_avail_list_48 : _GEN_879; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_881 = 6'h31 == buf_6_rs2_paddr ? io_avail_list_49 : _GEN_880; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_882 = 6'h32 == buf_6_rs2_paddr ? io_avail_list_50 : _GEN_881; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_883 = 6'h33 == buf_6_rs2_paddr ? io_avail_list_51 : _GEN_882; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_884 = 6'h34 == buf_6_rs2_paddr ? io_avail_list_52 : _GEN_883; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_885 = 6'h35 == buf_6_rs2_paddr ? io_avail_list_53 : _GEN_884; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_886 = 6'h36 == buf_6_rs2_paddr ? io_avail_list_54 : _GEN_885; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_887 = 6'h37 == buf_6_rs2_paddr ? io_avail_list_55 : _GEN_886; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_888 = 6'h38 == buf_6_rs2_paddr ? io_avail_list_56 : _GEN_887; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_889 = 6'h39 == buf_6_rs2_paddr ? io_avail_list_57 : _GEN_888; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_890 = 6'h3a == buf_6_rs2_paddr ? io_avail_list_58 : _GEN_889; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_891 = 6'h3b == buf_6_rs2_paddr ? io_avail_list_59 : _GEN_890; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_892 = 6'h3c == buf_6_rs2_paddr ? io_avail_list_60 : _GEN_891; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_893 = 6'h3d == buf_6_rs2_paddr ? io_avail_list_61 : _GEN_892; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_894 = 6'h3e == buf_6_rs2_paddr ? io_avail_list_62 : _GEN_893; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_895 = 6'h3f == buf_6_rs2_paddr ? io_avail_list_63 : _GEN_894; // @[IssueUnit.scala 268:{32,32}]
  wire  ready_list_6 = _GEN_831 & _GEN_895 & io_fu_ready & store_mask_6; // @[IssueUnit.scala 268:57]
  wire  _GEN_897 = 6'h1 == buf_7_rs1_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_898 = 6'h2 == buf_7_rs1_paddr ? io_avail_list_2 : _GEN_897; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_899 = 6'h3 == buf_7_rs1_paddr ? io_avail_list_3 : _GEN_898; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_900 = 6'h4 == buf_7_rs1_paddr ? io_avail_list_4 : _GEN_899; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_901 = 6'h5 == buf_7_rs1_paddr ? io_avail_list_5 : _GEN_900; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_902 = 6'h6 == buf_7_rs1_paddr ? io_avail_list_6 : _GEN_901; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_903 = 6'h7 == buf_7_rs1_paddr ? io_avail_list_7 : _GEN_902; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_904 = 6'h8 == buf_7_rs1_paddr ? io_avail_list_8 : _GEN_903; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_905 = 6'h9 == buf_7_rs1_paddr ? io_avail_list_9 : _GEN_904; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_906 = 6'ha == buf_7_rs1_paddr ? io_avail_list_10 : _GEN_905; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_907 = 6'hb == buf_7_rs1_paddr ? io_avail_list_11 : _GEN_906; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_908 = 6'hc == buf_7_rs1_paddr ? io_avail_list_12 : _GEN_907; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_909 = 6'hd == buf_7_rs1_paddr ? io_avail_list_13 : _GEN_908; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_910 = 6'he == buf_7_rs1_paddr ? io_avail_list_14 : _GEN_909; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_911 = 6'hf == buf_7_rs1_paddr ? io_avail_list_15 : _GEN_910; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_912 = 6'h10 == buf_7_rs1_paddr ? io_avail_list_16 : _GEN_911; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_913 = 6'h11 == buf_7_rs1_paddr ? io_avail_list_17 : _GEN_912; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_914 = 6'h12 == buf_7_rs1_paddr ? io_avail_list_18 : _GEN_913; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_915 = 6'h13 == buf_7_rs1_paddr ? io_avail_list_19 : _GEN_914; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_916 = 6'h14 == buf_7_rs1_paddr ? io_avail_list_20 : _GEN_915; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_917 = 6'h15 == buf_7_rs1_paddr ? io_avail_list_21 : _GEN_916; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_918 = 6'h16 == buf_7_rs1_paddr ? io_avail_list_22 : _GEN_917; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_919 = 6'h17 == buf_7_rs1_paddr ? io_avail_list_23 : _GEN_918; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_920 = 6'h18 == buf_7_rs1_paddr ? io_avail_list_24 : _GEN_919; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_921 = 6'h19 == buf_7_rs1_paddr ? io_avail_list_25 : _GEN_920; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_922 = 6'h1a == buf_7_rs1_paddr ? io_avail_list_26 : _GEN_921; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_923 = 6'h1b == buf_7_rs1_paddr ? io_avail_list_27 : _GEN_922; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_924 = 6'h1c == buf_7_rs1_paddr ? io_avail_list_28 : _GEN_923; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_925 = 6'h1d == buf_7_rs1_paddr ? io_avail_list_29 : _GEN_924; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_926 = 6'h1e == buf_7_rs1_paddr ? io_avail_list_30 : _GEN_925; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_927 = 6'h1f == buf_7_rs1_paddr ? io_avail_list_31 : _GEN_926; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_928 = 6'h20 == buf_7_rs1_paddr ? io_avail_list_32 : _GEN_927; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_929 = 6'h21 == buf_7_rs1_paddr ? io_avail_list_33 : _GEN_928; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_930 = 6'h22 == buf_7_rs1_paddr ? io_avail_list_34 : _GEN_929; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_931 = 6'h23 == buf_7_rs1_paddr ? io_avail_list_35 : _GEN_930; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_932 = 6'h24 == buf_7_rs1_paddr ? io_avail_list_36 : _GEN_931; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_933 = 6'h25 == buf_7_rs1_paddr ? io_avail_list_37 : _GEN_932; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_934 = 6'h26 == buf_7_rs1_paddr ? io_avail_list_38 : _GEN_933; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_935 = 6'h27 == buf_7_rs1_paddr ? io_avail_list_39 : _GEN_934; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_936 = 6'h28 == buf_7_rs1_paddr ? io_avail_list_40 : _GEN_935; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_937 = 6'h29 == buf_7_rs1_paddr ? io_avail_list_41 : _GEN_936; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_938 = 6'h2a == buf_7_rs1_paddr ? io_avail_list_42 : _GEN_937; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_939 = 6'h2b == buf_7_rs1_paddr ? io_avail_list_43 : _GEN_938; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_940 = 6'h2c == buf_7_rs1_paddr ? io_avail_list_44 : _GEN_939; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_941 = 6'h2d == buf_7_rs1_paddr ? io_avail_list_45 : _GEN_940; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_942 = 6'h2e == buf_7_rs1_paddr ? io_avail_list_46 : _GEN_941; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_943 = 6'h2f == buf_7_rs1_paddr ? io_avail_list_47 : _GEN_942; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_944 = 6'h30 == buf_7_rs1_paddr ? io_avail_list_48 : _GEN_943; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_945 = 6'h31 == buf_7_rs1_paddr ? io_avail_list_49 : _GEN_944; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_946 = 6'h32 == buf_7_rs1_paddr ? io_avail_list_50 : _GEN_945; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_947 = 6'h33 == buf_7_rs1_paddr ? io_avail_list_51 : _GEN_946; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_948 = 6'h34 == buf_7_rs1_paddr ? io_avail_list_52 : _GEN_947; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_949 = 6'h35 == buf_7_rs1_paddr ? io_avail_list_53 : _GEN_948; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_950 = 6'h36 == buf_7_rs1_paddr ? io_avail_list_54 : _GEN_949; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_951 = 6'h37 == buf_7_rs1_paddr ? io_avail_list_55 : _GEN_950; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_952 = 6'h38 == buf_7_rs1_paddr ? io_avail_list_56 : _GEN_951; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_953 = 6'h39 == buf_7_rs1_paddr ? io_avail_list_57 : _GEN_952; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_954 = 6'h3a == buf_7_rs1_paddr ? io_avail_list_58 : _GEN_953; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_955 = 6'h3b == buf_7_rs1_paddr ? io_avail_list_59 : _GEN_954; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_956 = 6'h3c == buf_7_rs1_paddr ? io_avail_list_60 : _GEN_955; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_957 = 6'h3d == buf_7_rs1_paddr ? io_avail_list_61 : _GEN_956; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_958 = 6'h3e == buf_7_rs1_paddr ? io_avail_list_62 : _GEN_957; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_959 = 6'h3f == buf_7_rs1_paddr ? io_avail_list_63 : _GEN_958; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_961 = 6'h1 == buf_7_rs2_paddr ? io_avail_list_1 : io_avail_list_0; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_962 = 6'h2 == buf_7_rs2_paddr ? io_avail_list_2 : _GEN_961; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_963 = 6'h3 == buf_7_rs2_paddr ? io_avail_list_3 : _GEN_962; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_964 = 6'h4 == buf_7_rs2_paddr ? io_avail_list_4 : _GEN_963; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_965 = 6'h5 == buf_7_rs2_paddr ? io_avail_list_5 : _GEN_964; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_966 = 6'h6 == buf_7_rs2_paddr ? io_avail_list_6 : _GEN_965; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_967 = 6'h7 == buf_7_rs2_paddr ? io_avail_list_7 : _GEN_966; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_968 = 6'h8 == buf_7_rs2_paddr ? io_avail_list_8 : _GEN_967; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_969 = 6'h9 == buf_7_rs2_paddr ? io_avail_list_9 : _GEN_968; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_970 = 6'ha == buf_7_rs2_paddr ? io_avail_list_10 : _GEN_969; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_971 = 6'hb == buf_7_rs2_paddr ? io_avail_list_11 : _GEN_970; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_972 = 6'hc == buf_7_rs2_paddr ? io_avail_list_12 : _GEN_971; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_973 = 6'hd == buf_7_rs2_paddr ? io_avail_list_13 : _GEN_972; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_974 = 6'he == buf_7_rs2_paddr ? io_avail_list_14 : _GEN_973; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_975 = 6'hf == buf_7_rs2_paddr ? io_avail_list_15 : _GEN_974; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_976 = 6'h10 == buf_7_rs2_paddr ? io_avail_list_16 : _GEN_975; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_977 = 6'h11 == buf_7_rs2_paddr ? io_avail_list_17 : _GEN_976; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_978 = 6'h12 == buf_7_rs2_paddr ? io_avail_list_18 : _GEN_977; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_979 = 6'h13 == buf_7_rs2_paddr ? io_avail_list_19 : _GEN_978; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_980 = 6'h14 == buf_7_rs2_paddr ? io_avail_list_20 : _GEN_979; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_981 = 6'h15 == buf_7_rs2_paddr ? io_avail_list_21 : _GEN_980; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_982 = 6'h16 == buf_7_rs2_paddr ? io_avail_list_22 : _GEN_981; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_983 = 6'h17 == buf_7_rs2_paddr ? io_avail_list_23 : _GEN_982; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_984 = 6'h18 == buf_7_rs2_paddr ? io_avail_list_24 : _GEN_983; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_985 = 6'h19 == buf_7_rs2_paddr ? io_avail_list_25 : _GEN_984; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_986 = 6'h1a == buf_7_rs2_paddr ? io_avail_list_26 : _GEN_985; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_987 = 6'h1b == buf_7_rs2_paddr ? io_avail_list_27 : _GEN_986; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_988 = 6'h1c == buf_7_rs2_paddr ? io_avail_list_28 : _GEN_987; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_989 = 6'h1d == buf_7_rs2_paddr ? io_avail_list_29 : _GEN_988; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_990 = 6'h1e == buf_7_rs2_paddr ? io_avail_list_30 : _GEN_989; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_991 = 6'h1f == buf_7_rs2_paddr ? io_avail_list_31 : _GEN_990; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_992 = 6'h20 == buf_7_rs2_paddr ? io_avail_list_32 : _GEN_991; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_993 = 6'h21 == buf_7_rs2_paddr ? io_avail_list_33 : _GEN_992; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_994 = 6'h22 == buf_7_rs2_paddr ? io_avail_list_34 : _GEN_993; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_995 = 6'h23 == buf_7_rs2_paddr ? io_avail_list_35 : _GEN_994; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_996 = 6'h24 == buf_7_rs2_paddr ? io_avail_list_36 : _GEN_995; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_997 = 6'h25 == buf_7_rs2_paddr ? io_avail_list_37 : _GEN_996; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_998 = 6'h26 == buf_7_rs2_paddr ? io_avail_list_38 : _GEN_997; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_999 = 6'h27 == buf_7_rs2_paddr ? io_avail_list_39 : _GEN_998; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1000 = 6'h28 == buf_7_rs2_paddr ? io_avail_list_40 : _GEN_999; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1001 = 6'h29 == buf_7_rs2_paddr ? io_avail_list_41 : _GEN_1000; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1002 = 6'h2a == buf_7_rs2_paddr ? io_avail_list_42 : _GEN_1001; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1003 = 6'h2b == buf_7_rs2_paddr ? io_avail_list_43 : _GEN_1002; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1004 = 6'h2c == buf_7_rs2_paddr ? io_avail_list_44 : _GEN_1003; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1005 = 6'h2d == buf_7_rs2_paddr ? io_avail_list_45 : _GEN_1004; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1006 = 6'h2e == buf_7_rs2_paddr ? io_avail_list_46 : _GEN_1005; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1007 = 6'h2f == buf_7_rs2_paddr ? io_avail_list_47 : _GEN_1006; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1008 = 6'h30 == buf_7_rs2_paddr ? io_avail_list_48 : _GEN_1007; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1009 = 6'h31 == buf_7_rs2_paddr ? io_avail_list_49 : _GEN_1008; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1010 = 6'h32 == buf_7_rs2_paddr ? io_avail_list_50 : _GEN_1009; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1011 = 6'h33 == buf_7_rs2_paddr ? io_avail_list_51 : _GEN_1010; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1012 = 6'h34 == buf_7_rs2_paddr ? io_avail_list_52 : _GEN_1011; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1013 = 6'h35 == buf_7_rs2_paddr ? io_avail_list_53 : _GEN_1012; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1014 = 6'h36 == buf_7_rs2_paddr ? io_avail_list_54 : _GEN_1013; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1015 = 6'h37 == buf_7_rs2_paddr ? io_avail_list_55 : _GEN_1014; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1016 = 6'h38 == buf_7_rs2_paddr ? io_avail_list_56 : _GEN_1015; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1017 = 6'h39 == buf_7_rs2_paddr ? io_avail_list_57 : _GEN_1016; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1018 = 6'h3a == buf_7_rs2_paddr ? io_avail_list_58 : _GEN_1017; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1019 = 6'h3b == buf_7_rs2_paddr ? io_avail_list_59 : _GEN_1018; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1020 = 6'h3c == buf_7_rs2_paddr ? io_avail_list_60 : _GEN_1019; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1021 = 6'h3d == buf_7_rs2_paddr ? io_avail_list_61 : _GEN_1020; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1022 = 6'h3e == buf_7_rs2_paddr ? io_avail_list_62 : _GEN_1021; // @[IssueUnit.scala 268:{32,32}]
  wire  _GEN_1023 = 6'h3f == buf_7_rs2_paddr ? io_avail_list_63 : _GEN_1022; // @[IssueUnit.scala 268:{32,32}]
  wire  ready_list_7 = _GEN_959 & _GEN_1023 & io_fu_ready & store_mask_7; // @[IssueUnit.scala 268:57]
  wire [7:0] rl0 = {ready_list_7,ready_list_6,ready_list_5,ready_list_4,ready_list_3,ready_list_2,ready_list_1,
    ready_list_0}; // @[Cat.scala 30:58]
  wire [2:0] _T_70 = rl0[6] ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _T_71 = rl0[5] ? 3'h5 : _T_70; // @[Mux.scala 47:69]
  wire [2:0] _T_72 = rl0[4] ? 3'h4 : _T_71; // @[Mux.scala 47:69]
  wire [2:0] _T_73 = rl0[3] ? 3'h3 : _T_72; // @[Mux.scala 47:69]
  wire [2:0] _T_74 = rl0[2] ? 3'h2 : _T_73; // @[Mux.scala 47:69]
  wire [2:0] _T_75 = rl0[1] ? 3'h1 : _T_74; // @[Mux.scala 47:69]
  wire [2:0] deq_vec_0 = rl0[0] ? 3'h0 : _T_75; // @[Mux.scala 47:69]
  wire  _GEN_1025 = 3'h1 == deq_vec_0 ? ready_list_1 : ready_list_0; // @[IssueUnit.scala 274:{20,20}]
  wire  _GEN_1026 = 3'h2 == deq_vec_0 ? ready_list_2 : _GEN_1025; // @[IssueUnit.scala 274:{20,20}]
  wire  _GEN_1027 = 3'h3 == deq_vec_0 ? ready_list_3 : _GEN_1026; // @[IssueUnit.scala 274:{20,20}]
  wire  _GEN_1028 = 3'h4 == deq_vec_0 ? ready_list_4 : _GEN_1027; // @[IssueUnit.scala 274:{20,20}]
  wire  _GEN_1029 = 3'h5 == deq_vec_0 ? ready_list_5 : _GEN_1028; // @[IssueUnit.scala 274:{20,20}]
  wire  _GEN_1030 = 3'h6 == deq_vec_0 ? ready_list_6 : _GEN_1029; // @[IssueUnit.scala 274:{20,20}]
  wire  deq_vec_valid_0 = 3'h7 == deq_vec_0 ? ready_list_7 : _GEN_1030; // @[IssueUnit.scala 274:{20,20}]
  wire [3:0] _GEN_1033 = 3'h1 == deq_vec_0 ? buf_1_rob_addr : buf_0_rob_addr; // @[IssueUnit.scala 278:{15,15}]
  wire [3:0] _GEN_1034 = 3'h2 == deq_vec_0 ? buf_2_rob_addr : _GEN_1033; // @[IssueUnit.scala 278:{15,15}]
  wire [3:0] _GEN_1035 = 3'h3 == deq_vec_0 ? buf_3_rob_addr : _GEN_1034; // @[IssueUnit.scala 278:{15,15}]
  wire [3:0] _GEN_1036 = 3'h4 == deq_vec_0 ? buf_4_rob_addr : _GEN_1035; // @[IssueUnit.scala 278:{15,15}]
  wire [3:0] _GEN_1037 = 3'h5 == deq_vec_0 ? buf_5_rob_addr : _GEN_1036; // @[IssueUnit.scala 278:{15,15}]
  wire [3:0] _GEN_1038 = 3'h6 == deq_vec_0 ? buf_6_rob_addr : _GEN_1037; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1049 = 3'h1 == deq_vec_0 ? buf_1_rd_paddr : buf_0_rd_paddr; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1050 = 3'h2 == deq_vec_0 ? buf_2_rd_paddr : _GEN_1049; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1051 = 3'h3 == deq_vec_0 ? buf_3_rd_paddr : _GEN_1050; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1052 = 3'h4 == deq_vec_0 ? buf_4_rd_paddr : _GEN_1051; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1053 = 3'h5 == deq_vec_0 ? buf_5_rd_paddr : _GEN_1052; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1054 = 3'h6 == deq_vec_0 ? buf_6_rd_paddr : _GEN_1053; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1057 = 3'h1 == deq_vec_0 ? buf_1_rs2_paddr : buf_0_rs2_paddr; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1058 = 3'h2 == deq_vec_0 ? buf_2_rs2_paddr : _GEN_1057; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1059 = 3'h3 == deq_vec_0 ? buf_3_rs2_paddr : _GEN_1058; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1060 = 3'h4 == deq_vec_0 ? buf_4_rs2_paddr : _GEN_1059; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1061 = 3'h5 == deq_vec_0 ? buf_5_rs2_paddr : _GEN_1060; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1062 = 3'h6 == deq_vec_0 ? buf_6_rs2_paddr : _GEN_1061; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1065 = 3'h1 == deq_vec_0 ? buf_1_rs1_paddr : buf_0_rs1_paddr; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1066 = 3'h2 == deq_vec_0 ? buf_2_rs1_paddr : _GEN_1065; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1067 = 3'h3 == deq_vec_0 ? buf_3_rs1_paddr : _GEN_1066; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1068 = 3'h4 == deq_vec_0 ? buf_4_rs1_paddr : _GEN_1067; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1069 = 3'h5 == deq_vec_0 ? buf_5_rs1_paddr : _GEN_1068; // @[IssueUnit.scala 278:{15,15}]
  wire [5:0] _GEN_1070 = 3'h6 == deq_vec_0 ? buf_6_rs1_paddr : _GEN_1069; // @[IssueUnit.scala 278:{15,15}]
  wire [31:0] _GEN_1089 = 3'h1 == deq_vec_0 ? buf_1_imm : buf_0_imm; // @[IssueUnit.scala 278:{15,15}]
  wire [31:0] _GEN_1090 = 3'h2 == deq_vec_0 ? buf_2_imm : _GEN_1089; // @[IssueUnit.scala 278:{15,15}]
  wire [31:0] _GEN_1091 = 3'h3 == deq_vec_0 ? buf_3_imm : _GEN_1090; // @[IssueUnit.scala 278:{15,15}]
  wire [31:0] _GEN_1092 = 3'h4 == deq_vec_0 ? buf_4_imm : _GEN_1091; // @[IssueUnit.scala 278:{15,15}]
  wire [31:0] _GEN_1093 = 3'h5 == deq_vec_0 ? buf_5_imm : _GEN_1092; // @[IssueUnit.scala 278:{15,15}]
  wire [31:0] _GEN_1094 = 3'h6 == deq_vec_0 ? buf_6_imm : _GEN_1093; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1097 = 3'h1 == deq_vec_0 ? buf_1_rd_en : buf_0_rd_en; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1098 = 3'h2 == deq_vec_0 ? buf_2_rd_en : _GEN_1097; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1099 = 3'h3 == deq_vec_0 ? buf_3_rd_en : _GEN_1098; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1100 = 3'h4 == deq_vec_0 ? buf_4_rd_en : _GEN_1099; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1101 = 3'h5 == deq_vec_0 ? buf_5_rd_en : _GEN_1100; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1102 = 3'h6 == deq_vec_0 ? buf_6_rd_en : _GEN_1101; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1129 = 3'h1 == deq_vec_0 ? buf_1_rs2_src : buf_0_rs2_src; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1130 = 3'h2 == deq_vec_0 ? buf_2_rs2_src : _GEN_1129; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1131 = 3'h3 == deq_vec_0 ? buf_3_rs2_src : _GEN_1130; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1132 = 3'h4 == deq_vec_0 ? buf_4_rs2_src : _GEN_1131; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1133 = 3'h5 == deq_vec_0 ? buf_5_rs2_src : _GEN_1132; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1134 = 3'h6 == deq_vec_0 ? buf_6_rs2_src : _GEN_1133; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1137 = 3'h1 == deq_vec_0 ? buf_1_rs1_src : buf_0_rs1_src; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1138 = 3'h2 == deq_vec_0 ? buf_2_rs1_src : _GEN_1137; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1139 = 3'h3 == deq_vec_0 ? buf_3_rs1_src : _GEN_1138; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1140 = 3'h4 == deq_vec_0 ? buf_4_rs1_src : _GEN_1139; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1141 = 3'h5 == deq_vec_0 ? buf_5_rs1_src : _GEN_1140; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1142 = 3'h6 == deq_vec_0 ? buf_6_rs1_src : _GEN_1141; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1145 = 3'h1 == deq_vec_0 ? buf_1_w_type : buf_0_w_type; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1146 = 3'h2 == deq_vec_0 ? buf_2_w_type : _GEN_1145; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1147 = 3'h3 == deq_vec_0 ? buf_3_w_type : _GEN_1146; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1148 = 3'h4 == deq_vec_0 ? buf_4_w_type : _GEN_1147; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1149 = 3'h5 == deq_vec_0 ? buf_5_w_type : _GEN_1148; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1150 = 3'h6 == deq_vec_0 ? buf_6_w_type : _GEN_1149; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1161 = 3'h1 == deq_vec_0 ? buf_1_mem_size : buf_0_mem_size; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1162 = 3'h2 == deq_vec_0 ? buf_2_mem_size : _GEN_1161; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1163 = 3'h3 == deq_vec_0 ? buf_3_mem_size : _GEN_1162; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1164 = 3'h4 == deq_vec_0 ? buf_4_mem_size : _GEN_1163; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1165 = 3'h5 == deq_vec_0 ? buf_5_mem_size : _GEN_1164; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1166 = 3'h6 == deq_vec_0 ? buf_6_mem_size : _GEN_1165; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1169 = 3'h1 == deq_vec_0 ? buf_1_mem_code : buf_0_mem_code; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1170 = 3'h2 == deq_vec_0 ? buf_2_mem_code : _GEN_1169; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1171 = 3'h3 == deq_vec_0 ? buf_3_mem_code : _GEN_1170; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1172 = 3'h4 == deq_vec_0 ? buf_4_mem_code : _GEN_1171; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1173 = 3'h5 == deq_vec_0 ? buf_5_mem_code : _GEN_1172; // @[IssueUnit.scala 278:{15,15}]
  wire [1:0] _GEN_1174 = 3'h6 == deq_vec_0 ? buf_6_mem_code : _GEN_1173; // @[IssueUnit.scala 278:{15,15}]
  wire [3:0] _GEN_1185 = 3'h1 == deq_vec_0 ? buf_1_alu_code : buf_0_alu_code; // @[IssueUnit.scala 278:{15,15}]
  wire [3:0] _GEN_1186 = 3'h2 == deq_vec_0 ? buf_2_alu_code : _GEN_1185; // @[IssueUnit.scala 278:{15,15}]
  wire [3:0] _GEN_1187 = 3'h3 == deq_vec_0 ? buf_3_alu_code : _GEN_1186; // @[IssueUnit.scala 278:{15,15}]
  wire [3:0] _GEN_1188 = 3'h4 == deq_vec_0 ? buf_4_alu_code : _GEN_1187; // @[IssueUnit.scala 278:{15,15}]
  wire [3:0] _GEN_1189 = 3'h5 == deq_vec_0 ? buf_5_alu_code : _GEN_1188; // @[IssueUnit.scala 278:{15,15}]
  wire [3:0] _GEN_1190 = 3'h6 == deq_vec_0 ? buf_6_alu_code : _GEN_1189; // @[IssueUnit.scala 278:{15,15}]
  wire [2:0] _GEN_1193 = 3'h1 == deq_vec_0 ? buf_1_fu_code : buf_0_fu_code; // @[IssueUnit.scala 278:{15,15}]
  wire [2:0] _GEN_1194 = 3'h2 == deq_vec_0 ? buf_2_fu_code : _GEN_1193; // @[IssueUnit.scala 278:{15,15}]
  wire [2:0] _GEN_1195 = 3'h3 == deq_vec_0 ? buf_3_fu_code : _GEN_1194; // @[IssueUnit.scala 278:{15,15}]
  wire [2:0] _GEN_1196 = 3'h4 == deq_vec_0 ? buf_4_fu_code : _GEN_1195; // @[IssueUnit.scala 278:{15,15}]
  wire [2:0] _GEN_1197 = 3'h5 == deq_vec_0 ? buf_5_fu_code : _GEN_1196; // @[IssueUnit.scala 278:{15,15}]
  wire [2:0] _GEN_1198 = 3'h6 == deq_vec_0 ? buf_6_fu_code : _GEN_1197; // @[IssueUnit.scala 278:{15,15}]
  wire [31:0] _GEN_1217 = 3'h1 == deq_vec_0 ? buf_1_pc : buf_0_pc; // @[IssueUnit.scala 278:{15,15}]
  wire [31:0] _GEN_1218 = 3'h2 == deq_vec_0 ? buf_2_pc : _GEN_1217; // @[IssueUnit.scala 278:{15,15}]
  wire [31:0] _GEN_1219 = 3'h3 == deq_vec_0 ? buf_3_pc : _GEN_1218; // @[IssueUnit.scala 278:{15,15}]
  wire [31:0] _GEN_1220 = 3'h4 == deq_vec_0 ? buf_4_pc : _GEN_1219; // @[IssueUnit.scala 278:{15,15}]
  wire [31:0] _GEN_1221 = 3'h5 == deq_vec_0 ? buf_5_pc : _GEN_1220; // @[IssueUnit.scala 278:{15,15}]
  wire [31:0] _GEN_1222 = 3'h6 == deq_vec_0 ? buf_6_pc : _GEN_1221; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1225 = 3'h1 == deq_vec_0 ? buf_1_valid : buf_0_valid; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1226 = 3'h2 == deq_vec_0 ? buf_2_valid : _GEN_1225; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1227 = 3'h3 == deq_vec_0 ? buf_3_valid : _GEN_1226; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1228 = 3'h4 == deq_vec_0 ? buf_4_valid : _GEN_1227; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1229 = 3'h5 == deq_vec_0 ? buf_5_valid : _GEN_1228; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1230 = 3'h6 == deq_vec_0 ? buf_6_valid : _GEN_1229; // @[IssueUnit.scala 278:{15,15}]
  wire  _GEN_1231 = 3'h7 == deq_vec_0 ? buf_7_valid : _GEN_1230; // @[IssueUnit.scala 278:{15,15}]
  wire  up1_0 = 3'h0 >= deq_vec_0 & deq_vec_valid_0; // @[IssueUnit.scala 286:35]
  wire  up1_1 = 3'h1 >= deq_vec_0 & deq_vec_valid_0; // @[IssueUnit.scala 286:35]
  wire  up1_2 = 3'h2 >= deq_vec_0 & deq_vec_valid_0; // @[IssueUnit.scala 286:35]
  wire  up1_3 = 3'h3 >= deq_vec_0 & deq_vec_valid_0; // @[IssueUnit.scala 286:35]
  wire  up1_4 = 3'h4 >= deq_vec_0 & deq_vec_valid_0; // @[IssueUnit.scala 286:35]
  wire  up1_5 = 3'h5 >= deq_vec_0 & deq_vec_valid_0; // @[IssueUnit.scala 286:35]
  wire  up1_6 = 3'h6 >= deq_vec_0 & deq_vec_valid_0; // @[IssueUnit.scala 286:35]
  wire [3:0] _GEN_1232 = up1_0 ? buf_1_rob_addr : buf_0_rob_addr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1234 = up1_0 ? buf_1_rd_paddr : buf_0_rd_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1235 = up1_0 ? buf_1_rs2_paddr : buf_0_rs2_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1236 = up1_0 ? buf_1_rs1_paddr : buf_0_rs1_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [31:0] _GEN_1239 = up1_0 ? buf_1_imm : buf_0_imm; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1240 = up1_0 ? buf_1_rd_en : buf_0_rd_en; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1244 = up1_0 ? buf_1_rs2_src : buf_0_rs2_src; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1245 = up1_0 ? buf_1_rs1_src : buf_0_rs1_src; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1246 = up1_0 ? buf_1_w_type : buf_0_w_type; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1248 = up1_0 ? buf_1_mem_size : buf_0_mem_size; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1249 = up1_0 ? buf_1_mem_code : buf_0_mem_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [3:0] _GEN_1251 = up1_0 ? buf_1_alu_code : buf_0_alu_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [2:0] _GEN_1252 = up1_0 ? buf_1_fu_code : buf_0_fu_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [31:0] _GEN_1255 = up1_0 ? buf_1_pc : buf_0_pc; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1256 = up1_0 ? buf_1_valid : buf_0_valid; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [3:0] _GEN_1257 = up1_1 ? buf_2_rob_addr : buf_1_rob_addr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1259 = up1_1 ? buf_2_rd_paddr : buf_1_rd_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1260 = up1_1 ? buf_2_rs2_paddr : buf_1_rs2_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1261 = up1_1 ? buf_2_rs1_paddr : buf_1_rs1_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [31:0] _GEN_1264 = up1_1 ? buf_2_imm : buf_1_imm; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1265 = up1_1 ? buf_2_rd_en : buf_1_rd_en; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1269 = up1_1 ? buf_2_rs2_src : buf_1_rs2_src; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1270 = up1_1 ? buf_2_rs1_src : buf_1_rs1_src; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1271 = up1_1 ? buf_2_w_type : buf_1_w_type; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1273 = up1_1 ? buf_2_mem_size : buf_1_mem_size; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1274 = up1_1 ? buf_2_mem_code : buf_1_mem_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [3:0] _GEN_1276 = up1_1 ? buf_2_alu_code : buf_1_alu_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [2:0] _GEN_1277 = up1_1 ? buf_2_fu_code : buf_1_fu_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [31:0] _GEN_1280 = up1_1 ? buf_2_pc : buf_1_pc; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1281 = up1_1 ? buf_2_valid : buf_1_valid; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [3:0] _GEN_1282 = up1_2 ? buf_3_rob_addr : buf_2_rob_addr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1284 = up1_2 ? buf_3_rd_paddr : buf_2_rd_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1285 = up1_2 ? buf_3_rs2_paddr : buf_2_rs2_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1286 = up1_2 ? buf_3_rs1_paddr : buf_2_rs1_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [31:0] _GEN_1289 = up1_2 ? buf_3_imm : buf_2_imm; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1290 = up1_2 ? buf_3_rd_en : buf_2_rd_en; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1294 = up1_2 ? buf_3_rs2_src : buf_2_rs2_src; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1295 = up1_2 ? buf_3_rs1_src : buf_2_rs1_src; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1296 = up1_2 ? buf_3_w_type : buf_2_w_type; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1298 = up1_2 ? buf_3_mem_size : buf_2_mem_size; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1299 = up1_2 ? buf_3_mem_code : buf_2_mem_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [3:0] _GEN_1301 = up1_2 ? buf_3_alu_code : buf_2_alu_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [2:0] _GEN_1302 = up1_2 ? buf_3_fu_code : buf_2_fu_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [31:0] _GEN_1305 = up1_2 ? buf_3_pc : buf_2_pc; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1306 = up1_2 ? buf_3_valid : buf_2_valid; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [3:0] _GEN_1307 = up1_3 ? buf_4_rob_addr : buf_3_rob_addr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1309 = up1_3 ? buf_4_rd_paddr : buf_3_rd_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1310 = up1_3 ? buf_4_rs2_paddr : buf_3_rs2_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1311 = up1_3 ? buf_4_rs1_paddr : buf_3_rs1_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [31:0] _GEN_1314 = up1_3 ? buf_4_imm : buf_3_imm; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1315 = up1_3 ? buf_4_rd_en : buf_3_rd_en; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1319 = up1_3 ? buf_4_rs2_src : buf_3_rs2_src; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1320 = up1_3 ? buf_4_rs1_src : buf_3_rs1_src; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1321 = up1_3 ? buf_4_w_type : buf_3_w_type; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1323 = up1_3 ? buf_4_mem_size : buf_3_mem_size; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1324 = up1_3 ? buf_4_mem_code : buf_3_mem_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [3:0] _GEN_1326 = up1_3 ? buf_4_alu_code : buf_3_alu_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [2:0] _GEN_1327 = up1_3 ? buf_4_fu_code : buf_3_fu_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [31:0] _GEN_1330 = up1_3 ? buf_4_pc : buf_3_pc; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1331 = up1_3 ? buf_4_valid : buf_3_valid; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [3:0] _GEN_1332 = up1_4 ? buf_5_rob_addr : buf_4_rob_addr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1334 = up1_4 ? buf_5_rd_paddr : buf_4_rd_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1335 = up1_4 ? buf_5_rs2_paddr : buf_4_rs2_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1336 = up1_4 ? buf_5_rs1_paddr : buf_4_rs1_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [31:0] _GEN_1339 = up1_4 ? buf_5_imm : buf_4_imm; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1340 = up1_4 ? buf_5_rd_en : buf_4_rd_en; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1344 = up1_4 ? buf_5_rs2_src : buf_4_rs2_src; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1345 = up1_4 ? buf_5_rs1_src : buf_4_rs1_src; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1346 = up1_4 ? buf_5_w_type : buf_4_w_type; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1348 = up1_4 ? buf_5_mem_size : buf_4_mem_size; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1349 = up1_4 ? buf_5_mem_code : buf_4_mem_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [3:0] _GEN_1351 = up1_4 ? buf_5_alu_code : buf_4_alu_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [2:0] _GEN_1352 = up1_4 ? buf_5_fu_code : buf_4_fu_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [31:0] _GEN_1355 = up1_4 ? buf_5_pc : buf_4_pc; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1356 = up1_4 ? buf_5_valid : buf_4_valid; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [3:0] _GEN_1357 = up1_5 ? buf_6_rob_addr : buf_5_rob_addr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1359 = up1_5 ? buf_6_rd_paddr : buf_5_rd_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1360 = up1_5 ? buf_6_rs2_paddr : buf_5_rs2_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1361 = up1_5 ? buf_6_rs1_paddr : buf_5_rs1_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [31:0] _GEN_1364 = up1_5 ? buf_6_imm : buf_5_imm; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1365 = up1_5 ? buf_6_rd_en : buf_5_rd_en; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1369 = up1_5 ? buf_6_rs2_src : buf_5_rs2_src; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1370 = up1_5 ? buf_6_rs1_src : buf_5_rs1_src; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1371 = up1_5 ? buf_6_w_type : buf_5_w_type; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1373 = up1_5 ? buf_6_mem_size : buf_5_mem_size; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1374 = up1_5 ? buf_6_mem_code : buf_5_mem_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [3:0] _GEN_1376 = up1_5 ? buf_6_alu_code : buf_5_alu_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [2:0] _GEN_1377 = up1_5 ? buf_6_fu_code : buf_5_fu_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [31:0] _GEN_1380 = up1_5 ? buf_6_pc : buf_5_pc; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1381 = up1_5 ? buf_6_valid : buf_5_valid; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [3:0] _GEN_1382 = up1_6 ? buf_7_rob_addr : buf_6_rob_addr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1384 = up1_6 ? buf_7_rd_paddr : buf_6_rd_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1385 = up1_6 ? buf_7_rs2_paddr : buf_6_rs2_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [5:0] _GEN_1386 = up1_6 ? buf_7_rs1_paddr : buf_6_rs1_paddr; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [31:0] _GEN_1389 = up1_6 ? buf_7_imm : buf_6_imm; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1390 = up1_6 ? buf_7_rd_en : buf_6_rd_en; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1394 = up1_6 ? buf_7_rs2_src : buf_6_rs2_src; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1395 = up1_6 ? buf_7_rs1_src : buf_6_rs1_src; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1396 = up1_6 ? buf_7_w_type : buf_6_w_type; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1398 = up1_6 ? buf_7_mem_size : buf_6_mem_size; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [1:0] _GEN_1399 = up1_6 ? buf_7_mem_code : buf_6_mem_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [3:0] _GEN_1401 = up1_6 ? buf_7_alu_code : buf_6_alu_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [2:0] _GEN_1402 = up1_6 ? buf_7_fu_code : buf_6_fu_code; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [31:0] _GEN_1405 = up1_6 ? buf_7_pc : buf_6_pc; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire  _GEN_1406 = up1_6 ? buf_7_valid : buf_6_valid; // @[IssueUnit.scala 289:19 291:18 97:20]
  wire [3:0] _GEN_1407 = deq_vec_valid_0 ? 4'h0 : buf_7_rob_addr; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire [5:0] _GEN_1409 = deq_vec_valid_0 ? 6'h0 : buf_7_rd_paddr; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire [5:0] _GEN_1410 = deq_vec_valid_0 ? 6'h0 : buf_7_rs2_paddr; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire [5:0] _GEN_1411 = deq_vec_valid_0 ? 6'h0 : buf_7_rs1_paddr; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire [31:0] _GEN_1414 = deq_vec_valid_0 ? 32'h0 : buf_7_imm; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire  _GEN_1415 = deq_vec_valid_0 ? 1'h0 : buf_7_rd_en; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire [1:0] _GEN_1419 = deq_vec_valid_0 ? 2'h0 : buf_7_rs2_src; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire [1:0] _GEN_1420 = deq_vec_valid_0 ? 2'h0 : buf_7_rs1_src; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire  _GEN_1421 = deq_vec_valid_0 ? 1'h0 : buf_7_w_type; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire [1:0] _GEN_1423 = deq_vec_valid_0 ? 2'h0 : buf_7_mem_size; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire [1:0] _GEN_1424 = deq_vec_valid_0 ? 2'h0 : buf_7_mem_code; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire [3:0] _GEN_1426 = deq_vec_valid_0 ? 4'h0 : buf_7_alu_code; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire [2:0] _GEN_1427 = deq_vec_valid_0 ? 3'h0 : buf_7_fu_code; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire [31:0] _GEN_1430 = deq_vec_valid_0 ? 32'h0 : buf_7_pc; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire  _GEN_1431 = deq_vec_valid_0 ? 1'h0 : buf_7_valid; // @[IssueUnit.scala 289:19 293:18 97:20]
  wire  _T_97 = ~io_flush; // @[IssueUnit.scala 315:40]
  wire [3:0] _GEN_1434 = 3'h0 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1232; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1435 = 3'h1 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1257; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1436 = 3'h2 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1282; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1437 = 3'h3 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1307; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1438 = 3'h4 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1332; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1439 = 3'h5 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1357; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1440 = 3'h6 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1382; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1441 = 3'h7 == enq_vec_real_0[2:0] ? io_rob_addr_0 : _GEN_1407; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1450 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1234; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1451 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1259; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1452 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1284; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1453 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1309; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1454 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1334; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1455 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1359; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1456 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1384; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1457 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_paddr : _GEN_1409; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1458 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1235; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1459 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1260; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1460 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1285; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1461 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1310; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1462 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1335; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1463 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1360; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1464 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1385; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1465 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_paddr : _GEN_1410; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1466 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1236; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1467 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1261; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1468 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1286; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1469 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1311; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1470 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1336; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1471 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1361; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1472 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1386; // @[IssueUnit.scala 316:{48,48}]
  wire [5:0] _GEN_1473 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_paddr : _GEN_1411; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1490 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1239; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1491 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1264; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1492 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1289; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1493 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1314; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1494 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1339; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1495 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1364; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1496 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1389; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1497 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_imm : _GEN_1414; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1498 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1240; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1499 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1265; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1500 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1290; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1501 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1315; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1502 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1340; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1503 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1365; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1504 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1390; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1505 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rd_en : _GEN_1415; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1530 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1244; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1531 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1269; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1532 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1294; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1533 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1319; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1534 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1344; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1535 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1369; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1536 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1394; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1537 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs2_src : _GEN_1419; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1538 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1245; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1539 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1270; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1540 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1295; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1541 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1320; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1542 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1345; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1543 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1370; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1544 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1395; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1545 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_rs1_src : _GEN_1420; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1546 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1246; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1547 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1271; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1548 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1296; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1549 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1321; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1550 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1346; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1551 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1371; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1552 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1396; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1553 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_w_type : _GEN_1421; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1562 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_size : _GEN_1248; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1563 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_size : _GEN_1273; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1564 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_size : _GEN_1298; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1565 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_size : _GEN_1323; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1566 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_size : _GEN_1348; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1567 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_size : _GEN_1373; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1568 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_size : _GEN_1398; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1569 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_size : _GEN_1423; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1570 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_code : _GEN_1249; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1571 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_code : _GEN_1274; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1572 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_code : _GEN_1299; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1573 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_code : _GEN_1324; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1574 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_code : _GEN_1349; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1575 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_code : _GEN_1374; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1576 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_code : _GEN_1399; // @[IssueUnit.scala 316:{48,48}]
  wire [1:0] _GEN_1577 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_mem_code : _GEN_1424; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1586 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1251; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1587 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1276; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1588 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1301; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1589 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1326; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1590 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1351; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1591 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1376; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1592 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1401; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1593 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_alu_code : _GEN_1426; // @[IssueUnit.scala 316:{48,48}]
  wire [2:0] _GEN_1594 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1252; // @[IssueUnit.scala 316:{48,48}]
  wire [2:0] _GEN_1595 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1277; // @[IssueUnit.scala 316:{48,48}]
  wire [2:0] _GEN_1596 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1302; // @[IssueUnit.scala 316:{48,48}]
  wire [2:0] _GEN_1597 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1327; // @[IssueUnit.scala 316:{48,48}]
  wire [2:0] _GEN_1598 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1352; // @[IssueUnit.scala 316:{48,48}]
  wire [2:0] _GEN_1599 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1377; // @[IssueUnit.scala 316:{48,48}]
  wire [2:0] _GEN_1600 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1402; // @[IssueUnit.scala 316:{48,48}]
  wire [2:0] _GEN_1601 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_fu_code : _GEN_1427; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1618 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1255; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1619 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1280; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1620 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1305; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1621 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1330; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1622 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1355; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1623 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1380; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1624 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1405; // @[IssueUnit.scala 316:{48,48}]
  wire [31:0] _GEN_1625 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_pc : _GEN_1430; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1626 = 3'h0 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1256; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1627 = 3'h1 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1281; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1628 = 3'h2 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1306; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1629 = 3'h3 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1331; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1630 = 3'h4 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1356; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1631 = 3'h5 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1381; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1632 = 3'h6 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1406; // @[IssueUnit.scala 316:{48,48}]
  wire  _GEN_1633 = 3'h7 == enq_vec_real_0[2:0] ? io_in_bits_vec_0_valid : _GEN_1431; // @[IssueUnit.scala 316:{48,48}]
  wire [3:0] _GEN_1634 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1434 : _GEN_1232; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1635 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1435 : _GEN_1257; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1636 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1436 : _GEN_1282; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1637 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1437 : _GEN_1307; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1638 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1438 : _GEN_1332; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1639 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1439 : _GEN_1357; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1640 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1440 : _GEN_1382; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1641 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1441 : _GEN_1407; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1650 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1450 : _GEN_1234; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1651 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1451 : _GEN_1259; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1652 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1452 : _GEN_1284; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1653 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1453 : _GEN_1309; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1654 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1454 : _GEN_1334; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1655 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1455 : _GEN_1359; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1656 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1456 : _GEN_1384; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1657 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1457 : _GEN_1409; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1658 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1458 : _GEN_1235; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1659 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1459 : _GEN_1260; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1660 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1460 : _GEN_1285; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1661 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1461 : _GEN_1310; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1662 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1462 : _GEN_1335; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1663 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1463 : _GEN_1360; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1664 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1464 : _GEN_1385; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1665 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1465 : _GEN_1410; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1666 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1466 : _GEN_1236; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1667 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1467 : _GEN_1261; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1668 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1468 : _GEN_1286; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1669 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1469 : _GEN_1311; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1670 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1470 : _GEN_1336; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1671 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1471 : _GEN_1361; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1672 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1472 : _GEN_1386; // @[IssueUnit.scala 315:51]
  wire [5:0] _GEN_1673 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1473 : _GEN_1411; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1690 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1490 : _GEN_1239; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1691 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1491 : _GEN_1264; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1692 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1492 : _GEN_1289; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1693 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1493 : _GEN_1314; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1694 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1494 : _GEN_1339; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1695 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1495 : _GEN_1364; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1696 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1496 : _GEN_1389; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1697 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1497 : _GEN_1414; // @[IssueUnit.scala 315:51]
  wire  _GEN_1698 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1498 : _GEN_1240; // @[IssueUnit.scala 315:51]
  wire  _GEN_1699 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1499 : _GEN_1265; // @[IssueUnit.scala 315:51]
  wire  _GEN_1700 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1500 : _GEN_1290; // @[IssueUnit.scala 315:51]
  wire  _GEN_1701 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1501 : _GEN_1315; // @[IssueUnit.scala 315:51]
  wire  _GEN_1702 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1502 : _GEN_1340; // @[IssueUnit.scala 315:51]
  wire  _GEN_1703 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1503 : _GEN_1365; // @[IssueUnit.scala 315:51]
  wire  _GEN_1704 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1504 : _GEN_1390; // @[IssueUnit.scala 315:51]
  wire  _GEN_1705 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1505 : _GEN_1415; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1730 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1530 : _GEN_1244; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1731 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1531 : _GEN_1269; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1732 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1532 : _GEN_1294; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1733 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1533 : _GEN_1319; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1734 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1534 : _GEN_1344; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1735 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1535 : _GEN_1369; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1736 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1536 : _GEN_1394; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1737 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1537 : _GEN_1419; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1738 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1538 : _GEN_1245; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1739 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1539 : _GEN_1270; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1740 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1540 : _GEN_1295; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1741 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1541 : _GEN_1320; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1742 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1542 : _GEN_1345; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1743 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1543 : _GEN_1370; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1744 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1544 : _GEN_1395; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1745 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1545 : _GEN_1420; // @[IssueUnit.scala 315:51]
  wire  _GEN_1746 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1546 : _GEN_1246; // @[IssueUnit.scala 315:51]
  wire  _GEN_1747 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1547 : _GEN_1271; // @[IssueUnit.scala 315:51]
  wire  _GEN_1748 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1548 : _GEN_1296; // @[IssueUnit.scala 315:51]
  wire  _GEN_1749 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1549 : _GEN_1321; // @[IssueUnit.scala 315:51]
  wire  _GEN_1750 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1550 : _GEN_1346; // @[IssueUnit.scala 315:51]
  wire  _GEN_1751 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1551 : _GEN_1371; // @[IssueUnit.scala 315:51]
  wire  _GEN_1752 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1552 : _GEN_1396; // @[IssueUnit.scala 315:51]
  wire  _GEN_1753 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1553 : _GEN_1421; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1762 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1562 : _GEN_1248; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1763 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1563 : _GEN_1273; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1764 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1564 : _GEN_1298; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1765 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1565 : _GEN_1323; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1766 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1566 : _GEN_1348; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1767 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1567 : _GEN_1373; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1768 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1568 : _GEN_1398; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1769 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1569 : _GEN_1423; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1770 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1570 : _GEN_1249; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1771 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1571 : _GEN_1274; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1772 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1572 : _GEN_1299; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1773 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1573 : _GEN_1324; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1774 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1574 : _GEN_1349; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1775 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1575 : _GEN_1374; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1776 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1576 : _GEN_1399; // @[IssueUnit.scala 315:51]
  wire [1:0] _GEN_1777 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1577 : _GEN_1424; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1786 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1586 : _GEN_1251; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1787 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1587 : _GEN_1276; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1788 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1588 : _GEN_1301; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1789 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1589 : _GEN_1326; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1790 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1590 : _GEN_1351; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1791 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1591 : _GEN_1376; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1792 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1592 : _GEN_1401; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1793 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1593 : _GEN_1426; // @[IssueUnit.scala 315:51]
  wire [2:0] _GEN_1794 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1594 : _GEN_1252; // @[IssueUnit.scala 315:51]
  wire [2:0] _GEN_1795 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1595 : _GEN_1277; // @[IssueUnit.scala 315:51]
  wire [2:0] _GEN_1796 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1596 : _GEN_1302; // @[IssueUnit.scala 315:51]
  wire [2:0] _GEN_1797 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1597 : _GEN_1327; // @[IssueUnit.scala 315:51]
  wire [2:0] _GEN_1798 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1598 : _GEN_1352; // @[IssueUnit.scala 315:51]
  wire [2:0] _GEN_1799 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1599 : _GEN_1377; // @[IssueUnit.scala 315:51]
  wire [2:0] _GEN_1800 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1600 : _GEN_1402; // @[IssueUnit.scala 315:51]
  wire [2:0] _GEN_1801 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1601 : _GEN_1427; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1818 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1618 : _GEN_1255; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1819 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1619 : _GEN_1280; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1820 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1620 : _GEN_1305; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1821 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1621 : _GEN_1330; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1822 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1622 : _GEN_1355; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1823 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1623 : _GEN_1380; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1824 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1624 : _GEN_1405; // @[IssueUnit.scala 315:51]
  wire [31:0] _GEN_1825 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1625 : _GEN_1430; // @[IssueUnit.scala 315:51]
  wire  _GEN_1826 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1626 : _GEN_1256; // @[IssueUnit.scala 315:51]
  wire  _GEN_1827 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1627 : _GEN_1281; // @[IssueUnit.scala 315:51]
  wire  _GEN_1828 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1628 : _GEN_1306; // @[IssueUnit.scala 315:51]
  wire  _GEN_1829 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1629 : _GEN_1331; // @[IssueUnit.scala 315:51]
  wire  _GEN_1830 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1630 : _GEN_1356; // @[IssueUnit.scala 315:51]
  wire  _GEN_1831 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1631 : _GEN_1381; // @[IssueUnit.scala 315:51]
  wire  _GEN_1832 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1632 : _GEN_1406; // @[IssueUnit.scala 315:51]
  wire  _GEN_1833 = io_in_bits_vec_0_valid & _T & ~io_flush ? _GEN_1633 : _GEN_1431; // @[IssueUnit.scala 315:51]
  wire [3:0] _GEN_1835 = io_in_bits_vec_0_valid ? enq_vec_real_1 : enq_vec_real_0; // @[IssueUnit.scala 95:{32,32}]
  wire [3:0] _GEN_2442 = {{2'd0}, num_enq}; // @[IssueUnit.scala 320:44]
  wire [3:0] _T_106 = enq_vec_0 + _GEN_2442; // @[IssueUnit.scala 320:44]
  wire [3:0] next_enq_vec_0 = _T_106 - _GEN_2440; // @[IssueUnit.scala 320:54]
  wire [3:0] _T_110 = enq_vec_1 + _GEN_2442; // @[IssueUnit.scala 320:44]
  wire [3:0] next_enq_vec_1 = _T_110 - _GEN_2440; // @[IssueUnit.scala 320:54]
  assign io_in_ready = enq_vec_real_0 <= 4'h6; // @[IssueUnit.scala 106:27]
  assign io_out_0_valid = _GEN_1231 & deq_vec_valid_0; // @[IssueUnit.scala 279:34]
  assign io_out_0_pc = 3'h7 == deq_vec_0 ? buf_7_pc : _GEN_1222; // @[IssueUnit.scala 278:{15,15}]
  assign io_out_0_fu_code = 3'h7 == deq_vec_0 ? buf_7_fu_code : _GEN_1198; // @[IssueUnit.scala 278:{15,15}]
  assign io_out_0_alu_code = 3'h7 == deq_vec_0 ? buf_7_alu_code : _GEN_1190; // @[IssueUnit.scala 278:{15,15}]
  assign io_out_0_mem_code = 3'h7 == deq_vec_0 ? buf_7_mem_code : _GEN_1174; // @[IssueUnit.scala 278:{15,15}]
  assign io_out_0_mem_size = 3'h7 == deq_vec_0 ? buf_7_mem_size : _GEN_1166; // @[IssueUnit.scala 278:{15,15}]
  assign io_out_0_w_type = 3'h7 == deq_vec_0 ? buf_7_w_type : _GEN_1150; // @[IssueUnit.scala 278:{15,15}]
  assign io_out_0_rs1_src = 3'h7 == deq_vec_0 ? buf_7_rs1_src : _GEN_1142; // @[IssueUnit.scala 278:{15,15}]
  assign io_out_0_rs2_src = 3'h7 == deq_vec_0 ? buf_7_rs2_src : _GEN_1134; // @[IssueUnit.scala 278:{15,15}]
  assign io_out_0_rd_en = 3'h7 == deq_vec_0 ? buf_7_rd_en : _GEN_1102; // @[IssueUnit.scala 278:{15,15}]
  assign io_out_0_imm = 3'h7 == deq_vec_0 ? buf_7_imm : _GEN_1094; // @[IssueUnit.scala 278:{15,15}]
  assign io_out_0_rs1_paddr = 3'h7 == deq_vec_0 ? buf_7_rs1_paddr : _GEN_1070; // @[IssueUnit.scala 278:{15,15}]
  assign io_out_0_rs2_paddr = 3'h7 == deq_vec_0 ? buf_7_rs2_paddr : _GEN_1062; // @[IssueUnit.scala 278:{15,15}]
  assign io_out_0_rd_paddr = 3'h7 == deq_vec_0 ? buf_7_rd_paddr : _GEN_1054; // @[IssueUnit.scala 278:{15,15}]
  assign io_out_0_rob_addr = 3'h7 == deq_vec_0 ? buf_7_rob_addr : _GEN_1038; // @[IssueUnit.scala 278:{15,15}]
  always @(posedge clock) begin
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_valid <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_valid <= _GEN_1826;
      end
    end else begin
      buf_0_valid <= _GEN_1826;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_pc <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_pc <= _GEN_1818;
      end
    end else begin
      buf_0_pc <= _GEN_1818;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_fu_code <= 3'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_fu_code <= _GEN_1794;
      end
    end else begin
      buf_0_fu_code <= _GEN_1794;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_alu_code <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_alu_code <= _GEN_1786;
      end
    end else begin
      buf_0_alu_code <= _GEN_1786;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_mem_code <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_mem_code <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_mem_code <= io_in_bits_vec_1_mem_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_mem_code <= _GEN_1770;
      end
    end else begin
      buf_0_mem_code <= _GEN_1770;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_mem_size <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_mem_size <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_mem_size <= io_in_bits_vec_1_mem_size; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_mem_size <= _GEN_1762;
      end
    end else begin
      buf_0_mem_size <= _GEN_1762;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_w_type <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_w_type <= _GEN_1746;
      end
    end else begin
      buf_0_w_type <= _GEN_1746;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_rs1_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_rs1_src <= _GEN_1738;
      end
    end else begin
      buf_0_rs1_src <= _GEN_1738;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_rs2_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_rs2_src <= _GEN_1730;
      end
    end else begin
      buf_0_rs2_src <= _GEN_1730;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_rd_en <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_rd_en <= _GEN_1698;
      end
    end else begin
      buf_0_rd_en <= _GEN_1698;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_imm <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_imm <= _GEN_1690;
      end
    end else begin
      buf_0_imm <= _GEN_1690;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_rs1_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_rs1_paddr <= _GEN_1666;
      end
    end else begin
      buf_0_rs1_paddr <= _GEN_1666;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_rs2_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_rs2_paddr <= _GEN_1658;
      end
    end else begin
      buf_0_rs2_paddr <= _GEN_1658;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_rd_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_rd_paddr <= _GEN_1650;
      end
    end else begin
      buf_0_rd_paddr <= _GEN_1650;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_0_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_0_rob_addr <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h0 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_0_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 316:48]
      end else begin
        buf_0_rob_addr <= _GEN_1634;
      end
    end else begin
      buf_0_rob_addr <= _GEN_1634;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_valid <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_valid <= _GEN_1827;
      end
    end else begin
      buf_1_valid <= _GEN_1827;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_pc <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_pc <= _GEN_1819;
      end
    end else begin
      buf_1_pc <= _GEN_1819;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_fu_code <= 3'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_fu_code <= _GEN_1795;
      end
    end else begin
      buf_1_fu_code <= _GEN_1795;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_alu_code <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_alu_code <= _GEN_1787;
      end
    end else begin
      buf_1_alu_code <= _GEN_1787;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_mem_code <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_mem_code <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_mem_code <= io_in_bits_vec_1_mem_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_mem_code <= _GEN_1771;
      end
    end else begin
      buf_1_mem_code <= _GEN_1771;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_mem_size <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_mem_size <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_mem_size <= io_in_bits_vec_1_mem_size; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_mem_size <= _GEN_1763;
      end
    end else begin
      buf_1_mem_size <= _GEN_1763;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_w_type <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_w_type <= _GEN_1747;
      end
    end else begin
      buf_1_w_type <= _GEN_1747;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_rs1_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_rs1_src <= _GEN_1739;
      end
    end else begin
      buf_1_rs1_src <= _GEN_1739;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_rs2_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_rs2_src <= _GEN_1731;
      end
    end else begin
      buf_1_rs2_src <= _GEN_1731;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_rd_en <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_rd_en <= _GEN_1699;
      end
    end else begin
      buf_1_rd_en <= _GEN_1699;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_imm <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_imm <= _GEN_1691;
      end
    end else begin
      buf_1_imm <= _GEN_1691;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_rs1_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_rs1_paddr <= _GEN_1667;
      end
    end else begin
      buf_1_rs1_paddr <= _GEN_1667;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_rs2_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_rs2_paddr <= _GEN_1659;
      end
    end else begin
      buf_1_rs2_paddr <= _GEN_1659;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_rd_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_rd_paddr <= _GEN_1651;
      end
    end else begin
      buf_1_rd_paddr <= _GEN_1651;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_1_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_1_rob_addr <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h1 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_1_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 316:48]
      end else begin
        buf_1_rob_addr <= _GEN_1635;
      end
    end else begin
      buf_1_rob_addr <= _GEN_1635;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_valid <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_valid <= _GEN_1828;
      end
    end else begin
      buf_2_valid <= _GEN_1828;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_pc <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_pc <= _GEN_1820;
      end
    end else begin
      buf_2_pc <= _GEN_1820;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_fu_code <= 3'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_fu_code <= _GEN_1796;
      end
    end else begin
      buf_2_fu_code <= _GEN_1796;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_alu_code <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_alu_code <= _GEN_1788;
      end
    end else begin
      buf_2_alu_code <= _GEN_1788;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_mem_code <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_mem_code <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_mem_code <= io_in_bits_vec_1_mem_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_mem_code <= _GEN_1772;
      end
    end else begin
      buf_2_mem_code <= _GEN_1772;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_mem_size <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_mem_size <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_mem_size <= io_in_bits_vec_1_mem_size; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_mem_size <= _GEN_1764;
      end
    end else begin
      buf_2_mem_size <= _GEN_1764;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_w_type <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_w_type <= _GEN_1748;
      end
    end else begin
      buf_2_w_type <= _GEN_1748;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_rs1_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_rs1_src <= _GEN_1740;
      end
    end else begin
      buf_2_rs1_src <= _GEN_1740;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_rs2_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_rs2_src <= _GEN_1732;
      end
    end else begin
      buf_2_rs2_src <= _GEN_1732;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_rd_en <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_rd_en <= _GEN_1700;
      end
    end else begin
      buf_2_rd_en <= _GEN_1700;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_imm <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_imm <= _GEN_1692;
      end
    end else begin
      buf_2_imm <= _GEN_1692;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_rs1_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_rs1_paddr <= _GEN_1668;
      end
    end else begin
      buf_2_rs1_paddr <= _GEN_1668;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_rs2_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_rs2_paddr <= _GEN_1660;
      end
    end else begin
      buf_2_rs2_paddr <= _GEN_1660;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_rd_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_rd_paddr <= _GEN_1652;
      end
    end else begin
      buf_2_rd_paddr <= _GEN_1652;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_2_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_2_rob_addr <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h2 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_2_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 316:48]
      end else begin
        buf_2_rob_addr <= _GEN_1636;
      end
    end else begin
      buf_2_rob_addr <= _GEN_1636;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_valid <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_valid <= _GEN_1829;
      end
    end else begin
      buf_3_valid <= _GEN_1829;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_pc <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_pc <= _GEN_1821;
      end
    end else begin
      buf_3_pc <= _GEN_1821;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_fu_code <= 3'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_fu_code <= _GEN_1797;
      end
    end else begin
      buf_3_fu_code <= _GEN_1797;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_alu_code <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_alu_code <= _GEN_1789;
      end
    end else begin
      buf_3_alu_code <= _GEN_1789;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_mem_code <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_mem_code <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_mem_code <= io_in_bits_vec_1_mem_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_mem_code <= _GEN_1773;
      end
    end else begin
      buf_3_mem_code <= _GEN_1773;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_mem_size <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_mem_size <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_mem_size <= io_in_bits_vec_1_mem_size; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_mem_size <= _GEN_1765;
      end
    end else begin
      buf_3_mem_size <= _GEN_1765;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_w_type <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_w_type <= _GEN_1749;
      end
    end else begin
      buf_3_w_type <= _GEN_1749;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_rs1_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_rs1_src <= _GEN_1741;
      end
    end else begin
      buf_3_rs1_src <= _GEN_1741;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_rs2_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_rs2_src <= _GEN_1733;
      end
    end else begin
      buf_3_rs2_src <= _GEN_1733;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_rd_en <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_rd_en <= _GEN_1701;
      end
    end else begin
      buf_3_rd_en <= _GEN_1701;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_imm <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_imm <= _GEN_1693;
      end
    end else begin
      buf_3_imm <= _GEN_1693;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_rs1_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_rs1_paddr <= _GEN_1669;
      end
    end else begin
      buf_3_rs1_paddr <= _GEN_1669;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_rs2_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_rs2_paddr <= _GEN_1661;
      end
    end else begin
      buf_3_rs2_paddr <= _GEN_1661;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_rd_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_rd_paddr <= _GEN_1653;
      end
    end else begin
      buf_3_rd_paddr <= _GEN_1653;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_3_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_3_rob_addr <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h3 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_3_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 316:48]
      end else begin
        buf_3_rob_addr <= _GEN_1637;
      end
    end else begin
      buf_3_rob_addr <= _GEN_1637;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_valid <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_valid <= _GEN_1830;
      end
    end else begin
      buf_4_valid <= _GEN_1830;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_pc <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_pc <= _GEN_1822;
      end
    end else begin
      buf_4_pc <= _GEN_1822;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_fu_code <= 3'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_fu_code <= _GEN_1798;
      end
    end else begin
      buf_4_fu_code <= _GEN_1798;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_alu_code <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_alu_code <= _GEN_1790;
      end
    end else begin
      buf_4_alu_code <= _GEN_1790;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_mem_code <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_mem_code <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_mem_code <= io_in_bits_vec_1_mem_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_mem_code <= _GEN_1774;
      end
    end else begin
      buf_4_mem_code <= _GEN_1774;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_mem_size <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_mem_size <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_mem_size <= io_in_bits_vec_1_mem_size; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_mem_size <= _GEN_1766;
      end
    end else begin
      buf_4_mem_size <= _GEN_1766;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_w_type <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_w_type <= _GEN_1750;
      end
    end else begin
      buf_4_w_type <= _GEN_1750;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_rs1_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_rs1_src <= _GEN_1742;
      end
    end else begin
      buf_4_rs1_src <= _GEN_1742;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_rs2_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_rs2_src <= _GEN_1734;
      end
    end else begin
      buf_4_rs2_src <= _GEN_1734;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_rd_en <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_rd_en <= _GEN_1702;
      end
    end else begin
      buf_4_rd_en <= _GEN_1702;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_imm <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_imm <= _GEN_1694;
      end
    end else begin
      buf_4_imm <= _GEN_1694;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_rs1_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_rs1_paddr <= _GEN_1670;
      end
    end else begin
      buf_4_rs1_paddr <= _GEN_1670;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_rs2_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_rs2_paddr <= _GEN_1662;
      end
    end else begin
      buf_4_rs2_paddr <= _GEN_1662;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_rd_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_rd_paddr <= _GEN_1654;
      end
    end else begin
      buf_4_rd_paddr <= _GEN_1654;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_4_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_4_rob_addr <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h4 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_4_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 316:48]
      end else begin
        buf_4_rob_addr <= _GEN_1638;
      end
    end else begin
      buf_4_rob_addr <= _GEN_1638;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_valid <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_valid <= _GEN_1831;
      end
    end else begin
      buf_5_valid <= _GEN_1831;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_pc <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_pc <= _GEN_1823;
      end
    end else begin
      buf_5_pc <= _GEN_1823;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_fu_code <= 3'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_fu_code <= _GEN_1799;
      end
    end else begin
      buf_5_fu_code <= _GEN_1799;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_alu_code <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_alu_code <= _GEN_1791;
      end
    end else begin
      buf_5_alu_code <= _GEN_1791;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_mem_code <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_mem_code <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_mem_code <= io_in_bits_vec_1_mem_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_mem_code <= _GEN_1775;
      end
    end else begin
      buf_5_mem_code <= _GEN_1775;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_mem_size <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_mem_size <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_mem_size <= io_in_bits_vec_1_mem_size; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_mem_size <= _GEN_1767;
      end
    end else begin
      buf_5_mem_size <= _GEN_1767;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_w_type <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_w_type <= _GEN_1751;
      end
    end else begin
      buf_5_w_type <= _GEN_1751;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_rs1_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_rs1_src <= _GEN_1743;
      end
    end else begin
      buf_5_rs1_src <= _GEN_1743;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_rs2_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_rs2_src <= _GEN_1735;
      end
    end else begin
      buf_5_rs2_src <= _GEN_1735;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_rd_en <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_rd_en <= _GEN_1703;
      end
    end else begin
      buf_5_rd_en <= _GEN_1703;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_imm <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_imm <= _GEN_1695;
      end
    end else begin
      buf_5_imm <= _GEN_1695;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_rs1_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_rs1_paddr <= _GEN_1671;
      end
    end else begin
      buf_5_rs1_paddr <= _GEN_1671;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_rs2_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_rs2_paddr <= _GEN_1663;
      end
    end else begin
      buf_5_rs2_paddr <= _GEN_1663;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_rd_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_rd_paddr <= _GEN_1655;
      end
    end else begin
      buf_5_rd_paddr <= _GEN_1655;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_5_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_5_rob_addr <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h5 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_5_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 316:48]
      end else begin
        buf_5_rob_addr <= _GEN_1639;
      end
    end else begin
      buf_5_rob_addr <= _GEN_1639;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_valid <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_valid <= _GEN_1832;
      end
    end else begin
      buf_6_valid <= _GEN_1832;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_pc <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_pc <= _GEN_1824;
      end
    end else begin
      buf_6_pc <= _GEN_1824;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_fu_code <= 3'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_fu_code <= _GEN_1800;
      end
    end else begin
      buf_6_fu_code <= _GEN_1800;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_alu_code <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_alu_code <= _GEN_1792;
      end
    end else begin
      buf_6_alu_code <= _GEN_1792;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_mem_code <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_mem_code <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_mem_code <= io_in_bits_vec_1_mem_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_mem_code <= _GEN_1776;
      end
    end else begin
      buf_6_mem_code <= _GEN_1776;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_mem_size <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_mem_size <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_mem_size <= io_in_bits_vec_1_mem_size; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_mem_size <= _GEN_1768;
      end
    end else begin
      buf_6_mem_size <= _GEN_1768;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_w_type <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_w_type <= _GEN_1752;
      end
    end else begin
      buf_6_w_type <= _GEN_1752;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_rs1_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_rs1_src <= _GEN_1744;
      end
    end else begin
      buf_6_rs1_src <= _GEN_1744;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_rs2_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_rs2_src <= _GEN_1736;
      end
    end else begin
      buf_6_rs2_src <= _GEN_1736;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_rd_en <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_rd_en <= _GEN_1704;
      end
    end else begin
      buf_6_rd_en <= _GEN_1704;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_imm <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_imm <= _GEN_1696;
      end
    end else begin
      buf_6_imm <= _GEN_1696;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_rs1_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_rs1_paddr <= _GEN_1672;
      end
    end else begin
      buf_6_rs1_paddr <= _GEN_1672;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_rs2_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_rs2_paddr <= _GEN_1664;
      end
    end else begin
      buf_6_rs2_paddr <= _GEN_1664;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_rd_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_rd_paddr <= _GEN_1656;
      end
    end else begin
      buf_6_rd_paddr <= _GEN_1656;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_6_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_6_rob_addr <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h6 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_6_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 316:48]
      end else begin
        buf_6_rob_addr <= _GEN_1640;
      end
    end else begin
      buf_6_rob_addr <= _GEN_1640;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_valid <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_valid <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_valid <= io_in_bits_vec_1_valid; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_valid <= _GEN_1833;
      end
    end else begin
      buf_7_valid <= _GEN_1833;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_pc <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_pc <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_pc <= io_in_bits_vec_1_pc; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_pc <= _GEN_1825;
      end
    end else begin
      buf_7_pc <= _GEN_1825;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_fu_code <= 3'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_fu_code <= 3'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_fu_code <= io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_fu_code <= _GEN_1801;
      end
    end else begin
      buf_7_fu_code <= _GEN_1801;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_alu_code <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_alu_code <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_alu_code <= io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_alu_code <= _GEN_1793;
      end
    end else begin
      buf_7_alu_code <= _GEN_1793;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_mem_code <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_mem_code <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_mem_code <= io_in_bits_vec_1_mem_code; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_mem_code <= _GEN_1777;
      end
    end else begin
      buf_7_mem_code <= _GEN_1777;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_mem_size <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_mem_size <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_mem_size <= io_in_bits_vec_1_mem_size; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_mem_size <= _GEN_1769;
      end
    end else begin
      buf_7_mem_size <= _GEN_1769;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_w_type <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_w_type <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_w_type <= io_in_bits_vec_1_w_type; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_w_type <= _GEN_1753;
      end
    end else begin
      buf_7_w_type <= _GEN_1753;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_rs1_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_rs1_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_rs1_src <= io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_rs1_src <= _GEN_1745;
      end
    end else begin
      buf_7_rs1_src <= _GEN_1745;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_rs2_src <= 2'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_rs2_src <= 2'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_rs2_src <= io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_rs2_src <= _GEN_1737;
      end
    end else begin
      buf_7_rs2_src <= _GEN_1737;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_rd_en <= 1'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_rd_en <= 1'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_rd_en <= io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_rd_en <= _GEN_1705;
      end
    end else begin
      buf_7_rd_en <= _GEN_1705;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_imm <= 32'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_imm <= 32'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_imm <= io_in_bits_vec_1_imm; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_imm <= _GEN_1697;
      end
    end else begin
      buf_7_imm <= _GEN_1697;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_rs1_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_rs1_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_rs1_paddr <= io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_rs1_paddr <= _GEN_1673;
      end
    end else begin
      buf_7_rs1_paddr <= _GEN_1673;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_rs2_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_rs2_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_rs2_paddr <= io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_rs2_paddr <= _GEN_1665;
      end
    end else begin
      buf_7_rs2_paddr <= _GEN_1665;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_rd_paddr <= 6'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_rd_paddr <= 6'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_rd_paddr <= io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_rd_paddr <= _GEN_1657;
      end
    end else begin
      buf_7_rd_paddr <= _GEN_1657;
    end
    if (reset) begin // @[IssueUnit.scala 97:20]
      buf_7_rob_addr <= 4'h0; // @[IssueUnit.scala 97:20]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      buf_7_rob_addr <= 4'h0; // @[IssueUnit.scala 332:14]
    end else if (io_in_bits_vec_1_valid & _T & ~io_flush) begin // @[IssueUnit.scala 315:51]
      if (3'h7 == _GEN_1835[2:0]) begin // @[IssueUnit.scala 316:48]
        buf_7_rob_addr <= io_rob_addr_1; // @[IssueUnit.scala 316:48]
      end else begin
        buf_7_rob_addr <= _GEN_1641;
      end
    end else begin
      buf_7_rob_addr <= _GEN_1641;
    end
    if (reset) begin // @[IssueUnit.scala 102:24]
      enq_vec_0 <= 4'h0; // @[IssueUnit.scala 102:24]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      enq_vec_0 <= 4'h0; // @[IssueUnit.scala 334:13]
    end else if ((_T | (|io_out_0_valid)) & _T_97) begin // @[IssueUnit.scala 322:70]
      enq_vec_0 <= next_enq_vec_0; // @[IssueUnit.scala 323:13]
    end
    if (reset) begin // @[IssueUnit.scala 102:24]
      enq_vec_1 <= 4'h1; // @[IssueUnit.scala 102:24]
    end else if (io_flush) begin // @[IssueUnit.scala 330:19]
      enq_vec_1 <= 4'h1; // @[IssueUnit.scala 334:13]
    end else if ((_T | (|io_out_0_valid)) & _T_97) begin // @[IssueUnit.scala 322:70]
      enq_vec_1 <= next_enq_vec_1; // @[IssueUnit.scala 323:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  buf_0_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  buf_0_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  buf_0_fu_code = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  buf_0_alu_code = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  buf_0_mem_code = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  buf_0_mem_size = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  buf_0_w_type = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  buf_0_rs1_src = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  buf_0_rs2_src = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  buf_0_rd_en = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  buf_0_imm = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  buf_0_rs1_paddr = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  buf_0_rs2_paddr = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  buf_0_rd_paddr = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  buf_0_rob_addr = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  buf_1_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  buf_1_pc = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  buf_1_fu_code = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  buf_1_alu_code = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  buf_1_mem_code = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  buf_1_mem_size = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  buf_1_w_type = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  buf_1_rs1_src = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  buf_1_rs2_src = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  buf_1_rd_en = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  buf_1_imm = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  buf_1_rs1_paddr = _RAND_26[5:0];
  _RAND_27 = {1{`RANDOM}};
  buf_1_rs2_paddr = _RAND_27[5:0];
  _RAND_28 = {1{`RANDOM}};
  buf_1_rd_paddr = _RAND_28[5:0];
  _RAND_29 = {1{`RANDOM}};
  buf_1_rob_addr = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  buf_2_valid = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  buf_2_pc = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  buf_2_fu_code = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  buf_2_alu_code = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  buf_2_mem_code = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  buf_2_mem_size = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  buf_2_w_type = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  buf_2_rs1_src = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  buf_2_rs2_src = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  buf_2_rd_en = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  buf_2_imm = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  buf_2_rs1_paddr = _RAND_41[5:0];
  _RAND_42 = {1{`RANDOM}};
  buf_2_rs2_paddr = _RAND_42[5:0];
  _RAND_43 = {1{`RANDOM}};
  buf_2_rd_paddr = _RAND_43[5:0];
  _RAND_44 = {1{`RANDOM}};
  buf_2_rob_addr = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  buf_3_valid = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  buf_3_pc = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  buf_3_fu_code = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  buf_3_alu_code = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  buf_3_mem_code = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  buf_3_mem_size = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  buf_3_w_type = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  buf_3_rs1_src = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  buf_3_rs2_src = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  buf_3_rd_en = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  buf_3_imm = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  buf_3_rs1_paddr = _RAND_56[5:0];
  _RAND_57 = {1{`RANDOM}};
  buf_3_rs2_paddr = _RAND_57[5:0];
  _RAND_58 = {1{`RANDOM}};
  buf_3_rd_paddr = _RAND_58[5:0];
  _RAND_59 = {1{`RANDOM}};
  buf_3_rob_addr = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  buf_4_valid = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  buf_4_pc = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  buf_4_fu_code = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  buf_4_alu_code = _RAND_63[3:0];
  _RAND_64 = {1{`RANDOM}};
  buf_4_mem_code = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  buf_4_mem_size = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  buf_4_w_type = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  buf_4_rs1_src = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  buf_4_rs2_src = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  buf_4_rd_en = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  buf_4_imm = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  buf_4_rs1_paddr = _RAND_71[5:0];
  _RAND_72 = {1{`RANDOM}};
  buf_4_rs2_paddr = _RAND_72[5:0];
  _RAND_73 = {1{`RANDOM}};
  buf_4_rd_paddr = _RAND_73[5:0];
  _RAND_74 = {1{`RANDOM}};
  buf_4_rob_addr = _RAND_74[3:0];
  _RAND_75 = {1{`RANDOM}};
  buf_5_valid = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  buf_5_pc = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  buf_5_fu_code = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  buf_5_alu_code = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  buf_5_mem_code = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  buf_5_mem_size = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  buf_5_w_type = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  buf_5_rs1_src = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  buf_5_rs2_src = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  buf_5_rd_en = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  buf_5_imm = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  buf_5_rs1_paddr = _RAND_86[5:0];
  _RAND_87 = {1{`RANDOM}};
  buf_5_rs2_paddr = _RAND_87[5:0];
  _RAND_88 = {1{`RANDOM}};
  buf_5_rd_paddr = _RAND_88[5:0];
  _RAND_89 = {1{`RANDOM}};
  buf_5_rob_addr = _RAND_89[3:0];
  _RAND_90 = {1{`RANDOM}};
  buf_6_valid = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  buf_6_pc = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  buf_6_fu_code = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  buf_6_alu_code = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  buf_6_mem_code = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  buf_6_mem_size = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  buf_6_w_type = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  buf_6_rs1_src = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  buf_6_rs2_src = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  buf_6_rd_en = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  buf_6_imm = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  buf_6_rs1_paddr = _RAND_101[5:0];
  _RAND_102 = {1{`RANDOM}};
  buf_6_rs2_paddr = _RAND_102[5:0];
  _RAND_103 = {1{`RANDOM}};
  buf_6_rd_paddr = _RAND_103[5:0];
  _RAND_104 = {1{`RANDOM}};
  buf_6_rob_addr = _RAND_104[3:0];
  _RAND_105 = {1{`RANDOM}};
  buf_7_valid = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  buf_7_pc = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  buf_7_fu_code = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  buf_7_alu_code = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  buf_7_mem_code = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  buf_7_mem_size = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  buf_7_w_type = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  buf_7_rs1_src = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  buf_7_rs2_src = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  buf_7_rd_en = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  buf_7_imm = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  buf_7_rs1_paddr = _RAND_116[5:0];
  _RAND_117 = {1{`RANDOM}};
  buf_7_rs2_paddr = _RAND_117[5:0];
  _RAND_118 = {1{`RANDOM}};
  buf_7_rd_paddr = _RAND_118[5:0];
  _RAND_119 = {1{`RANDOM}};
  buf_7_rob_addr = _RAND_119[3:0];
  _RAND_120 = {1{`RANDOM}};
  enq_vec_0 = _RAND_120[3:0];
  _RAND_121 = {1{`RANDOM}};
  enq_vec_1 = _RAND_121[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_IssueUnit(
  input         clock,
  input         reset,
  input         io_flush,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_vec_0_valid,
  input  [31:0] io_in_bits_vec_0_pc,
  input  [31:0] io_in_bits_vec_0_npc,
  input  [31:0] io_in_bits_vec_0_inst,
  input  [2:0]  io_in_bits_vec_0_fu_code,
  input  [3:0]  io_in_bits_vec_0_alu_code,
  input  [3:0]  io_in_bits_vec_0_jmp_code,
  input  [1:0]  io_in_bits_vec_0_mem_code,
  input  [1:0]  io_in_bits_vec_0_mem_size,
  input  [2:0]  io_in_bits_vec_0_sys_code,
  input         io_in_bits_vec_0_w_type,
  input  [1:0]  io_in_bits_vec_0_rs1_src,
  input  [1:0]  io_in_bits_vec_0_rs2_src,
  input         io_in_bits_vec_0_rd_en,
  input  [31:0] io_in_bits_vec_0_imm,
  input         io_in_bits_vec_0_pred_br,
  input  [31:0] io_in_bits_vec_0_pred_bpc,
  input  [5:0]  io_in_bits_vec_0_rs1_paddr,
  input  [5:0]  io_in_bits_vec_0_rs2_paddr,
  input  [5:0]  io_in_bits_vec_0_rd_paddr,
  input         io_in_bits_vec_1_valid,
  input  [31:0] io_in_bits_vec_1_pc,
  input  [31:0] io_in_bits_vec_1_npc,
  input  [31:0] io_in_bits_vec_1_inst,
  input  [2:0]  io_in_bits_vec_1_fu_code,
  input  [3:0]  io_in_bits_vec_1_alu_code,
  input  [3:0]  io_in_bits_vec_1_jmp_code,
  input  [1:0]  io_in_bits_vec_1_mem_code,
  input  [1:0]  io_in_bits_vec_1_mem_size,
  input  [2:0]  io_in_bits_vec_1_sys_code,
  input         io_in_bits_vec_1_w_type,
  input  [1:0]  io_in_bits_vec_1_rs1_src,
  input  [1:0]  io_in_bits_vec_1_rs2_src,
  input         io_in_bits_vec_1_rd_en,
  input  [31:0] io_in_bits_vec_1_imm,
  input         io_in_bits_vec_1_pred_br,
  input  [31:0] io_in_bits_vec_1_pred_bpc,
  input  [5:0]  io_in_bits_vec_1_rs1_paddr,
  input  [5:0]  io_in_bits_vec_1_rs2_paddr,
  input  [5:0]  io_in_bits_vec_1_rd_paddr,
  input  [3:0]  io_rob_addr_0,
  input  [3:0]  io_rob_addr_1,
  output        io_out_0_valid,
  output [31:0] io_out_0_pc,
  output [31:0] io_out_0_npc,
  output [31:0] io_out_0_inst,
  output [2:0]  io_out_0_fu_code,
  output [3:0]  io_out_0_alu_code,
  output [3:0]  io_out_0_jmp_code,
  output [2:0]  io_out_0_sys_code,
  output        io_out_0_w_type,
  output [1:0]  io_out_0_rs1_src,
  output [1:0]  io_out_0_rs2_src,
  output        io_out_0_rd_en,
  output [31:0] io_out_0_imm,
  output        io_out_0_pred_br,
  output [31:0] io_out_0_pred_bpc,
  output [5:0]  io_out_0_rs1_paddr,
  output [5:0]  io_out_0_rs2_paddr,
  output [5:0]  io_out_0_rd_paddr,
  output [3:0]  io_out_0_rob_addr,
  output        io_out_1_valid,
  output [31:0] io_out_1_pc,
  output [31:0] io_out_1_npc,
  output [2:0]  io_out_1_fu_code,
  output [3:0]  io_out_1_alu_code,
  output [3:0]  io_out_1_jmp_code,
  output        io_out_1_w_type,
  output [1:0]  io_out_1_rs1_src,
  output [1:0]  io_out_1_rs2_src,
  output        io_out_1_rd_en,
  output [31:0] io_out_1_imm,
  output        io_out_1_pred_br,
  output [31:0] io_out_1_pred_bpc,
  output [5:0]  io_out_1_rs1_paddr,
  output [5:0]  io_out_1_rs2_paddr,
  output [5:0]  io_out_1_rd_paddr,
  output [3:0]  io_out_1_rob_addr,
  output        io_out_2_valid,
  output [31:0] io_out_2_pc,
  output [2:0]  io_out_2_fu_code,
  output [3:0]  io_out_2_alu_code,
  output [1:0]  io_out_2_mem_code,
  output [1:0]  io_out_2_mem_size,
  output        io_out_2_w_type,
  output [1:0]  io_out_2_rs1_src,
  output [1:0]  io_out_2_rs2_src,
  output        io_out_2_rd_en,
  output [31:0] io_out_2_imm,
  output [5:0]  io_out_2_rs1_paddr,
  output [5:0]  io_out_2_rs2_paddr,
  output [5:0]  io_out_2_rd_paddr,
  output [3:0]  io_out_2_rob_addr,
  input  [63:0] io_avail_list,
  input         io_lsu_ready,
  input         io_sys_ready
);
  wire  int_iq_clock; // @[IssueUnit.scala 24:22]
  wire  int_iq_reset; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_flush; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_in_ready; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_in_valid; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_in_bits_vec_0_valid; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_in_bits_vec_0_pc; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_in_bits_vec_0_npc; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_in_bits_vec_0_inst; // @[IssueUnit.scala 24:22]
  wire [2:0] int_iq_io_in_bits_vec_0_fu_code; // @[IssueUnit.scala 24:22]
  wire [3:0] int_iq_io_in_bits_vec_0_alu_code; // @[IssueUnit.scala 24:22]
  wire [3:0] int_iq_io_in_bits_vec_0_jmp_code; // @[IssueUnit.scala 24:22]
  wire [2:0] int_iq_io_in_bits_vec_0_sys_code; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_in_bits_vec_0_w_type; // @[IssueUnit.scala 24:22]
  wire [1:0] int_iq_io_in_bits_vec_0_rs1_src; // @[IssueUnit.scala 24:22]
  wire [1:0] int_iq_io_in_bits_vec_0_rs2_src; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_in_bits_vec_0_rd_en; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_in_bits_vec_0_imm; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_in_bits_vec_0_pred_br; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_in_bits_vec_0_pred_bpc; // @[IssueUnit.scala 24:22]
  wire [5:0] int_iq_io_in_bits_vec_0_rs1_paddr; // @[IssueUnit.scala 24:22]
  wire [5:0] int_iq_io_in_bits_vec_0_rs2_paddr; // @[IssueUnit.scala 24:22]
  wire [5:0] int_iq_io_in_bits_vec_0_rd_paddr; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_in_bits_vec_1_valid; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_in_bits_vec_1_pc; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_in_bits_vec_1_npc; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_in_bits_vec_1_inst; // @[IssueUnit.scala 24:22]
  wire [2:0] int_iq_io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 24:22]
  wire [3:0] int_iq_io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 24:22]
  wire [3:0] int_iq_io_in_bits_vec_1_jmp_code; // @[IssueUnit.scala 24:22]
  wire [2:0] int_iq_io_in_bits_vec_1_sys_code; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_in_bits_vec_1_w_type; // @[IssueUnit.scala 24:22]
  wire [1:0] int_iq_io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 24:22]
  wire [1:0] int_iq_io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_in_bits_vec_1_imm; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_in_bits_vec_1_pred_br; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_in_bits_vec_1_pred_bpc; // @[IssueUnit.scala 24:22]
  wire [5:0] int_iq_io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 24:22]
  wire [5:0] int_iq_io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 24:22]
  wire [5:0] int_iq_io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 24:22]
  wire [3:0] int_iq_io_rob_addr_0; // @[IssueUnit.scala 24:22]
  wire [3:0] int_iq_io_rob_addr_1; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_out_0_valid; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_out_0_pc; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_out_0_npc; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_out_0_inst; // @[IssueUnit.scala 24:22]
  wire [2:0] int_iq_io_out_0_fu_code; // @[IssueUnit.scala 24:22]
  wire [3:0] int_iq_io_out_0_alu_code; // @[IssueUnit.scala 24:22]
  wire [3:0] int_iq_io_out_0_jmp_code; // @[IssueUnit.scala 24:22]
  wire [2:0] int_iq_io_out_0_sys_code; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_out_0_w_type; // @[IssueUnit.scala 24:22]
  wire [1:0] int_iq_io_out_0_rs1_src; // @[IssueUnit.scala 24:22]
  wire [1:0] int_iq_io_out_0_rs2_src; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_out_0_rd_en; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_out_0_imm; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_out_0_pred_br; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_out_0_pred_bpc; // @[IssueUnit.scala 24:22]
  wire [5:0] int_iq_io_out_0_rs1_paddr; // @[IssueUnit.scala 24:22]
  wire [5:0] int_iq_io_out_0_rs2_paddr; // @[IssueUnit.scala 24:22]
  wire [5:0] int_iq_io_out_0_rd_paddr; // @[IssueUnit.scala 24:22]
  wire [3:0] int_iq_io_out_0_rob_addr; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_out_1_valid; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_out_1_pc; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_out_1_npc; // @[IssueUnit.scala 24:22]
  wire [2:0] int_iq_io_out_1_fu_code; // @[IssueUnit.scala 24:22]
  wire [3:0] int_iq_io_out_1_alu_code; // @[IssueUnit.scala 24:22]
  wire [3:0] int_iq_io_out_1_jmp_code; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_out_1_w_type; // @[IssueUnit.scala 24:22]
  wire [1:0] int_iq_io_out_1_rs1_src; // @[IssueUnit.scala 24:22]
  wire [1:0] int_iq_io_out_1_rs2_src; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_out_1_rd_en; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_out_1_imm; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_out_1_pred_br; // @[IssueUnit.scala 24:22]
  wire [31:0] int_iq_io_out_1_pred_bpc; // @[IssueUnit.scala 24:22]
  wire [5:0] int_iq_io_out_1_rs1_paddr; // @[IssueUnit.scala 24:22]
  wire [5:0] int_iq_io_out_1_rs2_paddr; // @[IssueUnit.scala 24:22]
  wire [5:0] int_iq_io_out_1_rd_paddr; // @[IssueUnit.scala 24:22]
  wire [3:0] int_iq_io_out_1_rob_addr; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_0; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_1; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_2; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_3; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_4; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_5; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_6; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_7; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_8; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_9; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_10; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_11; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_12; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_13; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_14; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_15; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_16; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_17; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_18; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_19; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_20; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_21; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_22; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_23; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_24; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_25; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_26; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_27; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_28; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_29; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_30; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_31; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_32; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_33; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_34; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_35; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_36; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_37; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_38; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_39; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_40; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_41; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_42; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_43; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_44; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_45; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_46; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_47; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_48; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_49; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_50; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_51; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_52; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_53; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_54; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_55; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_56; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_57; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_58; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_59; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_60; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_61; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_62; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_avail_list_63; // @[IssueUnit.scala 24:22]
  wire  int_iq_io_sys_ready; // @[IssueUnit.scala 24:22]
  wire  mem_iq_clock; // @[IssueUnit.scala 32:22]
  wire  mem_iq_reset; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_flush; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_in_ready; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_in_valid; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_in_bits_vec_0_valid; // @[IssueUnit.scala 32:22]
  wire [31:0] mem_iq_io_in_bits_vec_0_pc; // @[IssueUnit.scala 32:22]
  wire [2:0] mem_iq_io_in_bits_vec_0_fu_code; // @[IssueUnit.scala 32:22]
  wire [3:0] mem_iq_io_in_bits_vec_0_alu_code; // @[IssueUnit.scala 32:22]
  wire [1:0] mem_iq_io_in_bits_vec_0_mem_code; // @[IssueUnit.scala 32:22]
  wire [1:0] mem_iq_io_in_bits_vec_0_mem_size; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_in_bits_vec_0_w_type; // @[IssueUnit.scala 32:22]
  wire [1:0] mem_iq_io_in_bits_vec_0_rs1_src; // @[IssueUnit.scala 32:22]
  wire [1:0] mem_iq_io_in_bits_vec_0_rs2_src; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_in_bits_vec_0_rd_en; // @[IssueUnit.scala 32:22]
  wire [31:0] mem_iq_io_in_bits_vec_0_imm; // @[IssueUnit.scala 32:22]
  wire [5:0] mem_iq_io_in_bits_vec_0_rs1_paddr; // @[IssueUnit.scala 32:22]
  wire [5:0] mem_iq_io_in_bits_vec_0_rs2_paddr; // @[IssueUnit.scala 32:22]
  wire [5:0] mem_iq_io_in_bits_vec_0_rd_paddr; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_in_bits_vec_1_valid; // @[IssueUnit.scala 32:22]
  wire [31:0] mem_iq_io_in_bits_vec_1_pc; // @[IssueUnit.scala 32:22]
  wire [2:0] mem_iq_io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 32:22]
  wire [3:0] mem_iq_io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 32:22]
  wire [1:0] mem_iq_io_in_bits_vec_1_mem_code; // @[IssueUnit.scala 32:22]
  wire [1:0] mem_iq_io_in_bits_vec_1_mem_size; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_in_bits_vec_1_w_type; // @[IssueUnit.scala 32:22]
  wire [1:0] mem_iq_io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 32:22]
  wire [1:0] mem_iq_io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 32:22]
  wire [31:0] mem_iq_io_in_bits_vec_1_imm; // @[IssueUnit.scala 32:22]
  wire [5:0] mem_iq_io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 32:22]
  wire [5:0] mem_iq_io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 32:22]
  wire [5:0] mem_iq_io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 32:22]
  wire [3:0] mem_iq_io_rob_addr_0; // @[IssueUnit.scala 32:22]
  wire [3:0] mem_iq_io_rob_addr_1; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_out_0_valid; // @[IssueUnit.scala 32:22]
  wire [31:0] mem_iq_io_out_0_pc; // @[IssueUnit.scala 32:22]
  wire [2:0] mem_iq_io_out_0_fu_code; // @[IssueUnit.scala 32:22]
  wire [3:0] mem_iq_io_out_0_alu_code; // @[IssueUnit.scala 32:22]
  wire [1:0] mem_iq_io_out_0_mem_code; // @[IssueUnit.scala 32:22]
  wire [1:0] mem_iq_io_out_0_mem_size; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_out_0_w_type; // @[IssueUnit.scala 32:22]
  wire [1:0] mem_iq_io_out_0_rs1_src; // @[IssueUnit.scala 32:22]
  wire [1:0] mem_iq_io_out_0_rs2_src; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_out_0_rd_en; // @[IssueUnit.scala 32:22]
  wire [31:0] mem_iq_io_out_0_imm; // @[IssueUnit.scala 32:22]
  wire [5:0] mem_iq_io_out_0_rs1_paddr; // @[IssueUnit.scala 32:22]
  wire [5:0] mem_iq_io_out_0_rs2_paddr; // @[IssueUnit.scala 32:22]
  wire [5:0] mem_iq_io_out_0_rd_paddr; // @[IssueUnit.scala 32:22]
  wire [3:0] mem_iq_io_out_0_rob_addr; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_0; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_1; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_2; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_3; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_4; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_5; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_6; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_7; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_8; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_9; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_10; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_11; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_12; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_13; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_14; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_15; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_16; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_17; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_18; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_19; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_20; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_21; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_22; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_23; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_24; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_25; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_26; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_27; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_28; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_29; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_30; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_31; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_32; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_33; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_34; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_35; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_36; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_37; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_38; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_39; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_40; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_41; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_42; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_43; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_44; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_45; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_46; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_47; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_48; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_49; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_50; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_51; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_52; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_53; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_54; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_55; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_56; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_57; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_58; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_59; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_60; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_61; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_62; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_avail_list_63; // @[IssueUnit.scala 32:22]
  wire  mem_iq_io_fu_ready; // @[IssueUnit.scala 32:22]
  wire  uop_int_0_valid = io_in_bits_vec_0_fu_code == 3'h4 ? 1'h0 : io_in_bits_vec_0_valid; // @[IssueUnit.scala 44:11 48:49 49:24]
  wire  uop_mem_0_valid = io_in_bits_vec_0_fu_code != 3'h4 ? 1'h0 : io_in_bits_vec_0_valid; // @[IssueUnit.scala 45:11 51:49 52:24]
  wire  uop_int_1_valid = io_in_bits_vec_1_fu_code == 3'h4 ? 1'h0 : io_in_bits_vec_1_valid; // @[IssueUnit.scala 44:11 48:49 49:24]
  wire  uop_mem_1_valid = io_in_bits_vec_1_fu_code != 3'h4 ? 1'h0 : io_in_bits_vec_1_valid; // @[IssueUnit.scala 45:11 51:49 52:24]
  wire [1:0] _T_260 = {uop_int_0_valid,uop_int_1_valid}; // @[Cat.scala 30:58]
  wire [1:0] _T_264 = {uop_mem_0_valid,uop_mem_1_valid}; // @[Cat.scala 30:58]
  ysyx_210128_IntIssueQueueOutOfOrder int_iq ( // @[IssueUnit.scala 24:22]
    .clock(int_iq_clock),
    .reset(int_iq_reset),
    .io_flush(int_iq_io_flush),
    .io_in_ready(int_iq_io_in_ready),
    .io_in_valid(int_iq_io_in_valid),
    .io_in_bits_vec_0_valid(int_iq_io_in_bits_vec_0_valid),
    .io_in_bits_vec_0_pc(int_iq_io_in_bits_vec_0_pc),
    .io_in_bits_vec_0_npc(int_iq_io_in_bits_vec_0_npc),
    .io_in_bits_vec_0_inst(int_iq_io_in_bits_vec_0_inst),
    .io_in_bits_vec_0_fu_code(int_iq_io_in_bits_vec_0_fu_code),
    .io_in_bits_vec_0_alu_code(int_iq_io_in_bits_vec_0_alu_code),
    .io_in_bits_vec_0_jmp_code(int_iq_io_in_bits_vec_0_jmp_code),
    .io_in_bits_vec_0_sys_code(int_iq_io_in_bits_vec_0_sys_code),
    .io_in_bits_vec_0_w_type(int_iq_io_in_bits_vec_0_w_type),
    .io_in_bits_vec_0_rs1_src(int_iq_io_in_bits_vec_0_rs1_src),
    .io_in_bits_vec_0_rs2_src(int_iq_io_in_bits_vec_0_rs2_src),
    .io_in_bits_vec_0_rd_en(int_iq_io_in_bits_vec_0_rd_en),
    .io_in_bits_vec_0_imm(int_iq_io_in_bits_vec_0_imm),
    .io_in_bits_vec_0_pred_br(int_iq_io_in_bits_vec_0_pred_br),
    .io_in_bits_vec_0_pred_bpc(int_iq_io_in_bits_vec_0_pred_bpc),
    .io_in_bits_vec_0_rs1_paddr(int_iq_io_in_bits_vec_0_rs1_paddr),
    .io_in_bits_vec_0_rs2_paddr(int_iq_io_in_bits_vec_0_rs2_paddr),
    .io_in_bits_vec_0_rd_paddr(int_iq_io_in_bits_vec_0_rd_paddr),
    .io_in_bits_vec_1_valid(int_iq_io_in_bits_vec_1_valid),
    .io_in_bits_vec_1_pc(int_iq_io_in_bits_vec_1_pc),
    .io_in_bits_vec_1_npc(int_iq_io_in_bits_vec_1_npc),
    .io_in_bits_vec_1_inst(int_iq_io_in_bits_vec_1_inst),
    .io_in_bits_vec_1_fu_code(int_iq_io_in_bits_vec_1_fu_code),
    .io_in_bits_vec_1_alu_code(int_iq_io_in_bits_vec_1_alu_code),
    .io_in_bits_vec_1_jmp_code(int_iq_io_in_bits_vec_1_jmp_code),
    .io_in_bits_vec_1_sys_code(int_iq_io_in_bits_vec_1_sys_code),
    .io_in_bits_vec_1_w_type(int_iq_io_in_bits_vec_1_w_type),
    .io_in_bits_vec_1_rs1_src(int_iq_io_in_bits_vec_1_rs1_src),
    .io_in_bits_vec_1_rs2_src(int_iq_io_in_bits_vec_1_rs2_src),
    .io_in_bits_vec_1_rd_en(int_iq_io_in_bits_vec_1_rd_en),
    .io_in_bits_vec_1_imm(int_iq_io_in_bits_vec_1_imm),
    .io_in_bits_vec_1_pred_br(int_iq_io_in_bits_vec_1_pred_br),
    .io_in_bits_vec_1_pred_bpc(int_iq_io_in_bits_vec_1_pred_bpc),
    .io_in_bits_vec_1_rs1_paddr(int_iq_io_in_bits_vec_1_rs1_paddr),
    .io_in_bits_vec_1_rs2_paddr(int_iq_io_in_bits_vec_1_rs2_paddr),
    .io_in_bits_vec_1_rd_paddr(int_iq_io_in_bits_vec_1_rd_paddr),
    .io_rob_addr_0(int_iq_io_rob_addr_0),
    .io_rob_addr_1(int_iq_io_rob_addr_1),
    .io_out_0_valid(int_iq_io_out_0_valid),
    .io_out_0_pc(int_iq_io_out_0_pc),
    .io_out_0_npc(int_iq_io_out_0_npc),
    .io_out_0_inst(int_iq_io_out_0_inst),
    .io_out_0_fu_code(int_iq_io_out_0_fu_code),
    .io_out_0_alu_code(int_iq_io_out_0_alu_code),
    .io_out_0_jmp_code(int_iq_io_out_0_jmp_code),
    .io_out_0_sys_code(int_iq_io_out_0_sys_code),
    .io_out_0_w_type(int_iq_io_out_0_w_type),
    .io_out_0_rs1_src(int_iq_io_out_0_rs1_src),
    .io_out_0_rs2_src(int_iq_io_out_0_rs2_src),
    .io_out_0_rd_en(int_iq_io_out_0_rd_en),
    .io_out_0_imm(int_iq_io_out_0_imm),
    .io_out_0_pred_br(int_iq_io_out_0_pred_br),
    .io_out_0_pred_bpc(int_iq_io_out_0_pred_bpc),
    .io_out_0_rs1_paddr(int_iq_io_out_0_rs1_paddr),
    .io_out_0_rs2_paddr(int_iq_io_out_0_rs2_paddr),
    .io_out_0_rd_paddr(int_iq_io_out_0_rd_paddr),
    .io_out_0_rob_addr(int_iq_io_out_0_rob_addr),
    .io_out_1_valid(int_iq_io_out_1_valid),
    .io_out_1_pc(int_iq_io_out_1_pc),
    .io_out_1_npc(int_iq_io_out_1_npc),
    .io_out_1_fu_code(int_iq_io_out_1_fu_code),
    .io_out_1_alu_code(int_iq_io_out_1_alu_code),
    .io_out_1_jmp_code(int_iq_io_out_1_jmp_code),
    .io_out_1_w_type(int_iq_io_out_1_w_type),
    .io_out_1_rs1_src(int_iq_io_out_1_rs1_src),
    .io_out_1_rs2_src(int_iq_io_out_1_rs2_src),
    .io_out_1_rd_en(int_iq_io_out_1_rd_en),
    .io_out_1_imm(int_iq_io_out_1_imm),
    .io_out_1_pred_br(int_iq_io_out_1_pred_br),
    .io_out_1_pred_bpc(int_iq_io_out_1_pred_bpc),
    .io_out_1_rs1_paddr(int_iq_io_out_1_rs1_paddr),
    .io_out_1_rs2_paddr(int_iq_io_out_1_rs2_paddr),
    .io_out_1_rd_paddr(int_iq_io_out_1_rd_paddr),
    .io_out_1_rob_addr(int_iq_io_out_1_rob_addr),
    .io_avail_list_0(int_iq_io_avail_list_0),
    .io_avail_list_1(int_iq_io_avail_list_1),
    .io_avail_list_2(int_iq_io_avail_list_2),
    .io_avail_list_3(int_iq_io_avail_list_3),
    .io_avail_list_4(int_iq_io_avail_list_4),
    .io_avail_list_5(int_iq_io_avail_list_5),
    .io_avail_list_6(int_iq_io_avail_list_6),
    .io_avail_list_7(int_iq_io_avail_list_7),
    .io_avail_list_8(int_iq_io_avail_list_8),
    .io_avail_list_9(int_iq_io_avail_list_9),
    .io_avail_list_10(int_iq_io_avail_list_10),
    .io_avail_list_11(int_iq_io_avail_list_11),
    .io_avail_list_12(int_iq_io_avail_list_12),
    .io_avail_list_13(int_iq_io_avail_list_13),
    .io_avail_list_14(int_iq_io_avail_list_14),
    .io_avail_list_15(int_iq_io_avail_list_15),
    .io_avail_list_16(int_iq_io_avail_list_16),
    .io_avail_list_17(int_iq_io_avail_list_17),
    .io_avail_list_18(int_iq_io_avail_list_18),
    .io_avail_list_19(int_iq_io_avail_list_19),
    .io_avail_list_20(int_iq_io_avail_list_20),
    .io_avail_list_21(int_iq_io_avail_list_21),
    .io_avail_list_22(int_iq_io_avail_list_22),
    .io_avail_list_23(int_iq_io_avail_list_23),
    .io_avail_list_24(int_iq_io_avail_list_24),
    .io_avail_list_25(int_iq_io_avail_list_25),
    .io_avail_list_26(int_iq_io_avail_list_26),
    .io_avail_list_27(int_iq_io_avail_list_27),
    .io_avail_list_28(int_iq_io_avail_list_28),
    .io_avail_list_29(int_iq_io_avail_list_29),
    .io_avail_list_30(int_iq_io_avail_list_30),
    .io_avail_list_31(int_iq_io_avail_list_31),
    .io_avail_list_32(int_iq_io_avail_list_32),
    .io_avail_list_33(int_iq_io_avail_list_33),
    .io_avail_list_34(int_iq_io_avail_list_34),
    .io_avail_list_35(int_iq_io_avail_list_35),
    .io_avail_list_36(int_iq_io_avail_list_36),
    .io_avail_list_37(int_iq_io_avail_list_37),
    .io_avail_list_38(int_iq_io_avail_list_38),
    .io_avail_list_39(int_iq_io_avail_list_39),
    .io_avail_list_40(int_iq_io_avail_list_40),
    .io_avail_list_41(int_iq_io_avail_list_41),
    .io_avail_list_42(int_iq_io_avail_list_42),
    .io_avail_list_43(int_iq_io_avail_list_43),
    .io_avail_list_44(int_iq_io_avail_list_44),
    .io_avail_list_45(int_iq_io_avail_list_45),
    .io_avail_list_46(int_iq_io_avail_list_46),
    .io_avail_list_47(int_iq_io_avail_list_47),
    .io_avail_list_48(int_iq_io_avail_list_48),
    .io_avail_list_49(int_iq_io_avail_list_49),
    .io_avail_list_50(int_iq_io_avail_list_50),
    .io_avail_list_51(int_iq_io_avail_list_51),
    .io_avail_list_52(int_iq_io_avail_list_52),
    .io_avail_list_53(int_iq_io_avail_list_53),
    .io_avail_list_54(int_iq_io_avail_list_54),
    .io_avail_list_55(int_iq_io_avail_list_55),
    .io_avail_list_56(int_iq_io_avail_list_56),
    .io_avail_list_57(int_iq_io_avail_list_57),
    .io_avail_list_58(int_iq_io_avail_list_58),
    .io_avail_list_59(int_iq_io_avail_list_59),
    .io_avail_list_60(int_iq_io_avail_list_60),
    .io_avail_list_61(int_iq_io_avail_list_61),
    .io_avail_list_62(int_iq_io_avail_list_62),
    .io_avail_list_63(int_iq_io_avail_list_63),
    .io_sys_ready(int_iq_io_sys_ready)
  );
  ysyx_210128_MemIssueQueueOutOfOrder mem_iq ( // @[IssueUnit.scala 32:22]
    .clock(mem_iq_clock),
    .reset(mem_iq_reset),
    .io_flush(mem_iq_io_flush),
    .io_in_ready(mem_iq_io_in_ready),
    .io_in_valid(mem_iq_io_in_valid),
    .io_in_bits_vec_0_valid(mem_iq_io_in_bits_vec_0_valid),
    .io_in_bits_vec_0_pc(mem_iq_io_in_bits_vec_0_pc),
    .io_in_bits_vec_0_fu_code(mem_iq_io_in_bits_vec_0_fu_code),
    .io_in_bits_vec_0_alu_code(mem_iq_io_in_bits_vec_0_alu_code),
    .io_in_bits_vec_0_mem_code(mem_iq_io_in_bits_vec_0_mem_code),
    .io_in_bits_vec_0_mem_size(mem_iq_io_in_bits_vec_0_mem_size),
    .io_in_bits_vec_0_w_type(mem_iq_io_in_bits_vec_0_w_type),
    .io_in_bits_vec_0_rs1_src(mem_iq_io_in_bits_vec_0_rs1_src),
    .io_in_bits_vec_0_rs2_src(mem_iq_io_in_bits_vec_0_rs2_src),
    .io_in_bits_vec_0_rd_en(mem_iq_io_in_bits_vec_0_rd_en),
    .io_in_bits_vec_0_imm(mem_iq_io_in_bits_vec_0_imm),
    .io_in_bits_vec_0_rs1_paddr(mem_iq_io_in_bits_vec_0_rs1_paddr),
    .io_in_bits_vec_0_rs2_paddr(mem_iq_io_in_bits_vec_0_rs2_paddr),
    .io_in_bits_vec_0_rd_paddr(mem_iq_io_in_bits_vec_0_rd_paddr),
    .io_in_bits_vec_1_valid(mem_iq_io_in_bits_vec_1_valid),
    .io_in_bits_vec_1_pc(mem_iq_io_in_bits_vec_1_pc),
    .io_in_bits_vec_1_fu_code(mem_iq_io_in_bits_vec_1_fu_code),
    .io_in_bits_vec_1_alu_code(mem_iq_io_in_bits_vec_1_alu_code),
    .io_in_bits_vec_1_mem_code(mem_iq_io_in_bits_vec_1_mem_code),
    .io_in_bits_vec_1_mem_size(mem_iq_io_in_bits_vec_1_mem_size),
    .io_in_bits_vec_1_w_type(mem_iq_io_in_bits_vec_1_w_type),
    .io_in_bits_vec_1_rs1_src(mem_iq_io_in_bits_vec_1_rs1_src),
    .io_in_bits_vec_1_rs2_src(mem_iq_io_in_bits_vec_1_rs2_src),
    .io_in_bits_vec_1_rd_en(mem_iq_io_in_bits_vec_1_rd_en),
    .io_in_bits_vec_1_imm(mem_iq_io_in_bits_vec_1_imm),
    .io_in_bits_vec_1_rs1_paddr(mem_iq_io_in_bits_vec_1_rs1_paddr),
    .io_in_bits_vec_1_rs2_paddr(mem_iq_io_in_bits_vec_1_rs2_paddr),
    .io_in_bits_vec_1_rd_paddr(mem_iq_io_in_bits_vec_1_rd_paddr),
    .io_rob_addr_0(mem_iq_io_rob_addr_0),
    .io_rob_addr_1(mem_iq_io_rob_addr_1),
    .io_out_0_valid(mem_iq_io_out_0_valid),
    .io_out_0_pc(mem_iq_io_out_0_pc),
    .io_out_0_fu_code(mem_iq_io_out_0_fu_code),
    .io_out_0_alu_code(mem_iq_io_out_0_alu_code),
    .io_out_0_mem_code(mem_iq_io_out_0_mem_code),
    .io_out_0_mem_size(mem_iq_io_out_0_mem_size),
    .io_out_0_w_type(mem_iq_io_out_0_w_type),
    .io_out_0_rs1_src(mem_iq_io_out_0_rs1_src),
    .io_out_0_rs2_src(mem_iq_io_out_0_rs2_src),
    .io_out_0_rd_en(mem_iq_io_out_0_rd_en),
    .io_out_0_imm(mem_iq_io_out_0_imm),
    .io_out_0_rs1_paddr(mem_iq_io_out_0_rs1_paddr),
    .io_out_0_rs2_paddr(mem_iq_io_out_0_rs2_paddr),
    .io_out_0_rd_paddr(mem_iq_io_out_0_rd_paddr),
    .io_out_0_rob_addr(mem_iq_io_out_0_rob_addr),
    .io_avail_list_0(mem_iq_io_avail_list_0),
    .io_avail_list_1(mem_iq_io_avail_list_1),
    .io_avail_list_2(mem_iq_io_avail_list_2),
    .io_avail_list_3(mem_iq_io_avail_list_3),
    .io_avail_list_4(mem_iq_io_avail_list_4),
    .io_avail_list_5(mem_iq_io_avail_list_5),
    .io_avail_list_6(mem_iq_io_avail_list_6),
    .io_avail_list_7(mem_iq_io_avail_list_7),
    .io_avail_list_8(mem_iq_io_avail_list_8),
    .io_avail_list_9(mem_iq_io_avail_list_9),
    .io_avail_list_10(mem_iq_io_avail_list_10),
    .io_avail_list_11(mem_iq_io_avail_list_11),
    .io_avail_list_12(mem_iq_io_avail_list_12),
    .io_avail_list_13(mem_iq_io_avail_list_13),
    .io_avail_list_14(mem_iq_io_avail_list_14),
    .io_avail_list_15(mem_iq_io_avail_list_15),
    .io_avail_list_16(mem_iq_io_avail_list_16),
    .io_avail_list_17(mem_iq_io_avail_list_17),
    .io_avail_list_18(mem_iq_io_avail_list_18),
    .io_avail_list_19(mem_iq_io_avail_list_19),
    .io_avail_list_20(mem_iq_io_avail_list_20),
    .io_avail_list_21(mem_iq_io_avail_list_21),
    .io_avail_list_22(mem_iq_io_avail_list_22),
    .io_avail_list_23(mem_iq_io_avail_list_23),
    .io_avail_list_24(mem_iq_io_avail_list_24),
    .io_avail_list_25(mem_iq_io_avail_list_25),
    .io_avail_list_26(mem_iq_io_avail_list_26),
    .io_avail_list_27(mem_iq_io_avail_list_27),
    .io_avail_list_28(mem_iq_io_avail_list_28),
    .io_avail_list_29(mem_iq_io_avail_list_29),
    .io_avail_list_30(mem_iq_io_avail_list_30),
    .io_avail_list_31(mem_iq_io_avail_list_31),
    .io_avail_list_32(mem_iq_io_avail_list_32),
    .io_avail_list_33(mem_iq_io_avail_list_33),
    .io_avail_list_34(mem_iq_io_avail_list_34),
    .io_avail_list_35(mem_iq_io_avail_list_35),
    .io_avail_list_36(mem_iq_io_avail_list_36),
    .io_avail_list_37(mem_iq_io_avail_list_37),
    .io_avail_list_38(mem_iq_io_avail_list_38),
    .io_avail_list_39(mem_iq_io_avail_list_39),
    .io_avail_list_40(mem_iq_io_avail_list_40),
    .io_avail_list_41(mem_iq_io_avail_list_41),
    .io_avail_list_42(mem_iq_io_avail_list_42),
    .io_avail_list_43(mem_iq_io_avail_list_43),
    .io_avail_list_44(mem_iq_io_avail_list_44),
    .io_avail_list_45(mem_iq_io_avail_list_45),
    .io_avail_list_46(mem_iq_io_avail_list_46),
    .io_avail_list_47(mem_iq_io_avail_list_47),
    .io_avail_list_48(mem_iq_io_avail_list_48),
    .io_avail_list_49(mem_iq_io_avail_list_49),
    .io_avail_list_50(mem_iq_io_avail_list_50),
    .io_avail_list_51(mem_iq_io_avail_list_51),
    .io_avail_list_52(mem_iq_io_avail_list_52),
    .io_avail_list_53(mem_iq_io_avail_list_53),
    .io_avail_list_54(mem_iq_io_avail_list_54),
    .io_avail_list_55(mem_iq_io_avail_list_55),
    .io_avail_list_56(mem_iq_io_avail_list_56),
    .io_avail_list_57(mem_iq_io_avail_list_57),
    .io_avail_list_58(mem_iq_io_avail_list_58),
    .io_avail_list_59(mem_iq_io_avail_list_59),
    .io_avail_list_60(mem_iq_io_avail_list_60),
    .io_avail_list_61(mem_iq_io_avail_list_61),
    .io_avail_list_62(mem_iq_io_avail_list_62),
    .io_avail_list_63(mem_iq_io_avail_list_63),
    .io_fu_ready(mem_iq_io_fu_ready)
  );
  assign io_in_ready = int_iq_io_in_ready & mem_iq_io_in_ready; // @[IssueUnit.scala 68:37]
  assign io_out_0_valid = int_iq_io_out_0_valid; // @[IssueUnit.scala 64:15]
  assign io_out_0_pc = int_iq_io_out_0_pc; // @[IssueUnit.scala 64:15]
  assign io_out_0_npc = int_iq_io_out_0_npc; // @[IssueUnit.scala 64:15]
  assign io_out_0_inst = int_iq_io_out_0_inst; // @[IssueUnit.scala 64:15]
  assign io_out_0_fu_code = int_iq_io_out_0_fu_code; // @[IssueUnit.scala 64:15]
  assign io_out_0_alu_code = int_iq_io_out_0_alu_code; // @[IssueUnit.scala 64:15]
  assign io_out_0_jmp_code = int_iq_io_out_0_jmp_code; // @[IssueUnit.scala 64:15]
  assign io_out_0_sys_code = int_iq_io_out_0_sys_code; // @[IssueUnit.scala 64:15]
  assign io_out_0_w_type = int_iq_io_out_0_w_type; // @[IssueUnit.scala 64:15]
  assign io_out_0_rs1_src = int_iq_io_out_0_rs1_src; // @[IssueUnit.scala 64:15]
  assign io_out_0_rs2_src = int_iq_io_out_0_rs2_src; // @[IssueUnit.scala 64:15]
  assign io_out_0_rd_en = int_iq_io_out_0_rd_en; // @[IssueUnit.scala 64:15]
  assign io_out_0_imm = int_iq_io_out_0_imm; // @[IssueUnit.scala 64:15]
  assign io_out_0_pred_br = int_iq_io_out_0_pred_br; // @[IssueUnit.scala 64:15]
  assign io_out_0_pred_bpc = int_iq_io_out_0_pred_bpc; // @[IssueUnit.scala 64:15]
  assign io_out_0_rs1_paddr = int_iq_io_out_0_rs1_paddr; // @[IssueUnit.scala 64:15]
  assign io_out_0_rs2_paddr = int_iq_io_out_0_rs2_paddr; // @[IssueUnit.scala 64:15]
  assign io_out_0_rd_paddr = int_iq_io_out_0_rd_paddr; // @[IssueUnit.scala 64:15]
  assign io_out_0_rob_addr = int_iq_io_out_0_rob_addr; // @[IssueUnit.scala 64:15]
  assign io_out_1_valid = int_iq_io_out_1_valid; // @[IssueUnit.scala 64:15]
  assign io_out_1_pc = int_iq_io_out_1_pc; // @[IssueUnit.scala 64:15]
  assign io_out_1_npc = int_iq_io_out_1_npc; // @[IssueUnit.scala 64:15]
  assign io_out_1_fu_code = int_iq_io_out_1_fu_code; // @[IssueUnit.scala 64:15]
  assign io_out_1_alu_code = int_iq_io_out_1_alu_code; // @[IssueUnit.scala 64:15]
  assign io_out_1_jmp_code = int_iq_io_out_1_jmp_code; // @[IssueUnit.scala 64:15]
  assign io_out_1_w_type = int_iq_io_out_1_w_type; // @[IssueUnit.scala 64:15]
  assign io_out_1_rs1_src = int_iq_io_out_1_rs1_src; // @[IssueUnit.scala 64:15]
  assign io_out_1_rs2_src = int_iq_io_out_1_rs2_src; // @[IssueUnit.scala 64:15]
  assign io_out_1_rd_en = int_iq_io_out_1_rd_en; // @[IssueUnit.scala 64:15]
  assign io_out_1_imm = int_iq_io_out_1_imm; // @[IssueUnit.scala 64:15]
  assign io_out_1_pred_br = int_iq_io_out_1_pred_br; // @[IssueUnit.scala 64:15]
  assign io_out_1_pred_bpc = int_iq_io_out_1_pred_bpc; // @[IssueUnit.scala 64:15]
  assign io_out_1_rs1_paddr = int_iq_io_out_1_rs1_paddr; // @[IssueUnit.scala 64:15]
  assign io_out_1_rs2_paddr = int_iq_io_out_1_rs2_paddr; // @[IssueUnit.scala 64:15]
  assign io_out_1_rd_paddr = int_iq_io_out_1_rd_paddr; // @[IssueUnit.scala 64:15]
  assign io_out_1_rob_addr = int_iq_io_out_1_rob_addr; // @[IssueUnit.scala 64:15]
  assign io_out_2_valid = mem_iq_io_out_0_valid; // @[IssueUnit.scala 66:26]
  assign io_out_2_pc = mem_iq_io_out_0_pc; // @[IssueUnit.scala 66:26]
  assign io_out_2_fu_code = mem_iq_io_out_0_fu_code; // @[IssueUnit.scala 66:26]
  assign io_out_2_alu_code = mem_iq_io_out_0_alu_code; // @[IssueUnit.scala 66:26]
  assign io_out_2_mem_code = mem_iq_io_out_0_mem_code; // @[IssueUnit.scala 66:26]
  assign io_out_2_mem_size = mem_iq_io_out_0_mem_size; // @[IssueUnit.scala 66:26]
  assign io_out_2_w_type = mem_iq_io_out_0_w_type; // @[IssueUnit.scala 66:26]
  assign io_out_2_rs1_src = mem_iq_io_out_0_rs1_src; // @[IssueUnit.scala 66:26]
  assign io_out_2_rs2_src = mem_iq_io_out_0_rs2_src; // @[IssueUnit.scala 66:26]
  assign io_out_2_rd_en = mem_iq_io_out_0_rd_en; // @[IssueUnit.scala 66:26]
  assign io_out_2_imm = mem_iq_io_out_0_imm; // @[IssueUnit.scala 66:26]
  assign io_out_2_rs1_paddr = mem_iq_io_out_0_rs1_paddr; // @[IssueUnit.scala 66:26]
  assign io_out_2_rs2_paddr = mem_iq_io_out_0_rs2_paddr; // @[IssueUnit.scala 66:26]
  assign io_out_2_rd_paddr = mem_iq_io_out_0_rd_paddr; // @[IssueUnit.scala 66:26]
  assign io_out_2_rob_addr = mem_iq_io_out_0_rob_addr; // @[IssueUnit.scala 66:26]
  assign int_iq_clock = clock;
  assign int_iq_reset = reset;
  assign int_iq_io_flush = io_flush; // @[IssueUnit.scala 25:19]
  assign int_iq_io_in_valid = io_in_valid & |_T_260 & mem_iq_io_in_ready; // @[IssueUnit.scala 57:70]
  assign int_iq_io_in_bits_vec_0_valid = io_in_bits_vec_0_fu_code == 3'h4 ? 1'h0 : io_in_bits_vec_0_valid; // @[IssueUnit.scala 44:11 48:49 49:24]
  assign int_iq_io_in_bits_vec_0_pc = io_in_bits_vec_0_pc; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_npc = io_in_bits_vec_0_npc; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_inst = io_in_bits_vec_0_inst; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_fu_code = io_in_bits_vec_0_fu_code; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_alu_code = io_in_bits_vec_0_alu_code; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_jmp_code = io_in_bits_vec_0_jmp_code; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_sys_code = io_in_bits_vec_0_sys_code; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_w_type = io_in_bits_vec_0_w_type; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_rs1_src = io_in_bits_vec_0_rs1_src; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_rs2_src = io_in_bits_vec_0_rs2_src; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_rd_en = io_in_bits_vec_0_rd_en; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_imm = io_in_bits_vec_0_imm; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_pred_br = io_in_bits_vec_0_pred_br; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_pred_bpc = io_in_bits_vec_0_pred_bpc; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_rs1_paddr = io_in_bits_vec_0_rs1_paddr; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_rs2_paddr = io_in_bits_vec_0_rs2_paddr; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_0_rd_paddr = io_in_bits_vec_0_rd_paddr; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_valid = io_in_bits_vec_1_fu_code == 3'h4 ? 1'h0 : io_in_bits_vec_1_valid; // @[IssueUnit.scala 44:11 48:49 49:24]
  assign int_iq_io_in_bits_vec_1_pc = io_in_bits_vec_1_pc; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_npc = io_in_bits_vec_1_npc; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_inst = io_in_bits_vec_1_inst; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_fu_code = io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_alu_code = io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_jmp_code = io_in_bits_vec_1_jmp_code; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_sys_code = io_in_bits_vec_1_sys_code; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_w_type = io_in_bits_vec_1_w_type; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_rs1_src = io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_rs2_src = io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_rd_en = io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_imm = io_in_bits_vec_1_imm; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_pred_br = io_in_bits_vec_1_pred_br; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_pred_bpc = io_in_bits_vec_1_pred_bpc; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_rs1_paddr = io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_rs2_paddr = io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 56:25]
  assign int_iq_io_in_bits_vec_1_rd_paddr = io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 56:25]
  assign int_iq_io_rob_addr_0 = io_rob_addr_0; // @[IssueUnit.scala 26:22]
  assign int_iq_io_rob_addr_1 = io_rob_addr_1; // @[IssueUnit.scala 26:22]
  assign int_iq_io_avail_list_0 = io_avail_list[0]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_1 = io_avail_list[1]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_2 = io_avail_list[2]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_3 = io_avail_list[3]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_4 = io_avail_list[4]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_5 = io_avail_list[5]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_6 = io_avail_list[6]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_7 = io_avail_list[7]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_8 = io_avail_list[8]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_9 = io_avail_list[9]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_10 = io_avail_list[10]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_11 = io_avail_list[11]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_12 = io_avail_list[12]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_13 = io_avail_list[13]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_14 = io_avail_list[14]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_15 = io_avail_list[15]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_16 = io_avail_list[16]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_17 = io_avail_list[17]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_18 = io_avail_list[18]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_19 = io_avail_list[19]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_20 = io_avail_list[20]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_21 = io_avail_list[21]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_22 = io_avail_list[22]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_23 = io_avail_list[23]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_24 = io_avail_list[24]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_25 = io_avail_list[25]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_26 = io_avail_list[26]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_27 = io_avail_list[27]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_28 = io_avail_list[28]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_29 = io_avail_list[29]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_30 = io_avail_list[30]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_31 = io_avail_list[31]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_32 = io_avail_list[32]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_33 = io_avail_list[33]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_34 = io_avail_list[34]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_35 = io_avail_list[35]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_36 = io_avail_list[36]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_37 = io_avail_list[37]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_38 = io_avail_list[38]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_39 = io_avail_list[39]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_40 = io_avail_list[40]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_41 = io_avail_list[41]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_42 = io_avail_list[42]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_43 = io_avail_list[43]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_44 = io_avail_list[44]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_45 = io_avail_list[45]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_46 = io_avail_list[46]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_47 = io_avail_list[47]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_48 = io_avail_list[48]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_49 = io_avail_list[49]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_50 = io_avail_list[50]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_51 = io_avail_list[51]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_52 = io_avail_list[52]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_53 = io_avail_list[53]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_54 = io_avail_list[54]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_55 = io_avail_list[55]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_56 = io_avail_list[56]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_57 = io_avail_list[57]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_58 = io_avail_list[58]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_59 = io_avail_list[59]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_60 = io_avail_list[60]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_61 = io_avail_list[61]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_62 = io_avail_list[62]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_avail_list_63 = io_avail_list[63]; // @[IssueUnit.scala 28:45]
  assign int_iq_io_sys_ready = io_sys_ready; // @[IssueUnit.scala 58:23]
  assign mem_iq_clock = clock;
  assign mem_iq_reset = reset;
  assign mem_iq_io_flush = io_flush; // @[IssueUnit.scala 33:19]
  assign mem_iq_io_in_valid = io_in_valid & |_T_264 & int_iq_io_in_ready; // @[IssueUnit.scala 60:70]
  assign mem_iq_io_in_bits_vec_0_valid = io_in_bits_vec_0_fu_code != 3'h4 ? 1'h0 : io_in_bits_vec_0_valid; // @[IssueUnit.scala 45:11 51:49 52:24]
  assign mem_iq_io_in_bits_vec_0_pc = io_in_bits_vec_0_pc; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_0_fu_code = io_in_bits_vec_0_fu_code; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_0_alu_code = io_in_bits_vec_0_alu_code; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_0_mem_code = io_in_bits_vec_0_mem_code; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_0_mem_size = io_in_bits_vec_0_mem_size; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_0_w_type = io_in_bits_vec_0_w_type; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_0_rs1_src = io_in_bits_vec_0_rs1_src; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_0_rs2_src = io_in_bits_vec_0_rs2_src; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_0_rd_en = io_in_bits_vec_0_rd_en; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_0_imm = io_in_bits_vec_0_imm; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_0_rs1_paddr = io_in_bits_vec_0_rs1_paddr; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_0_rs2_paddr = io_in_bits_vec_0_rs2_paddr; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_0_rd_paddr = io_in_bits_vec_0_rd_paddr; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_1_valid = io_in_bits_vec_1_fu_code != 3'h4 ? 1'h0 : io_in_bits_vec_1_valid; // @[IssueUnit.scala 45:11 51:49 52:24]
  assign mem_iq_io_in_bits_vec_1_pc = io_in_bits_vec_1_pc; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_1_fu_code = io_in_bits_vec_1_fu_code; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_1_alu_code = io_in_bits_vec_1_alu_code; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_1_mem_code = io_in_bits_vec_1_mem_code; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_1_mem_size = io_in_bits_vec_1_mem_size; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_1_w_type = io_in_bits_vec_1_w_type; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_1_rs1_src = io_in_bits_vec_1_rs1_src; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_1_rs2_src = io_in_bits_vec_1_rs2_src; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_1_rd_en = io_in_bits_vec_1_rd_en; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_1_imm = io_in_bits_vec_1_imm; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_1_rs1_paddr = io_in_bits_vec_1_rs1_paddr; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_1_rs2_paddr = io_in_bits_vec_1_rs2_paddr; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_in_bits_vec_1_rd_paddr = io_in_bits_vec_1_rd_paddr; // @[IssueUnit.scala 59:25]
  assign mem_iq_io_rob_addr_0 = io_rob_addr_0; // @[IssueUnit.scala 34:22]
  assign mem_iq_io_rob_addr_1 = io_rob_addr_1; // @[IssueUnit.scala 34:22]
  assign mem_iq_io_avail_list_0 = io_avail_list[0]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_1 = io_avail_list[1]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_2 = io_avail_list[2]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_3 = io_avail_list[3]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_4 = io_avail_list[4]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_5 = io_avail_list[5]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_6 = io_avail_list[6]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_7 = io_avail_list[7]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_8 = io_avail_list[8]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_9 = io_avail_list[9]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_10 = io_avail_list[10]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_11 = io_avail_list[11]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_12 = io_avail_list[12]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_13 = io_avail_list[13]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_14 = io_avail_list[14]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_15 = io_avail_list[15]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_16 = io_avail_list[16]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_17 = io_avail_list[17]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_18 = io_avail_list[18]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_19 = io_avail_list[19]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_20 = io_avail_list[20]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_21 = io_avail_list[21]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_22 = io_avail_list[22]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_23 = io_avail_list[23]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_24 = io_avail_list[24]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_25 = io_avail_list[25]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_26 = io_avail_list[26]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_27 = io_avail_list[27]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_28 = io_avail_list[28]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_29 = io_avail_list[29]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_30 = io_avail_list[30]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_31 = io_avail_list[31]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_32 = io_avail_list[32]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_33 = io_avail_list[33]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_34 = io_avail_list[34]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_35 = io_avail_list[35]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_36 = io_avail_list[36]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_37 = io_avail_list[37]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_38 = io_avail_list[38]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_39 = io_avail_list[39]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_40 = io_avail_list[40]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_41 = io_avail_list[41]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_42 = io_avail_list[42]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_43 = io_avail_list[43]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_44 = io_avail_list[44]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_45 = io_avail_list[45]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_46 = io_avail_list[46]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_47 = io_avail_list[47]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_48 = io_avail_list[48]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_49 = io_avail_list[49]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_50 = io_avail_list[50]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_51 = io_avail_list[51]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_52 = io_avail_list[52]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_53 = io_avail_list[53]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_54 = io_avail_list[54]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_55 = io_avail_list[55]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_56 = io_avail_list[56]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_57 = io_avail_list[57]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_58 = io_avail_list[58]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_59 = io_avail_list[59]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_60 = io_avail_list[60]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_61 = io_avail_list[61]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_62 = io_avail_list[62]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_avail_list_63 = io_avail_list[63]; // @[IssueUnit.scala 36:45]
  assign mem_iq_io_fu_ready = io_lsu_ready; // @[IssueUnit.scala 38:22]
endmodule
module ysyx_210128_Prf(
  input         clock,
  input         reset,
  input         io_in_0_valid,
  input  [31:0] io_in_0_pc,
  input  [31:0] io_in_0_npc,
  input  [31:0] io_in_0_inst,
  input  [2:0]  io_in_0_fu_code,
  input  [3:0]  io_in_0_alu_code,
  input  [3:0]  io_in_0_jmp_code,
  input  [2:0]  io_in_0_sys_code,
  input         io_in_0_w_type,
  input  [1:0]  io_in_0_rs1_src,
  input  [1:0]  io_in_0_rs2_src,
  input         io_in_0_rd_en,
  input  [31:0] io_in_0_imm,
  input         io_in_0_pred_br,
  input  [31:0] io_in_0_pred_bpc,
  input  [5:0]  io_in_0_rs1_paddr,
  input  [5:0]  io_in_0_rs2_paddr,
  input  [5:0]  io_in_0_rd_paddr,
  input  [3:0]  io_in_0_rob_addr,
  input         io_in_1_valid,
  input  [31:0] io_in_1_pc,
  input  [31:0] io_in_1_npc,
  input  [2:0]  io_in_1_fu_code,
  input  [3:0]  io_in_1_alu_code,
  input  [3:0]  io_in_1_jmp_code,
  input         io_in_1_w_type,
  input  [1:0]  io_in_1_rs1_src,
  input  [1:0]  io_in_1_rs2_src,
  input         io_in_1_rd_en,
  input  [31:0] io_in_1_imm,
  input         io_in_1_pred_br,
  input  [31:0] io_in_1_pred_bpc,
  input  [5:0]  io_in_1_rs1_paddr,
  input  [5:0]  io_in_1_rs2_paddr,
  input  [5:0]  io_in_1_rd_paddr,
  input  [3:0]  io_in_1_rob_addr,
  input         io_in_2_valid,
  input  [31:0] io_in_2_pc,
  input  [2:0]  io_in_2_fu_code,
  input  [3:0]  io_in_2_alu_code,
  input  [1:0]  io_in_2_mem_code,
  input  [1:0]  io_in_2_mem_size,
  input         io_in_2_w_type,
  input  [1:0]  io_in_2_rs1_src,
  input  [1:0]  io_in_2_rs2_src,
  input         io_in_2_rd_en,
  input  [31:0] io_in_2_imm,
  input  [5:0]  io_in_2_rs1_paddr,
  input  [5:0]  io_in_2_rs2_paddr,
  input  [5:0]  io_in_2_rd_paddr,
  input  [3:0]  io_in_2_rob_addr,
  output        io_out_0_valid,
  output [31:0] io_out_0_pc,
  output [31:0] io_out_0_npc,
  output [31:0] io_out_0_inst,
  output [2:0]  io_out_0_fu_code,
  output [3:0]  io_out_0_alu_code,
  output [3:0]  io_out_0_jmp_code,
  output [2:0]  io_out_0_sys_code,
  output        io_out_0_w_type,
  output [1:0]  io_out_0_rs1_src,
  output [1:0]  io_out_0_rs2_src,
  output        io_out_0_rd_en,
  output [31:0] io_out_0_imm,
  output        io_out_0_pred_br,
  output [31:0] io_out_0_pred_bpc,
  output [5:0]  io_out_0_rd_paddr,
  output [3:0]  io_out_0_rob_addr,
  output        io_out_1_valid,
  output [31:0] io_out_1_pc,
  output [31:0] io_out_1_npc,
  output [2:0]  io_out_1_fu_code,
  output [3:0]  io_out_1_alu_code,
  output [3:0]  io_out_1_jmp_code,
  output        io_out_1_w_type,
  output [1:0]  io_out_1_rs1_src,
  output [1:0]  io_out_1_rs2_src,
  output        io_out_1_rd_en,
  output [31:0] io_out_1_imm,
  output        io_out_1_pred_br,
  output [31:0] io_out_1_pred_bpc,
  output [5:0]  io_out_1_rd_paddr,
  output [3:0]  io_out_1_rob_addr,
  output        io_out_2_valid,
  output [31:0] io_out_2_pc,
  output [2:0]  io_out_2_fu_code,
  output [3:0]  io_out_2_alu_code,
  output [1:0]  io_out_2_mem_code,
  output [1:0]  io_out_2_mem_size,
  output        io_out_2_w_type,
  output [1:0]  io_out_2_rs1_src,
  output [1:0]  io_out_2_rs2_src,
  output        io_out_2_rd_en,
  output [31:0] io_out_2_imm,
  output [5:0]  io_out_2_rd_paddr,
  output [3:0]  io_out_2_rob_addr,
  output [63:0] io_rs1_data_0,
  output [63:0] io_rs1_data_1,
  output [63:0] io_rs1_data_2,
  output [63:0] io_rs2_data_0,
  output [63:0] io_rs2_data_1,
  output [63:0] io_rs2_data_2,
  input         io_rd_en_0,
  input         io_rd_en_1,
  input         io_rd_en_2,
  input  [5:0]  io_rd_paddr_0,
  input  [5:0]  io_rd_paddr_1,
  input  [5:0]  io_rd_paddr_2,
  input  [63:0] io_rd_data_0,
  input  [63:0] io_rd_data_1,
  input  [63:0] io_rd_data_2,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] prf [0:63]; // @[Prf.scala 20:16]
//   wire  prf_MPORT_3_en; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_3_addr; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_3_data; // @[Prf.scala 20:16]
//   wire  prf_MPORT_4_en; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_4_addr; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_4_data; // @[Prf.scala 20:16]
//   wire  prf_MPORT_5_en; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_5_addr; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_5_data; // @[Prf.scala 20:16]
//   wire  prf_MPORT_6_en; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_6_addr; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_6_data; // @[Prf.scala 20:16]
//   wire  prf_MPORT_7_en; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_7_addr; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_7_data; // @[Prf.scala 20:16]
//   wire  prf_MPORT_8_en; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_8_addr; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_8_data; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_1_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_1_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_1_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_1_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_2_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_2_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_2_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_2_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_9_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_9_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_9_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_9_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_10_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_10_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_10_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_10_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_11_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_11_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_11_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_11_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_12_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_12_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_12_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_12_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_13_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_13_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_13_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_13_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_14_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_14_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_14_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_14_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_15_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_15_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_15_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_15_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_16_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_16_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_16_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_16_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_17_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_17_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_17_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_17_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_18_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_18_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_18_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_18_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_19_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_19_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_19_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_19_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_20_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_20_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_20_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_20_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_21_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_21_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_21_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_21_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_22_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_22_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_22_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_22_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_23_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_23_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_23_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_23_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_24_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_24_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_24_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_24_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_25_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_25_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_25_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_25_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_26_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_26_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_26_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_26_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_27_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_27_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_27_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_27_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_28_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_28_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_28_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_28_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_29_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_29_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_29_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_29_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_30_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_30_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_30_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_30_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_31_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_31_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_31_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_31_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_32_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_32_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_32_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_32_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_33_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_33_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_33_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_33_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_34_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_34_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_34_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_34_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_35_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_35_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_35_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_35_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_36_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_36_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_36_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_36_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_37_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_37_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_37_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_37_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_38_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_38_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_38_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_38_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_39_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_39_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_39_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_39_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_40_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_40_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_40_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_40_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_41_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_41_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_41_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_41_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_42_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_42_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_42_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_42_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_43_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_43_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_43_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_43_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_44_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_44_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_44_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_44_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_45_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_45_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_45_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_45_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_46_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_46_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_46_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_46_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_47_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_47_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_47_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_47_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_48_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_48_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_48_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_48_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_49_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_49_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_49_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_49_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_50_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_50_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_50_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_50_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_51_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_51_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_51_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_51_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_52_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_52_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_52_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_52_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_53_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_53_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_53_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_53_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_54_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_54_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_54_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_54_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_55_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_55_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_55_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_55_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_56_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_56_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_56_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_56_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_57_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_57_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_57_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_57_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_58_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_58_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_58_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_58_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_59_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_59_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_59_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_59_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_60_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_60_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_60_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_60_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_61_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_61_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_61_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_61_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_62_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_62_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_62_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_62_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_63_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_63_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_63_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_63_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_64_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_64_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_64_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_64_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_65_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_65_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_65_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_65_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_66_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_66_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_66_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_66_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_67_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_67_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_67_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_67_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_68_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_68_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_68_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_68_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_69_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_69_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_69_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_69_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_70_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_70_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_70_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_70_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_71_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_71_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_71_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_71_en; // @[Prf.scala 20:16]
  wire [63:0] prf_MPORT_72_data; // @[Prf.scala 20:16]
  wire [5:0] prf_MPORT_72_addr; // @[Prf.scala 20:16]
  wire  prf_MPORT_72_mask; // @[Prf.scala 20:16]
  wire  prf_MPORT_72_en; // @[Prf.scala 20:16]
  wire  _T = io_rd_paddr_0 != 6'h0; // @[Prf.scala 23:42]
  wire  _T_1 = io_rd_en_0 & io_rd_paddr_0 != 6'h0; // @[Prf.scala 23:23]
  wire  _T_2 = io_rd_paddr_1 != 6'h0; // @[Prf.scala 23:42]
  wire  _T_3 = io_rd_en_1 & io_rd_paddr_1 != 6'h0; // @[Prf.scala 23:23]
  wire  _T_4 = io_rd_paddr_2 != 6'h0; // @[Prf.scala 23:42]
  wire [63:0] _T_7 = io_in_0_rs1_paddr != 6'h0 ? prf_MPORT_3_data : 64'h0; // @[Prf.scala 34:23]
  wire [63:0] _T_9 = io_in_0_rs2_paddr != 6'h0 ? prf_MPORT_4_data : 64'h0; // @[Prf.scala 35:23]
  wire [63:0] _T_11 = io_in_1_rs1_paddr != 6'h0 ? prf_MPORT_5_data : 64'h0; // @[Prf.scala 34:23]
  wire [63:0] _T_13 = io_in_1_rs2_paddr != 6'h0 ? prf_MPORT_6_data : 64'h0; // @[Prf.scala 35:23]
  wire [63:0] _T_15 = io_in_2_rs1_paddr != 6'h0 ? prf_MPORT_7_data : 64'h0; // @[Prf.scala 34:23]
  wire [63:0] _T_17 = io_in_2_rs2_paddr != 6'h0 ? prf_MPORT_8_data : 64'h0; // @[Prf.scala 35:23]
  wire [63:0] _GEN_15 = io_rd_paddr_0 == io_in_0_rs1_paddr ? io_rd_data_0 : _T_7; // @[Prf.scala 34:17 42:48 43:23]
  wire [63:0] _GEN_16 = io_rd_paddr_0 == io_in_0_rs2_paddr ? io_rd_data_0 : _T_9; // @[Prf.scala 35:17 45:48 46:23]
  wire [63:0] _GEN_17 = _T_1 ? _GEN_15 : _T_7; // @[Prf.scala 34:17 41:54]
  wire [63:0] _GEN_18 = _T_1 ? _GEN_16 : _T_9; // @[Prf.scala 35:17 41:54]
  wire [63:0] _GEN_23 = io_rd_paddr_0 == io_in_1_rs1_paddr ? io_rd_data_0 : _T_11; // @[Prf.scala 34:17 42:48 43:23]
  wire [63:0] _GEN_24 = io_rd_paddr_0 == io_in_1_rs2_paddr ? io_rd_data_0 : _T_13; // @[Prf.scala 35:17 45:48 46:23]
  wire [63:0] _GEN_25 = _T_1 ? _GEN_23 : _T_11; // @[Prf.scala 34:17 41:54]
  wire [63:0] _GEN_26 = _T_1 ? _GEN_24 : _T_13; // @[Prf.scala 35:17 41:54]
  wire [63:0] _GEN_31 = io_rd_paddr_0 == io_in_2_rs1_paddr ? io_rd_data_0 : _T_15; // @[Prf.scala 34:17 42:48 43:23]
  wire [63:0] _GEN_32 = io_rd_paddr_0 == io_in_2_rs2_paddr ? io_rd_data_0 : _T_17; // @[Prf.scala 35:17 45:48 46:23]
  wire [63:0] _GEN_33 = _T_1 ? _GEN_31 : _T_15; // @[Prf.scala 34:17 41:54]
  wire [63:0] _GEN_34 = _T_1 ? _GEN_32 : _T_17; // @[Prf.scala 35:17 41:54]
  reg  out_uop_0_valid; // @[Prf.scala 60:24]
  reg [31:0] out_uop_0_pc; // @[Prf.scala 60:24]
  reg [31:0] out_uop_0_npc; // @[Prf.scala 60:24]
  reg [31:0] out_uop_0_inst; // @[Prf.scala 60:24]
  reg [2:0] out_uop_0_fu_code; // @[Prf.scala 60:24]
  reg [3:0] out_uop_0_alu_code; // @[Prf.scala 60:24]
  reg [3:0] out_uop_0_jmp_code; // @[Prf.scala 60:24]
  reg [2:0] out_uop_0_sys_code; // @[Prf.scala 60:24]
  reg  out_uop_0_w_type; // @[Prf.scala 60:24]
  reg [1:0] out_uop_0_rs1_src; // @[Prf.scala 60:24]
  reg [1:0] out_uop_0_rs2_src; // @[Prf.scala 60:24]
  reg  out_uop_0_rd_en; // @[Prf.scala 60:24]
  reg [31:0] out_uop_0_imm; // @[Prf.scala 60:24]
  reg  out_uop_0_pred_br; // @[Prf.scala 60:24]
  reg [31:0] out_uop_0_pred_bpc; // @[Prf.scala 60:24]
  reg [5:0] out_uop_0_rd_paddr; // @[Prf.scala 60:24]
  reg [3:0] out_uop_0_rob_addr; // @[Prf.scala 60:24]
  reg  out_uop_1_valid; // @[Prf.scala 60:24]
  reg [31:0] out_uop_1_pc; // @[Prf.scala 60:24]
  reg [31:0] out_uop_1_npc; // @[Prf.scala 60:24]
  reg [2:0] out_uop_1_fu_code; // @[Prf.scala 60:24]
  reg [3:0] out_uop_1_alu_code; // @[Prf.scala 60:24]
  reg [3:0] out_uop_1_jmp_code; // @[Prf.scala 60:24]
  reg  out_uop_1_w_type; // @[Prf.scala 60:24]
  reg [1:0] out_uop_1_rs1_src; // @[Prf.scala 60:24]
  reg [1:0] out_uop_1_rs2_src; // @[Prf.scala 60:24]
  reg  out_uop_1_rd_en; // @[Prf.scala 60:24]
  reg [31:0] out_uop_1_imm; // @[Prf.scala 60:24]
  reg  out_uop_1_pred_br; // @[Prf.scala 60:24]
  reg [31:0] out_uop_1_pred_bpc; // @[Prf.scala 60:24]
  reg [5:0] out_uop_1_rd_paddr; // @[Prf.scala 60:24]
  reg [3:0] out_uop_1_rob_addr; // @[Prf.scala 60:24]
  reg  out_uop_2_valid; // @[Prf.scala 60:24]
  reg [31:0] out_uop_2_pc; // @[Prf.scala 60:24]
  reg [2:0] out_uop_2_fu_code; // @[Prf.scala 60:24]
  reg [3:0] out_uop_2_alu_code; // @[Prf.scala 60:24]
  reg [1:0] out_uop_2_mem_code; // @[Prf.scala 60:24]
  reg [1:0] out_uop_2_mem_size; // @[Prf.scala 60:24]
  reg  out_uop_2_w_type; // @[Prf.scala 60:24]
  reg [1:0] out_uop_2_rs1_src; // @[Prf.scala 60:24]
  reg [1:0] out_uop_2_rs2_src; // @[Prf.scala 60:24]
  reg  out_uop_2_rd_en; // @[Prf.scala 60:24]
  reg [31:0] out_uop_2_imm; // @[Prf.scala 60:24]
  reg [5:0] out_uop_2_rd_paddr; // @[Prf.scala 60:24]
  reg [3:0] out_uop_2_rob_addr; // @[Prf.scala 60:24]
  reg [63:0] out_rs1_data_0; // @[Prf.scala 61:29]
  reg [63:0] out_rs1_data_1; // @[Prf.scala 61:29]
  reg [63:0] out_rs1_data_2; // @[Prf.scala 61:29]
  reg [63:0] out_rs2_data_0; // @[Prf.scala 62:29]
  reg [63:0] out_rs2_data_1; // @[Prf.scala 62:29]
  reg [63:0] out_rs2_data_2; // @[Prf.scala 62:29]
//   assign prf_MPORT_3_en = 1'h1;
  assign prf_MPORT_3_addr = io_in_0_rs1_paddr;
  assign prf_MPORT_3_data = prf[prf_MPORT_3_addr]; // @[Prf.scala 20:16]
//   assign prf_MPORT_4_en = 1'h1;
  assign prf_MPORT_4_addr = io_in_0_rs2_paddr;
  assign prf_MPORT_4_data = prf[prf_MPORT_4_addr]; // @[Prf.scala 20:16]
//   assign prf_MPORT_5_en = 1'h1;
  assign prf_MPORT_5_addr = io_in_1_rs1_paddr;
  assign prf_MPORT_5_data = prf[prf_MPORT_5_addr]; // @[Prf.scala 20:16]
//   assign prf_MPORT_6_en = 1'h1;
  assign prf_MPORT_6_addr = io_in_1_rs2_paddr;
  assign prf_MPORT_6_data = prf[prf_MPORT_6_addr]; // @[Prf.scala 20:16]
//   assign prf_MPORT_7_en = 1'h1;
  assign prf_MPORT_7_addr = io_in_2_rs1_paddr;
  assign prf_MPORT_7_data = prf[prf_MPORT_7_addr]; // @[Prf.scala 20:16]
//   assign prf_MPORT_8_en = 1'h1;
  assign prf_MPORT_8_addr = io_in_2_rs2_paddr;
  assign prf_MPORT_8_data = prf[prf_MPORT_8_addr]; // @[Prf.scala 20:16]
  assign prf_MPORT_data = io_rd_data_0;
  assign prf_MPORT_addr = io_rd_paddr_0;
  assign prf_MPORT_mask = 1'h1;
  assign prf_MPORT_en = io_rd_en_0 & _T;
  assign prf_MPORT_1_data = io_rd_data_1;
  assign prf_MPORT_1_addr = io_rd_paddr_1;
  assign prf_MPORT_1_mask = 1'h1;
  assign prf_MPORT_1_en = io_rd_en_1 & _T_2;
  assign prf_MPORT_2_data = io_rd_data_2;
  assign prf_MPORT_2_addr = io_rd_paddr_2;
  assign prf_MPORT_2_mask = 1'h1;
  assign prf_MPORT_2_en = io_rd_en_2 & _T_4;
  assign prf_MPORT_9_data = 64'h0;
  assign prf_MPORT_9_addr = 6'h0;
  assign prf_MPORT_9_mask = 1'h1;
  assign prf_MPORT_9_en = reset;
  assign prf_MPORT_10_data = 64'h0;
  assign prf_MPORT_10_addr = 6'h1;
  assign prf_MPORT_10_mask = 1'h1;
  assign prf_MPORT_10_en = reset;
  assign prf_MPORT_11_data = 64'h0;
  assign prf_MPORT_11_addr = 6'h2;
  assign prf_MPORT_11_mask = 1'h1;
  assign prf_MPORT_11_en = reset;
  assign prf_MPORT_12_data = 64'h0;
  assign prf_MPORT_12_addr = 6'h3;
  assign prf_MPORT_12_mask = 1'h1;
  assign prf_MPORT_12_en = reset;
  assign prf_MPORT_13_data = 64'h0;
  assign prf_MPORT_13_addr = 6'h4;
  assign prf_MPORT_13_mask = 1'h1;
  assign prf_MPORT_13_en = reset;
  assign prf_MPORT_14_data = 64'h0;
  assign prf_MPORT_14_addr = 6'h5;
  assign prf_MPORT_14_mask = 1'h1;
  assign prf_MPORT_14_en = reset;
  assign prf_MPORT_15_data = 64'h0;
  assign prf_MPORT_15_addr = 6'h6;
  assign prf_MPORT_15_mask = 1'h1;
  assign prf_MPORT_15_en = reset;
  assign prf_MPORT_16_data = 64'h0;
  assign prf_MPORT_16_addr = 6'h7;
  assign prf_MPORT_16_mask = 1'h1;
  assign prf_MPORT_16_en = reset;
  assign prf_MPORT_17_data = 64'h0;
  assign prf_MPORT_17_addr = 6'h8;
  assign prf_MPORT_17_mask = 1'h1;
  assign prf_MPORT_17_en = reset;
  assign prf_MPORT_18_data = 64'h0;
  assign prf_MPORT_18_addr = 6'h9;
  assign prf_MPORT_18_mask = 1'h1;
  assign prf_MPORT_18_en = reset;
  assign prf_MPORT_19_data = 64'h0;
  assign prf_MPORT_19_addr = 6'ha;
  assign prf_MPORT_19_mask = 1'h1;
  assign prf_MPORT_19_en = reset;
  assign prf_MPORT_20_data = 64'h0;
  assign prf_MPORT_20_addr = 6'hb;
  assign prf_MPORT_20_mask = 1'h1;
  assign prf_MPORT_20_en = reset;
  assign prf_MPORT_21_data = 64'h0;
  assign prf_MPORT_21_addr = 6'hc;
  assign prf_MPORT_21_mask = 1'h1;
  assign prf_MPORT_21_en = reset;
  assign prf_MPORT_22_data = 64'h0;
  assign prf_MPORT_22_addr = 6'hd;
  assign prf_MPORT_22_mask = 1'h1;
  assign prf_MPORT_22_en = reset;
  assign prf_MPORT_23_data = 64'h0;
  assign prf_MPORT_23_addr = 6'he;
  assign prf_MPORT_23_mask = 1'h1;
  assign prf_MPORT_23_en = reset;
  assign prf_MPORT_24_data = 64'h0;
  assign prf_MPORT_24_addr = 6'hf;
  assign prf_MPORT_24_mask = 1'h1;
  assign prf_MPORT_24_en = reset;
  assign prf_MPORT_25_data = 64'h0;
  assign prf_MPORT_25_addr = 6'h10;
  assign prf_MPORT_25_mask = 1'h1;
  assign prf_MPORT_25_en = reset;
  assign prf_MPORT_26_data = 64'h0;
  assign prf_MPORT_26_addr = 6'h11;
  assign prf_MPORT_26_mask = 1'h1;
  assign prf_MPORT_26_en = reset;
  assign prf_MPORT_27_data = 64'h0;
  assign prf_MPORT_27_addr = 6'h12;
  assign prf_MPORT_27_mask = 1'h1;
  assign prf_MPORT_27_en = reset;
  assign prf_MPORT_28_data = 64'h0;
  assign prf_MPORT_28_addr = 6'h13;
  assign prf_MPORT_28_mask = 1'h1;
  assign prf_MPORT_28_en = reset;
  assign prf_MPORT_29_data = 64'h0;
  assign prf_MPORT_29_addr = 6'h14;
  assign prf_MPORT_29_mask = 1'h1;
  assign prf_MPORT_29_en = reset;
  assign prf_MPORT_30_data = 64'h0;
  assign prf_MPORT_30_addr = 6'h15;
  assign prf_MPORT_30_mask = 1'h1;
  assign prf_MPORT_30_en = reset;
  assign prf_MPORT_31_data = 64'h0;
  assign prf_MPORT_31_addr = 6'h16;
  assign prf_MPORT_31_mask = 1'h1;
  assign prf_MPORT_31_en = reset;
  assign prf_MPORT_32_data = 64'h0;
  assign prf_MPORT_32_addr = 6'h17;
  assign prf_MPORT_32_mask = 1'h1;
  assign prf_MPORT_32_en = reset;
  assign prf_MPORT_33_data = 64'h0;
  assign prf_MPORT_33_addr = 6'h18;
  assign prf_MPORT_33_mask = 1'h1;
  assign prf_MPORT_33_en = reset;
  assign prf_MPORT_34_data = 64'h0;
  assign prf_MPORT_34_addr = 6'h19;
  assign prf_MPORT_34_mask = 1'h1;
  assign prf_MPORT_34_en = reset;
  assign prf_MPORT_35_data = 64'h0;
  assign prf_MPORT_35_addr = 6'h1a;
  assign prf_MPORT_35_mask = 1'h1;
  assign prf_MPORT_35_en = reset;
  assign prf_MPORT_36_data = 64'h0;
  assign prf_MPORT_36_addr = 6'h1b;
  assign prf_MPORT_36_mask = 1'h1;
  assign prf_MPORT_36_en = reset;
  assign prf_MPORT_37_data = 64'h0;
  assign prf_MPORT_37_addr = 6'h1c;
  assign prf_MPORT_37_mask = 1'h1;
  assign prf_MPORT_37_en = reset;
  assign prf_MPORT_38_data = 64'h0;
  assign prf_MPORT_38_addr = 6'h1d;
  assign prf_MPORT_38_mask = 1'h1;
  assign prf_MPORT_38_en = reset;
  assign prf_MPORT_39_data = 64'h0;
  assign prf_MPORT_39_addr = 6'h1e;
  assign prf_MPORT_39_mask = 1'h1;
  assign prf_MPORT_39_en = reset;
  assign prf_MPORT_40_data = 64'h0;
  assign prf_MPORT_40_addr = 6'h1f;
  assign prf_MPORT_40_mask = 1'h1;
  assign prf_MPORT_40_en = reset;
  assign prf_MPORT_41_data = 64'h0;
  assign prf_MPORT_41_addr = 6'h20;
  assign prf_MPORT_41_mask = 1'h1;
  assign prf_MPORT_41_en = reset;
  assign prf_MPORT_42_data = 64'h0;
  assign prf_MPORT_42_addr = 6'h21;
  assign prf_MPORT_42_mask = 1'h1;
  assign prf_MPORT_42_en = reset;
  assign prf_MPORT_43_data = 64'h0;
  assign prf_MPORT_43_addr = 6'h22;
  assign prf_MPORT_43_mask = 1'h1;
  assign prf_MPORT_43_en = reset;
  assign prf_MPORT_44_data = 64'h0;
  assign prf_MPORT_44_addr = 6'h23;
  assign prf_MPORT_44_mask = 1'h1;
  assign prf_MPORT_44_en = reset;
  assign prf_MPORT_45_data = 64'h0;
  assign prf_MPORT_45_addr = 6'h24;
  assign prf_MPORT_45_mask = 1'h1;
  assign prf_MPORT_45_en = reset;
  assign prf_MPORT_46_data = 64'h0;
  assign prf_MPORT_46_addr = 6'h25;
  assign prf_MPORT_46_mask = 1'h1;
  assign prf_MPORT_46_en = reset;
  assign prf_MPORT_47_data = 64'h0;
  assign prf_MPORT_47_addr = 6'h26;
  assign prf_MPORT_47_mask = 1'h1;
  assign prf_MPORT_47_en = reset;
  assign prf_MPORT_48_data = 64'h0;
  assign prf_MPORT_48_addr = 6'h27;
  assign prf_MPORT_48_mask = 1'h1;
  assign prf_MPORT_48_en = reset;
  assign prf_MPORT_49_data = 64'h0;
  assign prf_MPORT_49_addr = 6'h28;
  assign prf_MPORT_49_mask = 1'h1;
  assign prf_MPORT_49_en = reset;
  assign prf_MPORT_50_data = 64'h0;
  assign prf_MPORT_50_addr = 6'h29;
  assign prf_MPORT_50_mask = 1'h1;
  assign prf_MPORT_50_en = reset;
  assign prf_MPORT_51_data = 64'h0;
  assign prf_MPORT_51_addr = 6'h2a;
  assign prf_MPORT_51_mask = 1'h1;
  assign prf_MPORT_51_en = reset;
  assign prf_MPORT_52_data = 64'h0;
  assign prf_MPORT_52_addr = 6'h2b;
  assign prf_MPORT_52_mask = 1'h1;
  assign prf_MPORT_52_en = reset;
  assign prf_MPORT_53_data = 64'h0;
  assign prf_MPORT_53_addr = 6'h2c;
  assign prf_MPORT_53_mask = 1'h1;
  assign prf_MPORT_53_en = reset;
  assign prf_MPORT_54_data = 64'h0;
  assign prf_MPORT_54_addr = 6'h2d;
  assign prf_MPORT_54_mask = 1'h1;
  assign prf_MPORT_54_en = reset;
  assign prf_MPORT_55_data = 64'h0;
  assign prf_MPORT_55_addr = 6'h2e;
  assign prf_MPORT_55_mask = 1'h1;
  assign prf_MPORT_55_en = reset;
  assign prf_MPORT_56_data = 64'h0;
  assign prf_MPORT_56_addr = 6'h2f;
  assign prf_MPORT_56_mask = 1'h1;
  assign prf_MPORT_56_en = reset;
  assign prf_MPORT_57_data = 64'h0;
  assign prf_MPORT_57_addr = 6'h30;
  assign prf_MPORT_57_mask = 1'h1;
  assign prf_MPORT_57_en = reset;
  assign prf_MPORT_58_data = 64'h0;
  assign prf_MPORT_58_addr = 6'h31;
  assign prf_MPORT_58_mask = 1'h1;
  assign prf_MPORT_58_en = reset;
  assign prf_MPORT_59_data = 64'h0;
  assign prf_MPORT_59_addr = 6'h32;
  assign prf_MPORT_59_mask = 1'h1;
  assign prf_MPORT_59_en = reset;
  assign prf_MPORT_60_data = 64'h0;
  assign prf_MPORT_60_addr = 6'h33;
  assign prf_MPORT_60_mask = 1'h1;
  assign prf_MPORT_60_en = reset;
  assign prf_MPORT_61_data = 64'h0;
  assign prf_MPORT_61_addr = 6'h34;
  assign prf_MPORT_61_mask = 1'h1;
  assign prf_MPORT_61_en = reset;
  assign prf_MPORT_62_data = 64'h0;
  assign prf_MPORT_62_addr = 6'h35;
  assign prf_MPORT_62_mask = 1'h1;
  assign prf_MPORT_62_en = reset;
  assign prf_MPORT_63_data = 64'h0;
  assign prf_MPORT_63_addr = 6'h36;
  assign prf_MPORT_63_mask = 1'h1;
  assign prf_MPORT_63_en = reset;
  assign prf_MPORT_64_data = 64'h0;
  assign prf_MPORT_64_addr = 6'h37;
  assign prf_MPORT_64_mask = 1'h1;
  assign prf_MPORT_64_en = reset;
  assign prf_MPORT_65_data = 64'h0;
  assign prf_MPORT_65_addr = 6'h38;
  assign prf_MPORT_65_mask = 1'h1;
  assign prf_MPORT_65_en = reset;
  assign prf_MPORT_66_data = 64'h0;
  assign prf_MPORT_66_addr = 6'h39;
  assign prf_MPORT_66_mask = 1'h1;
  assign prf_MPORT_66_en = reset;
  assign prf_MPORT_67_data = 64'h0;
  assign prf_MPORT_67_addr = 6'h3a;
  assign prf_MPORT_67_mask = 1'h1;
  assign prf_MPORT_67_en = reset;
  assign prf_MPORT_68_data = 64'h0;
  assign prf_MPORT_68_addr = 6'h3b;
  assign prf_MPORT_68_mask = 1'h1;
  assign prf_MPORT_68_en = reset;
  assign prf_MPORT_69_data = 64'h0;
  assign prf_MPORT_69_addr = 6'h3c;
  assign prf_MPORT_69_mask = 1'h1;
  assign prf_MPORT_69_en = reset;
  assign prf_MPORT_70_data = 64'h0;
  assign prf_MPORT_70_addr = 6'h3d;
  assign prf_MPORT_70_mask = 1'h1;
  assign prf_MPORT_70_en = reset;
  assign prf_MPORT_71_data = 64'h0;
  assign prf_MPORT_71_addr = 6'h3e;
  assign prf_MPORT_71_mask = 1'h1;
  assign prf_MPORT_71_en = reset;
  assign prf_MPORT_72_data = 64'h0;
  assign prf_MPORT_72_addr = 6'h3f;
  assign prf_MPORT_72_mask = 1'h1;
  assign prf_MPORT_72_en = reset;
  assign io_out_0_valid = out_uop_0_valid; // @[Prf.scala 79:10]
  assign io_out_0_pc = out_uop_0_pc; // @[Prf.scala 79:10]
  assign io_out_0_npc = out_uop_0_npc; // @[Prf.scala 79:10]
  assign io_out_0_inst = out_uop_0_inst; // @[Prf.scala 79:10]
  assign io_out_0_fu_code = out_uop_0_fu_code; // @[Prf.scala 79:10]
  assign io_out_0_alu_code = out_uop_0_alu_code; // @[Prf.scala 79:10]
  assign io_out_0_jmp_code = out_uop_0_jmp_code; // @[Prf.scala 79:10]
  assign io_out_0_sys_code = out_uop_0_sys_code; // @[Prf.scala 79:10]
  assign io_out_0_w_type = out_uop_0_w_type; // @[Prf.scala 79:10]
  assign io_out_0_rs1_src = out_uop_0_rs1_src; // @[Prf.scala 79:10]
  assign io_out_0_rs2_src = out_uop_0_rs2_src; // @[Prf.scala 79:10]
  assign io_out_0_rd_en = out_uop_0_rd_en; // @[Prf.scala 79:10]
  assign io_out_0_imm = out_uop_0_imm; // @[Prf.scala 79:10]
  assign io_out_0_pred_br = out_uop_0_pred_br; // @[Prf.scala 79:10]
  assign io_out_0_pred_bpc = out_uop_0_pred_bpc; // @[Prf.scala 79:10]
  assign io_out_0_rd_paddr = out_uop_0_rd_paddr; // @[Prf.scala 79:10]
  assign io_out_0_rob_addr = out_uop_0_rob_addr; // @[Prf.scala 79:10]
  assign io_out_1_valid = out_uop_1_valid; // @[Prf.scala 79:10]
  assign io_out_1_pc = out_uop_1_pc; // @[Prf.scala 79:10]
  assign io_out_1_npc = out_uop_1_npc; // @[Prf.scala 79:10]
  assign io_out_1_fu_code = out_uop_1_fu_code; // @[Prf.scala 79:10]
  assign io_out_1_alu_code = out_uop_1_alu_code; // @[Prf.scala 79:10]
  assign io_out_1_jmp_code = out_uop_1_jmp_code; // @[Prf.scala 79:10]
  assign io_out_1_w_type = out_uop_1_w_type; // @[Prf.scala 79:10]
  assign io_out_1_rs1_src = out_uop_1_rs1_src; // @[Prf.scala 79:10]
  assign io_out_1_rs2_src = out_uop_1_rs2_src; // @[Prf.scala 79:10]
  assign io_out_1_rd_en = out_uop_1_rd_en; // @[Prf.scala 79:10]
  assign io_out_1_imm = out_uop_1_imm; // @[Prf.scala 79:10]
  assign io_out_1_pred_br = out_uop_1_pred_br; // @[Prf.scala 79:10]
  assign io_out_1_pred_bpc = out_uop_1_pred_bpc; // @[Prf.scala 79:10]
  assign io_out_1_rd_paddr = out_uop_1_rd_paddr; // @[Prf.scala 79:10]
  assign io_out_1_rob_addr = out_uop_1_rob_addr; // @[Prf.scala 79:10]
  assign io_out_2_valid = out_uop_2_valid; // @[Prf.scala 79:10]
  assign io_out_2_pc = out_uop_2_pc; // @[Prf.scala 79:10]
  assign io_out_2_fu_code = out_uop_2_fu_code; // @[Prf.scala 79:10]
  assign io_out_2_alu_code = out_uop_2_alu_code; // @[Prf.scala 79:10]
  assign io_out_2_mem_code = out_uop_2_mem_code; // @[Prf.scala 79:10]
  assign io_out_2_mem_size = out_uop_2_mem_size; // @[Prf.scala 79:10]
  assign io_out_2_w_type = out_uop_2_w_type; // @[Prf.scala 79:10]
  assign io_out_2_rs1_src = out_uop_2_rs1_src; // @[Prf.scala 79:10]
  assign io_out_2_rs2_src = out_uop_2_rs2_src; // @[Prf.scala 79:10]
  assign io_out_2_rd_en = out_uop_2_rd_en; // @[Prf.scala 79:10]
  assign io_out_2_imm = out_uop_2_imm; // @[Prf.scala 79:10]
  assign io_out_2_rd_paddr = out_uop_2_rd_paddr; // @[Prf.scala 79:10]
  assign io_out_2_rob_addr = out_uop_2_rob_addr; // @[Prf.scala 79:10]
  assign io_rs1_data_0 = out_rs1_data_0; // @[Prf.scala 80:15]
  assign io_rs1_data_1 = out_rs1_data_1; // @[Prf.scala 80:15]
  assign io_rs1_data_2 = out_rs1_data_2; // @[Prf.scala 80:15]
  assign io_rs2_data_0 = out_rs2_data_0; // @[Prf.scala 81:15]
  assign io_rs2_data_1 = out_rs2_data_1; // @[Prf.scala 81:15]
  assign io_rs2_data_2 = out_rs2_data_2; // @[Prf.scala 81:15]
  always @(posedge clock) begin
    if (prf_MPORT_en & prf_MPORT_mask) begin
      prf[prf_MPORT_addr] <= prf_MPORT_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_1_en & prf_MPORT_1_mask) begin
      prf[prf_MPORT_1_addr] <= prf_MPORT_1_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_2_en & prf_MPORT_2_mask) begin
      prf[prf_MPORT_2_addr] <= prf_MPORT_2_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_9_en & prf_MPORT_9_mask) begin
      prf[prf_MPORT_9_addr] <= prf_MPORT_9_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_10_en & prf_MPORT_10_mask) begin
      prf[prf_MPORT_10_addr] <= prf_MPORT_10_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_11_en & prf_MPORT_11_mask) begin
      prf[prf_MPORT_11_addr] <= prf_MPORT_11_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_12_en & prf_MPORT_12_mask) begin
      prf[prf_MPORT_12_addr] <= prf_MPORT_12_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_13_en & prf_MPORT_13_mask) begin
      prf[prf_MPORT_13_addr] <= prf_MPORT_13_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_14_en & prf_MPORT_14_mask) begin
      prf[prf_MPORT_14_addr] <= prf_MPORT_14_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_15_en & prf_MPORT_15_mask) begin
      prf[prf_MPORT_15_addr] <= prf_MPORT_15_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_16_en & prf_MPORT_16_mask) begin
      prf[prf_MPORT_16_addr] <= prf_MPORT_16_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_17_en & prf_MPORT_17_mask) begin
      prf[prf_MPORT_17_addr] <= prf_MPORT_17_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_18_en & prf_MPORT_18_mask) begin
      prf[prf_MPORT_18_addr] <= prf_MPORT_18_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_19_en & prf_MPORT_19_mask) begin
      prf[prf_MPORT_19_addr] <= prf_MPORT_19_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_20_en & prf_MPORT_20_mask) begin
      prf[prf_MPORT_20_addr] <= prf_MPORT_20_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_21_en & prf_MPORT_21_mask) begin
      prf[prf_MPORT_21_addr] <= prf_MPORT_21_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_22_en & prf_MPORT_22_mask) begin
      prf[prf_MPORT_22_addr] <= prf_MPORT_22_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_23_en & prf_MPORT_23_mask) begin
      prf[prf_MPORT_23_addr] <= prf_MPORT_23_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_24_en & prf_MPORT_24_mask) begin
      prf[prf_MPORT_24_addr] <= prf_MPORT_24_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_25_en & prf_MPORT_25_mask) begin
      prf[prf_MPORT_25_addr] <= prf_MPORT_25_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_26_en & prf_MPORT_26_mask) begin
      prf[prf_MPORT_26_addr] <= prf_MPORT_26_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_27_en & prf_MPORT_27_mask) begin
      prf[prf_MPORT_27_addr] <= prf_MPORT_27_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_28_en & prf_MPORT_28_mask) begin
      prf[prf_MPORT_28_addr] <= prf_MPORT_28_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_29_en & prf_MPORT_29_mask) begin
      prf[prf_MPORT_29_addr] <= prf_MPORT_29_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_30_en & prf_MPORT_30_mask) begin
      prf[prf_MPORT_30_addr] <= prf_MPORT_30_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_31_en & prf_MPORT_31_mask) begin
      prf[prf_MPORT_31_addr] <= prf_MPORT_31_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_32_en & prf_MPORT_32_mask) begin
      prf[prf_MPORT_32_addr] <= prf_MPORT_32_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_33_en & prf_MPORT_33_mask) begin
      prf[prf_MPORT_33_addr] <= prf_MPORT_33_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_34_en & prf_MPORT_34_mask) begin
      prf[prf_MPORT_34_addr] <= prf_MPORT_34_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_35_en & prf_MPORT_35_mask) begin
      prf[prf_MPORT_35_addr] <= prf_MPORT_35_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_36_en & prf_MPORT_36_mask) begin
      prf[prf_MPORT_36_addr] <= prf_MPORT_36_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_37_en & prf_MPORT_37_mask) begin
      prf[prf_MPORT_37_addr] <= prf_MPORT_37_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_38_en & prf_MPORT_38_mask) begin
      prf[prf_MPORT_38_addr] <= prf_MPORT_38_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_39_en & prf_MPORT_39_mask) begin
      prf[prf_MPORT_39_addr] <= prf_MPORT_39_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_40_en & prf_MPORT_40_mask) begin
      prf[prf_MPORT_40_addr] <= prf_MPORT_40_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_41_en & prf_MPORT_41_mask) begin
      prf[prf_MPORT_41_addr] <= prf_MPORT_41_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_42_en & prf_MPORT_42_mask) begin
      prf[prf_MPORT_42_addr] <= prf_MPORT_42_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_43_en & prf_MPORT_43_mask) begin
      prf[prf_MPORT_43_addr] <= prf_MPORT_43_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_44_en & prf_MPORT_44_mask) begin
      prf[prf_MPORT_44_addr] <= prf_MPORT_44_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_45_en & prf_MPORT_45_mask) begin
      prf[prf_MPORT_45_addr] <= prf_MPORT_45_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_46_en & prf_MPORT_46_mask) begin
      prf[prf_MPORT_46_addr] <= prf_MPORT_46_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_47_en & prf_MPORT_47_mask) begin
      prf[prf_MPORT_47_addr] <= prf_MPORT_47_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_48_en & prf_MPORT_48_mask) begin
      prf[prf_MPORT_48_addr] <= prf_MPORT_48_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_49_en & prf_MPORT_49_mask) begin
      prf[prf_MPORT_49_addr] <= prf_MPORT_49_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_50_en & prf_MPORT_50_mask) begin
      prf[prf_MPORT_50_addr] <= prf_MPORT_50_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_51_en & prf_MPORT_51_mask) begin
      prf[prf_MPORT_51_addr] <= prf_MPORT_51_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_52_en & prf_MPORT_52_mask) begin
      prf[prf_MPORT_52_addr] <= prf_MPORT_52_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_53_en & prf_MPORT_53_mask) begin
      prf[prf_MPORT_53_addr] <= prf_MPORT_53_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_54_en & prf_MPORT_54_mask) begin
      prf[prf_MPORT_54_addr] <= prf_MPORT_54_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_55_en & prf_MPORT_55_mask) begin
      prf[prf_MPORT_55_addr] <= prf_MPORT_55_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_56_en & prf_MPORT_56_mask) begin
      prf[prf_MPORT_56_addr] <= prf_MPORT_56_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_57_en & prf_MPORT_57_mask) begin
      prf[prf_MPORT_57_addr] <= prf_MPORT_57_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_58_en & prf_MPORT_58_mask) begin
      prf[prf_MPORT_58_addr] <= prf_MPORT_58_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_59_en & prf_MPORT_59_mask) begin
      prf[prf_MPORT_59_addr] <= prf_MPORT_59_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_60_en & prf_MPORT_60_mask) begin
      prf[prf_MPORT_60_addr] <= prf_MPORT_60_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_61_en & prf_MPORT_61_mask) begin
      prf[prf_MPORT_61_addr] <= prf_MPORT_61_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_62_en & prf_MPORT_62_mask) begin
      prf[prf_MPORT_62_addr] <= prf_MPORT_62_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_63_en & prf_MPORT_63_mask) begin
      prf[prf_MPORT_63_addr] <= prf_MPORT_63_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_64_en & prf_MPORT_64_mask) begin
      prf[prf_MPORT_64_addr] <= prf_MPORT_64_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_65_en & prf_MPORT_65_mask) begin
      prf[prf_MPORT_65_addr] <= prf_MPORT_65_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_66_en & prf_MPORT_66_mask) begin
      prf[prf_MPORT_66_addr] <= prf_MPORT_66_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_67_en & prf_MPORT_67_mask) begin
      prf[prf_MPORT_67_addr] <= prf_MPORT_67_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_68_en & prf_MPORT_68_mask) begin
      prf[prf_MPORT_68_addr] <= prf_MPORT_68_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_69_en & prf_MPORT_69_mask) begin
      prf[prf_MPORT_69_addr] <= prf_MPORT_69_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_70_en & prf_MPORT_70_mask) begin
      prf[prf_MPORT_70_addr] <= prf_MPORT_70_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_71_en & prf_MPORT_71_mask) begin
      prf[prf_MPORT_71_addr] <= prf_MPORT_71_data; // @[Prf.scala 20:16]
    end
    if (prf_MPORT_72_en & prf_MPORT_72_mask) begin
      prf[prf_MPORT_72_addr] <= prf_MPORT_72_data; // @[Prf.scala 20:16]
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_valid <= 1'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_valid <= 1'h0; // @[Prf.scala 67:18]
    end else begin
      out_uop_0_valid <= io_in_0_valid; // @[Prf.scala 73:18]
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_pc <= 32'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_pc <= 32'h0; // @[Prf.scala 67:18]
    end else if (io_in_0_valid) begin // @[Prf.scala 73:24]
      out_uop_0_pc <= io_in_0_pc;
    end else begin
      out_uop_0_pc <= 32'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_npc <= 32'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_npc <= 32'h0; // @[Prf.scala 67:18]
    end else if (io_in_0_valid) begin // @[Prf.scala 73:24]
      out_uop_0_npc <= io_in_0_npc;
    end else begin
      out_uop_0_npc <= 32'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_inst <= 32'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_inst <= 32'h0; // @[Prf.scala 67:18]
    end else if (io_in_0_valid) begin // @[Prf.scala 73:24]
      out_uop_0_inst <= io_in_0_inst;
    end else begin
      out_uop_0_inst <= 32'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_fu_code <= 3'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_fu_code <= 3'h0; // @[Prf.scala 67:18]
    end else if (io_in_0_valid) begin // @[Prf.scala 73:24]
      out_uop_0_fu_code <= io_in_0_fu_code;
    end else begin
      out_uop_0_fu_code <= 3'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_alu_code <= 4'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_alu_code <= 4'h0; // @[Prf.scala 67:18]
    end else if (io_in_0_valid) begin // @[Prf.scala 73:24]
      out_uop_0_alu_code <= io_in_0_alu_code;
    end else begin
      out_uop_0_alu_code <= 4'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_jmp_code <= 4'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_jmp_code <= 4'h0; // @[Prf.scala 67:18]
    end else if (io_in_0_valid) begin // @[Prf.scala 73:24]
      out_uop_0_jmp_code <= io_in_0_jmp_code;
    end else begin
      out_uop_0_jmp_code <= 4'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_sys_code <= 3'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_sys_code <= 3'h0; // @[Prf.scala 67:18]
    end else if (io_in_0_valid) begin // @[Prf.scala 73:24]
      out_uop_0_sys_code <= io_in_0_sys_code;
    end else begin
      out_uop_0_sys_code <= 3'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_w_type <= 1'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_w_type <= 1'h0; // @[Prf.scala 67:18]
    end else begin
      out_uop_0_w_type <= io_in_0_valid & io_in_0_w_type; // @[Prf.scala 73:18]
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_rs1_src <= 2'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_rs1_src <= 2'h0; // @[Prf.scala 67:18]
    end else if (io_in_0_valid) begin // @[Prf.scala 73:24]
      out_uop_0_rs1_src <= io_in_0_rs1_src;
    end else begin
      out_uop_0_rs1_src <= 2'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_rs2_src <= 2'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_rs2_src <= 2'h0; // @[Prf.scala 67:18]
    end else if (io_in_0_valid) begin // @[Prf.scala 73:24]
      out_uop_0_rs2_src <= io_in_0_rs2_src;
    end else begin
      out_uop_0_rs2_src <= 2'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_rd_en <= 1'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_rd_en <= 1'h0; // @[Prf.scala 67:18]
    end else begin
      out_uop_0_rd_en <= io_in_0_valid & io_in_0_rd_en; // @[Prf.scala 73:18]
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_imm <= 32'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_imm <= 32'h0; // @[Prf.scala 67:18]
    end else if (io_in_0_valid) begin // @[Prf.scala 73:24]
      out_uop_0_imm <= io_in_0_imm;
    end else begin
      out_uop_0_imm <= 32'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_pred_br <= 1'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_pred_br <= 1'h0; // @[Prf.scala 67:18]
    end else begin
      out_uop_0_pred_br <= io_in_0_valid & io_in_0_pred_br; // @[Prf.scala 73:18]
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_pred_bpc <= 32'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_pred_bpc <= 32'h0; // @[Prf.scala 67:18]
    end else if (io_in_0_valid) begin // @[Prf.scala 73:24]
      out_uop_0_pred_bpc <= io_in_0_pred_bpc;
    end else begin
      out_uop_0_pred_bpc <= 32'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_rd_paddr <= 6'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_rd_paddr <= 6'h0; // @[Prf.scala 67:18]
    end else if (io_in_0_valid) begin // @[Prf.scala 73:24]
      out_uop_0_rd_paddr <= io_in_0_rd_paddr;
    end else begin
      out_uop_0_rd_paddr <= 6'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_0_rob_addr <= 4'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_0_rob_addr <= 4'h0; // @[Prf.scala 67:18]
    end else if (io_in_0_valid) begin // @[Prf.scala 73:24]
      out_uop_0_rob_addr <= io_in_0_rob_addr;
    end else begin
      out_uop_0_rob_addr <= 4'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_valid <= 1'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_valid <= 1'h0; // @[Prf.scala 67:18]
    end else begin
      out_uop_1_valid <= io_in_1_valid; // @[Prf.scala 73:18]
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_pc <= 32'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_pc <= 32'h0; // @[Prf.scala 67:18]
    end else if (io_in_1_valid) begin // @[Prf.scala 73:24]
      out_uop_1_pc <= io_in_1_pc;
    end else begin
      out_uop_1_pc <= 32'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_npc <= 32'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_npc <= 32'h0; // @[Prf.scala 67:18]
    end else if (io_in_1_valid) begin // @[Prf.scala 73:24]
      out_uop_1_npc <= io_in_1_npc;
    end else begin
      out_uop_1_npc <= 32'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_fu_code <= 3'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_fu_code <= 3'h0; // @[Prf.scala 67:18]
    end else if (io_in_1_valid) begin // @[Prf.scala 73:24]
      out_uop_1_fu_code <= io_in_1_fu_code;
    end else begin
      out_uop_1_fu_code <= 3'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_alu_code <= 4'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_alu_code <= 4'h0; // @[Prf.scala 67:18]
    end else if (io_in_1_valid) begin // @[Prf.scala 73:24]
      out_uop_1_alu_code <= io_in_1_alu_code;
    end else begin
      out_uop_1_alu_code <= 4'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_jmp_code <= 4'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_jmp_code <= 4'h0; // @[Prf.scala 67:18]
    end else if (io_in_1_valid) begin // @[Prf.scala 73:24]
      out_uop_1_jmp_code <= io_in_1_jmp_code;
    end else begin
      out_uop_1_jmp_code <= 4'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_w_type <= 1'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_w_type <= 1'h0; // @[Prf.scala 67:18]
    end else begin
      out_uop_1_w_type <= io_in_1_valid & io_in_1_w_type; // @[Prf.scala 73:18]
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_rs1_src <= 2'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_rs1_src <= 2'h0; // @[Prf.scala 67:18]
    end else if (io_in_1_valid) begin // @[Prf.scala 73:24]
      out_uop_1_rs1_src <= io_in_1_rs1_src;
    end else begin
      out_uop_1_rs1_src <= 2'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_rs2_src <= 2'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_rs2_src <= 2'h0; // @[Prf.scala 67:18]
    end else if (io_in_1_valid) begin // @[Prf.scala 73:24]
      out_uop_1_rs2_src <= io_in_1_rs2_src;
    end else begin
      out_uop_1_rs2_src <= 2'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_rd_en <= 1'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_rd_en <= 1'h0; // @[Prf.scala 67:18]
    end else begin
      out_uop_1_rd_en <= io_in_1_valid & io_in_1_rd_en; // @[Prf.scala 73:18]
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_imm <= 32'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_imm <= 32'h0; // @[Prf.scala 67:18]
    end else if (io_in_1_valid) begin // @[Prf.scala 73:24]
      out_uop_1_imm <= io_in_1_imm;
    end else begin
      out_uop_1_imm <= 32'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_pred_br <= 1'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_pred_br <= 1'h0; // @[Prf.scala 67:18]
    end else begin
      out_uop_1_pred_br <= io_in_1_valid & io_in_1_pred_br; // @[Prf.scala 73:18]
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_pred_bpc <= 32'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_pred_bpc <= 32'h0; // @[Prf.scala 67:18]
    end else if (io_in_1_valid) begin // @[Prf.scala 73:24]
      out_uop_1_pred_bpc <= io_in_1_pred_bpc;
    end else begin
      out_uop_1_pred_bpc <= 32'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_rd_paddr <= 6'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_rd_paddr <= 6'h0; // @[Prf.scala 67:18]
    end else if (io_in_1_valid) begin // @[Prf.scala 73:24]
      out_uop_1_rd_paddr <= io_in_1_rd_paddr;
    end else begin
      out_uop_1_rd_paddr <= 6'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_1_rob_addr <= 4'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_1_rob_addr <= 4'h0; // @[Prf.scala 67:18]
    end else if (io_in_1_valid) begin // @[Prf.scala 73:24]
      out_uop_1_rob_addr <= io_in_1_rob_addr;
    end else begin
      out_uop_1_rob_addr <= 4'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_2_valid <= 1'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_2_valid <= 1'h0; // @[Prf.scala 67:18]
    end else begin
      out_uop_2_valid <= io_in_2_valid; // @[Prf.scala 73:18]
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_2_pc <= 32'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_2_pc <= 32'h0; // @[Prf.scala 67:18]
    end else if (io_in_2_valid) begin // @[Prf.scala 73:24]
      out_uop_2_pc <= io_in_2_pc;
    end else begin
      out_uop_2_pc <= 32'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_2_fu_code <= 3'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_2_fu_code <= 3'h0; // @[Prf.scala 67:18]
    end else if (io_in_2_valid) begin // @[Prf.scala 73:24]
      out_uop_2_fu_code <= io_in_2_fu_code;
    end else begin
      out_uop_2_fu_code <= 3'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_2_alu_code <= 4'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_2_alu_code <= 4'h0; // @[Prf.scala 67:18]
    end else if (io_in_2_valid) begin // @[Prf.scala 73:24]
      out_uop_2_alu_code <= io_in_2_alu_code;
    end else begin
      out_uop_2_alu_code <= 4'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_2_mem_code <= 2'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_2_mem_code <= 2'h0; // @[Prf.scala 67:18]
    end else if (io_in_2_valid) begin // @[Prf.scala 73:24]
      out_uop_2_mem_code <= io_in_2_mem_code;
    end else begin
      out_uop_2_mem_code <= 2'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_2_mem_size <= 2'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_2_mem_size <= 2'h0; // @[Prf.scala 67:18]
    end else if (io_in_2_valid) begin // @[Prf.scala 73:24]
      out_uop_2_mem_size <= io_in_2_mem_size;
    end else begin
      out_uop_2_mem_size <= 2'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_2_w_type <= 1'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_2_w_type <= 1'h0; // @[Prf.scala 67:18]
    end else begin
      out_uop_2_w_type <= io_in_2_valid & io_in_2_w_type; // @[Prf.scala 73:18]
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_2_rs1_src <= 2'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_2_rs1_src <= 2'h0; // @[Prf.scala 67:18]
    end else if (io_in_2_valid) begin // @[Prf.scala 73:24]
      out_uop_2_rs1_src <= io_in_2_rs1_src;
    end else begin
      out_uop_2_rs1_src <= 2'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_2_rs2_src <= 2'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_2_rs2_src <= 2'h0; // @[Prf.scala 67:18]
    end else if (io_in_2_valid) begin // @[Prf.scala 73:24]
      out_uop_2_rs2_src <= io_in_2_rs2_src;
    end else begin
      out_uop_2_rs2_src <= 2'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_2_rd_en <= 1'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_2_rd_en <= 1'h0; // @[Prf.scala 67:18]
    end else begin
      out_uop_2_rd_en <= io_in_2_valid & io_in_2_rd_en; // @[Prf.scala 73:18]
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_2_imm <= 32'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_2_imm <= 32'h0; // @[Prf.scala 67:18]
    end else if (io_in_2_valid) begin // @[Prf.scala 73:24]
      out_uop_2_imm <= io_in_2_imm;
    end else begin
      out_uop_2_imm <= 32'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_2_rd_paddr <= 6'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_2_rd_paddr <= 6'h0; // @[Prf.scala 67:18]
    end else if (io_in_2_valid) begin // @[Prf.scala 73:24]
      out_uop_2_rd_paddr <= io_in_2_rd_paddr;
    end else begin
      out_uop_2_rd_paddr <= 6'h0;
    end
    if (reset) begin // @[Prf.scala 60:24]
      out_uop_2_rob_addr <= 4'h0; // @[Prf.scala 60:24]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_uop_2_rob_addr <= 4'h0; // @[Prf.scala 67:18]
    end else if (io_in_2_valid) begin // @[Prf.scala 73:24]
      out_uop_2_rob_addr <= io_in_2_rob_addr;
    end else begin
      out_uop_2_rob_addr <= 4'h0;
    end
    if (reset) begin // @[Prf.scala 61:29]
      out_rs1_data_0 <= 64'h0; // @[Prf.scala 61:29]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_rs1_data_0 <= 64'h0; // @[Prf.scala 68:23]
    end else if (_T_3) begin // @[Prf.scala 41:54]
      if (io_rd_paddr_1 == io_in_0_rs1_paddr) begin // @[Prf.scala 42:48]
        out_rs1_data_0 <= io_rd_data_1; // @[Prf.scala 43:23]
      end else begin
        out_rs1_data_0 <= _GEN_17;
      end
    end else begin
      out_rs1_data_0 <= _GEN_17;
    end
    if (reset) begin // @[Prf.scala 61:29]
      out_rs1_data_1 <= 64'h0; // @[Prf.scala 61:29]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_rs1_data_1 <= 64'h0; // @[Prf.scala 68:23]
    end else if (_T_3) begin // @[Prf.scala 41:54]
      if (io_rd_paddr_1 == io_in_1_rs1_paddr) begin // @[Prf.scala 42:48]
        out_rs1_data_1 <= io_rd_data_1; // @[Prf.scala 43:23]
      end else begin
        out_rs1_data_1 <= _GEN_25;
      end
    end else begin
      out_rs1_data_1 <= _GEN_25;
    end
    if (reset) begin // @[Prf.scala 61:29]
      out_rs1_data_2 <= 64'h0; // @[Prf.scala 61:29]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_rs1_data_2 <= 64'h0; // @[Prf.scala 68:23]
    end else if (_T_3) begin // @[Prf.scala 41:54]
      if (io_rd_paddr_1 == io_in_2_rs1_paddr) begin // @[Prf.scala 42:48]
        out_rs1_data_2 <= io_rd_data_1; // @[Prf.scala 43:23]
      end else begin
        out_rs1_data_2 <= _GEN_33;
      end
    end else begin
      out_rs1_data_2 <= _GEN_33;
    end
    if (reset) begin // @[Prf.scala 62:29]
      out_rs2_data_0 <= 64'h0; // @[Prf.scala 62:29]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_rs2_data_0 <= 64'h0; // @[Prf.scala 69:23]
    end else if (_T_3) begin // @[Prf.scala 41:54]
      if (io_rd_paddr_1 == io_in_0_rs2_paddr) begin // @[Prf.scala 45:48]
        out_rs2_data_0 <= io_rd_data_1; // @[Prf.scala 46:23]
      end else begin
        out_rs2_data_0 <= _GEN_18;
      end
    end else begin
      out_rs2_data_0 <= _GEN_18;
    end
    if (reset) begin // @[Prf.scala 62:29]
      out_rs2_data_1 <= 64'h0; // @[Prf.scala 62:29]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_rs2_data_1 <= 64'h0; // @[Prf.scala 69:23]
    end else if (_T_3) begin // @[Prf.scala 41:54]
      if (io_rd_paddr_1 == io_in_1_rs2_paddr) begin // @[Prf.scala 45:48]
        out_rs2_data_1 <= io_rd_data_1; // @[Prf.scala 46:23]
      end else begin
        out_rs2_data_1 <= _GEN_26;
      end
    end else begin
      out_rs2_data_1 <= _GEN_26;
    end
    if (reset) begin // @[Prf.scala 62:29]
      out_rs2_data_2 <= 64'h0; // @[Prf.scala 62:29]
    end else if (io_flush) begin // @[Prf.scala 65:19]
      out_rs2_data_2 <= 64'h0; // @[Prf.scala 69:23]
    end else if (_T_3) begin // @[Prf.scala 41:54]
      if (io_rd_paddr_1 == io_in_2_rs2_paddr) begin // @[Prf.scala 45:48]
        out_rs2_data_2 <= io_rd_data_1; // @[Prf.scala 46:23]
      end else begin
        out_rs2_data_2 <= _GEN_34;
      end
    end else begin
      out_rs2_data_2 <= _GEN_34;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    prf[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_uop_0_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_uop_0_pc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  out_uop_0_npc = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  out_uop_0_inst = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  out_uop_0_fu_code = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  out_uop_0_alu_code = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  out_uop_0_jmp_code = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  out_uop_0_sys_code = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  out_uop_0_w_type = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  out_uop_0_rs1_src = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  out_uop_0_rs2_src = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  out_uop_0_rd_en = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  out_uop_0_imm = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  out_uop_0_pred_br = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  out_uop_0_pred_bpc = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  out_uop_0_rd_paddr = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  out_uop_0_rob_addr = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  out_uop_1_valid = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  out_uop_1_pc = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  out_uop_1_npc = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  out_uop_1_fu_code = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  out_uop_1_alu_code = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  out_uop_1_jmp_code = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  out_uop_1_w_type = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  out_uop_1_rs1_src = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  out_uop_1_rs2_src = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  out_uop_1_rd_en = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  out_uop_1_imm = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  out_uop_1_pred_br = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  out_uop_1_pred_bpc = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  out_uop_1_rd_paddr = _RAND_31[5:0];
  _RAND_32 = {1{`RANDOM}};
  out_uop_1_rob_addr = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  out_uop_2_valid = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  out_uop_2_pc = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  out_uop_2_fu_code = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  out_uop_2_alu_code = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  out_uop_2_mem_code = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  out_uop_2_mem_size = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  out_uop_2_w_type = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  out_uop_2_rs1_src = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  out_uop_2_rs2_src = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  out_uop_2_rd_en = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  out_uop_2_imm = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  out_uop_2_rd_paddr = _RAND_44[5:0];
  _RAND_45 = {1{`RANDOM}};
  out_uop_2_rob_addr = _RAND_45[3:0];
  _RAND_46 = {2{`RANDOM}};
  out_rs1_data_0 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  out_rs1_data_1 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  out_rs1_data_2 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  out_rs2_data_0 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  out_rs2_data_1 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  out_rs2_data_2 = _RAND_51[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_Alu(
  input  [31:0] io_uop_pc,
  input  [31:0] io_uop_npc,
  input  [2:0]  io_uop_fu_code,
  input  [3:0]  io_uop_alu_code,
  input  [3:0]  io_uop_jmp_code,
  input         io_uop_w_type,
  input  [31:0] io_uop_imm,
  input         io_uop_pred_br,
  input  [31:0] io_uop_pred_bpc,
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output        io_ecp_jmp_valid,
  output        io_ecp_jmp,
  output [31:0] io_ecp_jmp_pc,
  output        io_ecp_mis,
  output [63:0] io_ecp_rd_data
);
  wire [5:0] shamt = io_uop_w_type ? {{1'd0}, io_in2[4:0]} : io_in2[5:0]; // @[Alu.scala 20:15]
  wire [63:0] _T_4 = io_in1 + io_in2; // @[Alu.scala 28:29]
  wire [63:0] _T_6 = io_in1 - io_in2; // @[Alu.scala 29:29]
  wire  _T_9 = $signed(io_in1) < $signed(io_in2); // @[Alu.scala 30:38]
  wire  _T_10 = io_in1 < io_in2; // @[Alu.scala 31:29]
  wire [63:0] _T_11 = io_in1 ^ io_in2; // @[Alu.scala 32:29]
  wire [63:0] _T_12 = io_in1 | io_in2; // @[Alu.scala 33:29]
  wire [63:0] _T_13 = io_in1 & io_in2; // @[Alu.scala 34:29]
  wire [126:0] _GEN_0 = {{63'd0}, io_in1}; // @[Alu.scala 35:30]
  wire [126:0] _T_14 = _GEN_0 << shamt; // @[Alu.scala 35:30]
  wire [63:0] _T_16 = io_in1 >> shamt; // @[Alu.scala 36:38]
  wire [63:0] _T_19 = $signed(io_in1) >>> shamt; // @[Alu.scala 37:54]
  wire [63:0] _T_21 = 4'h1 == io_uop_alu_code ? _T_4 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _T_23 = 4'h2 == io_uop_alu_code ? _T_6 : _T_21; // @[Mux.scala 80:57]
  wire [63:0] _T_25 = 4'h3 == io_uop_alu_code ? {{63'd0}, _T_9} : _T_23; // @[Mux.scala 80:57]
  wire [63:0] _T_27 = 4'h4 == io_uop_alu_code ? {{63'd0}, _T_10} : _T_25; // @[Mux.scala 80:57]
  wire [63:0] _T_29 = 4'h5 == io_uop_alu_code ? _T_11 : _T_27; // @[Mux.scala 80:57]
  wire [63:0] _T_31 = 4'h6 == io_uop_alu_code ? _T_12 : _T_29; // @[Mux.scala 80:57]
  wire [63:0] _T_33 = 4'h7 == io_uop_alu_code ? _T_13 : _T_31; // @[Mux.scala 80:57]
  wire [63:0] _T_35 = 4'h8 == io_uop_alu_code ? _T_14[63:0] : _T_33; // @[Mux.scala 80:57]
  wire [63:0] _T_37 = 4'h9 == io_uop_alu_code ? _T_16 : _T_35; // @[Mux.scala 80:57]
  wire [63:0] alu_out_0 = 4'ha == io_uop_alu_code ? _T_19 : _T_37; // @[Mux.scala 80:57]
  wire [31:0] _T_43 = alu_out_0[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_44 = {_T_43,alu_out_0[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] alu_out = io_uop_w_type ? _T_44 : alu_out_0; // @[Alu.scala 40:17]
  wire  _T_46 = io_in1 == io_in2; // @[Alu.scala 45:29]
  wire  _T_47 = io_in1 != io_in2; // @[Alu.scala 46:29]
  wire  _T_53 = $signed(io_in1) >= $signed(io_in2); // @[Alu.scala 48:38]
  wire  _T_55 = io_in1 >= io_in2; // @[Alu.scala 50:38]
  wire  _T_61 = 4'h3 == io_uop_jmp_code ? _T_46 : 4'h2 == io_uop_jmp_code | 4'h1 == io_uop_jmp_code; // @[Mux.scala 80:57]
  wire  _T_63 = 4'h4 == io_uop_jmp_code ? _T_47 : _T_61; // @[Mux.scala 80:57]
  wire  _T_65 = 4'h5 == io_uop_jmp_code ? _T_9 : _T_63; // @[Mux.scala 80:57]
  wire  _T_67 = 4'h6 == io_uop_jmp_code ? _T_53 : _T_65; // @[Mux.scala 80:57]
  wire  _T_69 = 4'h7 == io_uop_jmp_code ? _T_10 : _T_67; // @[Mux.scala 80:57]
  wire  jmp = 4'h8 == io_uop_jmp_code ? _T_55 : _T_69; // @[Mux.scala 80:57]
  wire [31:0] _T_74 = io_uop_jmp_code == 4'h2 ? io_in1[31:0] : io_uop_pc; // @[Alu.scala 53:16]
  wire [31:0] jmp_pc = _T_74 + io_uop_imm; // @[Alu.scala 53:71]
  wire [63:0] _T_78 = {32'h0,io_uop_npc}; // @[Cat.scala 30:58]
  wire [63:0] _T_82 = 4'h1 == io_uop_jmp_code ? _T_78 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] npc_to_rd = 4'h2 == io_uop_jmp_code ? _T_78 : _T_82; // @[Mux.scala 80:57]
  wire  _T_89 = io_uop_pred_br & jmp_pc != io_uop_pred_bpc | ~io_uop_pred_br; // @[Alu.scala 66:64]
  assign io_ecp_jmp_valid = io_uop_fu_code == 3'h2; // @[Alu.scala 62:36]
  assign io_ecp_jmp = 4'h8 == io_uop_jmp_code ? _T_55 : _T_69; // @[Mux.scala 80:57]
  assign io_ecp_jmp_pc = _T_74 + io_uop_imm; // @[Alu.scala 53:71]
  assign io_ecp_mis = jmp ? _T_89 : io_uop_pred_br; // @[Alu.scala 65:20]
  assign io_ecp_rd_data = io_uop_fu_code == 3'h1 ? alu_out : npc_to_rd; // @[Alu.scala 68:24]
endmodule
module ysyx_210128_Csr(
  input         clock,
  input         reset,
  input  [31:0] io_uop_pc,
  input  [31:0] io_uop_inst,
  input  [2:0]  io_uop_sys_code,
  input         io_uop_pred_br,
  input  [31:0] io_uop_pred_bpc,
  input  [63:0] io_in1,
  output        io_ecp_jmp_valid,
  output        io_ecp_jmp,
  output [31:0] io_ecp_jmp_pc,
  output        io_ecp_mis,
  output [63:0] io_ecp_rd_data,
  output        mtip_0,
  input  [63:0] intr_mcause_0,
  input  [63:0] csr_minstret,
  input  [63:0] intr_mstatus_0,
  output [29:0] _T_6_0,
  output        _T_5_0,
  input         intr_0,
  input  [63:0] csr_mcycle,
  output [63:0] mstatus_0,
  input  [63:0] intr_mepc_0,
  input         csr_mip_mtip
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  _T_1 = io_uop_sys_code == 3'h2; // @[Csr.scala 34:26]
  wire  _T_2 = io_uop_sys_code == 3'h1 | _T_1; // @[Csr.scala 33:48]
  wire  _T_3 = io_uop_sys_code == 3'h3; // @[Csr.scala 35:26]
  wire  csr_rw = _T_2 | _T_3; // @[Csr.scala 34:48]
  reg [63:0] mhartid; // @[Csr.scala 41:26]
  reg [63:0] mstatus; // @[Csr.scala 42:26]
  reg [63:0] mie; // @[Csr.scala 43:26]
  reg [63:0] mtvec; // @[Csr.scala 44:26]
  reg [63:0] mscratch; // @[Csr.scala 45:26]
  reg [63:0] mepc; // @[Csr.scala 46:26]
  reg [63:0] mcause; // @[Csr.scala 47:26]
//   wire  _T_5 = mie[7]; // @[Csr.scala 50:28]
//   wire [29:0] _T_6 = mtvec[31:2]; // @[Csr.scala 51:30]
  wire  _T_7 = io_uop_sys_code == 3'h4; // @[Csr.scala 75:18]
  wire [63:0] _T_12 = {mstatus[63:8],mstatus[3],mstatus[6:4],1'h0,mstatus[2:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_15 = {mtvec[31:2],2'h0}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_2 = io_uop_sys_code == 3'h4 ? _T_12 : mstatus; // @[Csr.scala 75:40 78:13 42:26]
  wire [31:0] _GEN_4 = io_uop_sys_code == 3'h4 ? _T_15 : 32'h0; // @[Csr.scala 75:40 80:16]
  wire [63:0] _T_21 = {mstatus[63:8],1'h1,mstatus[6:4],mstatus[7],mstatus[2:0]}; // @[Cat.scala 30:58]
  wire  csr_jmp = io_uop_sys_code == 3'h5 | _T_7; // @[Csr.scala 84:39 86:13]
  wire [31:0] csr_jmp_pc = io_uop_sys_code == 3'h5 ? mepc[31:0] : _GEN_4; // @[Csr.scala 84:39 87:16]
  wire [11:0] addr = io_uop_inst[31:20]; // @[Csr.scala 124:22]
  wire  _T_113 = addr == 12'h300; // @[RegMap.scala 42:18]
  wire  _T_105 = addr == 12'hf14; // @[RegMap.scala 42:18]
  wire  _T_97 = addr == 12'h342; // @[RegMap.scala 42:18]
  wire  _T_89 = addr == 12'h340; // @[RegMap.scala 42:18]
  wire  _T_81 = addr == 12'h305; // @[RegMap.scala 42:18]
  wire  _T_73 = addr == 12'h341; // @[RegMap.scala 42:18]
  wire  _T_65 = addr == 12'h304; // @[RegMap.scala 42:18]
  wire [63:0] _GEN_11 = addr == 12'hb02 ? csr_minstret : 64'h0; // @[RegMap.scala 42:25 43:15]
  wire [63:0] _GEN_13 = addr == 12'hb00 ? csr_mcycle : _GEN_11; // @[RegMap.scala 42:25 43:15]
  wire [63:0] _GEN_15 = addr == 12'h304 ? mie : _GEN_13; // @[RegMap.scala 42:25 43:15]
  wire [63:0] _GEN_17 = addr == 12'h341 ? mepc : _GEN_15; // @[RegMap.scala 42:25 43:15]
  wire [63:0] _GEN_19 = addr == 12'h305 ? mtvec : _GEN_17; // @[RegMap.scala 42:25 43:15]
  wire [63:0] _GEN_21 = addr == 12'h340 ? mscratch : _GEN_19; // @[RegMap.scala 42:25 43:15]
  wire [63:0] _GEN_23 = addr == 12'h342 ? mcause : _GEN_21; // @[RegMap.scala 42:25 43:15]
  wire [63:0] _GEN_25 = addr == 12'hf14 ? mhartid : _GEN_23; // @[RegMap.scala 42:25 43:15]
  wire [63:0] _GEN_27 = addr == 12'h300 ? mstatus : _GEN_25; // @[RegMap.scala 42:25 43:15]
  wire [63:0] rdata = 12'h344 == addr ? 64'h0 : _GEN_27; // @[Csr.scala 138:28 139:11]
  wire [63:0] _T_40 = rdata | io_in1; // @[Csr.scala 131:32]
  wire [63:0] _T_41 = ~io_in1; // @[Csr.scala 132:34]
  wire [63:0] _T_42 = rdata & _T_41; // @[Csr.scala 132:32]
  wire [63:0] _T_44 = 3'h1 == io_uop_sys_code ? io_in1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _T_46 = 3'h2 == io_uop_sys_code ? _T_40 : _T_44; // @[Mux.scala 80:57]
  wire [63:0] wdata = 3'h3 == io_uop_sys_code ? _T_42 : _T_46; // @[Mux.scala 80:57]
  wire  _T_125 = wdata[16:15] == 2'h3 | wdata[14:13] == 2'h3; // @[Csr.scala 69:61]
  wire [63:0] _T_127 = {_T_125,wdata[62:0]}; // @[Cat.scala 30:58]
  wire  _T_132 = io_uop_pred_br & csr_jmp_pc != io_uop_pred_bpc | ~io_uop_pred_br; // @[Csr.scala 148:68]
  wire  mtip = csr_mip_mtip;
  assign io_ecp_jmp_valid = io_uop_sys_code == 3'h5 | _T_7; // @[Csr.scala 84:39 86:13]
  assign io_ecp_jmp = io_uop_sys_code == 3'h5 | _T_7; // @[Csr.scala 84:39 86:13]
  assign io_ecp_jmp_pc = io_uop_sys_code == 3'h5 ? mepc[31:0] : _GEN_4; // @[Csr.scala 84:39 87:16]
  assign io_ecp_mis = csr_jmp ? _T_132 : io_uop_pred_br; // @[Csr.scala 147:20]
  assign io_ecp_rd_data = 12'h344 == addr ? 64'h0 : _GEN_27; // @[Csr.scala 138:28 139:11]
  assign mtip_0 = mtip;
  assign _T_6_0 = mtvec[31:2];
  assign _T_5_0 = mie[7];
  assign mstatus_0 = mstatus;
  always @(posedge clock) begin
    if (reset) begin // @[Csr.scala 41:26]
      mhartid <= 64'h0; // @[Csr.scala 41:26]
    end else if (_T_105 & csr_rw) begin // @[RegMap.scala 46:34]
      if (3'h3 == io_uop_sys_code) begin // @[Mux.scala 80:57]
        mhartid <= _T_42;
      end else if (3'h2 == io_uop_sys_code) begin // @[Mux.scala 80:57]
        mhartid <= _T_40;
      end else begin
        mhartid <= _T_44;
      end
    end
    if (reset) begin // @[Csr.scala 42:26]
      mstatus <= 64'h1800; // @[Csr.scala 42:26]
    end else if (_T_113 & csr_rw) begin // @[RegMap.scala 46:34]
      mstatus <= _T_127; // @[RegMap.scala 47:13]
    end else if (intr_0) begin // @[Csr.scala 101:15]
      mstatus <= intr_mstatus_0; // @[Csr.scala 102:13]
    end else if (io_uop_sys_code == 3'h5) begin // @[Csr.scala 84:39]
      mstatus <= _T_21; // @[Csr.scala 85:13]
    end else begin
      mstatus <= _GEN_2;
    end
    if (reset) begin // @[Csr.scala 43:26]
      mie <= 64'h0; // @[Csr.scala 43:26]
    end else if (_T_65 & csr_rw) begin // @[RegMap.scala 46:34]
      if (3'h3 == io_uop_sys_code) begin // @[Mux.scala 80:57]
        mie <= _T_42;
      end else if (3'h2 == io_uop_sys_code) begin // @[Mux.scala 80:57]
        mie <= _T_40;
      end else begin
        mie <= _T_44;
      end
    end
    if (reset) begin // @[Csr.scala 44:26]
      mtvec <= 64'h0; // @[Csr.scala 44:26]
    end else if (_T_81 & csr_rw) begin // @[RegMap.scala 46:34]
      if (3'h3 == io_uop_sys_code) begin // @[Mux.scala 80:57]
        mtvec <= _T_42;
      end else if (3'h2 == io_uop_sys_code) begin // @[Mux.scala 80:57]
        mtvec <= _T_40;
      end else begin
        mtvec <= _T_44;
      end
    end
    if (reset) begin // @[Csr.scala 45:26]
      mscratch <= 64'h0; // @[Csr.scala 45:26]
    end else if (_T_89 & csr_rw) begin // @[RegMap.scala 46:34]
      if (3'h3 == io_uop_sys_code) begin // @[Mux.scala 80:57]
        mscratch <= _T_42;
      end else if (3'h2 == io_uop_sys_code) begin // @[Mux.scala 80:57]
        mscratch <= _T_40;
      end else begin
        mscratch <= _T_44;
      end
    end
    if (reset) begin // @[Csr.scala 46:26]
      mepc <= 64'h0; // @[Csr.scala 46:26]
    end else if (_T_73 & csr_rw) begin // @[RegMap.scala 46:34]
      if (3'h3 == io_uop_sys_code) begin // @[Mux.scala 80:57]
        mepc <= _T_42;
      end else if (3'h2 == io_uop_sys_code) begin // @[Mux.scala 80:57]
        mepc <= _T_40;
      end else begin
        mepc <= _T_44;
      end
    end else if (intr_0) begin // @[Csr.scala 101:15]
      mepc <= intr_mepc_0; // @[Csr.scala 103:10]
    end else if (io_uop_sys_code == 3'h4) begin // @[Csr.scala 75:40]
      mepc <= {{32'd0}, io_uop_pc}; // @[Csr.scala 76:10]
    end
    if (reset) begin // @[Csr.scala 47:26]
      mcause <= 64'h0; // @[Csr.scala 47:26]
    end else if (_T_97 & csr_rw) begin // @[RegMap.scala 46:34]
      if (3'h3 == io_uop_sys_code) begin // @[Mux.scala 80:57]
        mcause <= _T_42;
      end else if (3'h2 == io_uop_sys_code) begin // @[Mux.scala 80:57]
        mcause <= _T_40;
      end else begin
        mcause <= _T_44;
      end
    end else if (intr_0) begin // @[Csr.scala 101:15]
      mcause <= intr_mcause_0; // @[Csr.scala 104:12]
    end else if (io_uop_sys_code == 3'h4) begin // @[Csr.scala 75:40]
      mcause <= 64'hb; // @[Csr.scala 77:12]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mhartid = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mstatus = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mie = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mtvec = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mscratch = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mepc = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mcause = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_Fence(
  input         io_uop_valid,
  input  [31:0] io_uop_npc,
  input  [2:0]  io_uop_fu_code,
  input  [2:0]  io_uop_sys_code,
  output [31:0] io_ecp_jmp_pc,
  output        fence_i_0
);
  wire  fence_i = io_uop_valid & io_uop_fu_code == 3'h3 & io_uop_sys_code == 3'h7; // @[Fence.scala 16:62]
  assign io_ecp_jmp_pc = io_uop_npc; // @[Fence.scala 28:17]
  assign fence_i_0 = fence_i;
endmodule
module ysyx_210128_ExPipe0(
  input         clock,
  input         reset,
  input         io_uop_valid,
  input  [31:0] io_uop_pc,
  input  [31:0] io_uop_npc,
  input  [31:0] io_uop_inst,
  input  [2:0]  io_uop_fu_code,
  input  [3:0]  io_uop_alu_code,
  input  [3:0]  io_uop_jmp_code,
  input  [2:0]  io_uop_sys_code,
  input         io_uop_w_type,
  input  [31:0] io_uop_imm,
  input         io_uop_pred_br,
  input  [31:0] io_uop_pred_bpc,
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output        io_ecp_jmp_valid,
  output        io_ecp_jmp,
  output [31:0] io_ecp_jmp_pc,
  output        io_ecp_mis,
  output [63:0] io_ecp_rd_data,
  output        mtip,
  input  [63:0] intr_mcause,
  input  [63:0] instr_cnt,
  input  [63:0] intr_mstatus,
  output [29:0] _T_6_0,
  output        _T_5_0,
  input         intr,
  output        fence_i,
  input  [63:0] cycle_cnt,
  output [63:0] mstatus,
  input  [63:0] intr_mepc,
  input         mtip_0
);
  wire [31:0] alu_io_uop_pc; // @[Execution.scala 150:19]
  wire [31:0] alu_io_uop_npc; // @[Execution.scala 150:19]
  wire [2:0] alu_io_uop_fu_code; // @[Execution.scala 150:19]
  wire [3:0] alu_io_uop_alu_code; // @[Execution.scala 150:19]
  wire [3:0] alu_io_uop_jmp_code; // @[Execution.scala 150:19]
  wire  alu_io_uop_w_type; // @[Execution.scala 150:19]
  wire [31:0] alu_io_uop_imm; // @[Execution.scala 150:19]
  wire  alu_io_uop_pred_br; // @[Execution.scala 150:19]
  wire [31:0] alu_io_uop_pred_bpc; // @[Execution.scala 150:19]
  wire [63:0] alu_io_in1; // @[Execution.scala 150:19]
  wire [63:0] alu_io_in2; // @[Execution.scala 150:19]
  wire  alu_io_ecp_jmp_valid; // @[Execution.scala 150:19]
  wire  alu_io_ecp_jmp; // @[Execution.scala 150:19]
  wire [31:0] alu_io_ecp_jmp_pc; // @[Execution.scala 150:19]
  wire  alu_io_ecp_mis; // @[Execution.scala 150:19]
  wire [63:0] alu_io_ecp_rd_data; // @[Execution.scala 150:19]
  wire  csr_clock; // @[Execution.scala 154:19]
  wire  csr_reset; // @[Execution.scala 154:19]
  wire [31:0] csr_io_uop_pc; // @[Execution.scala 154:19]
  wire [31:0] csr_io_uop_inst; // @[Execution.scala 154:19]
  wire [2:0] csr_io_uop_sys_code; // @[Execution.scala 154:19]
  wire  csr_io_uop_pred_br; // @[Execution.scala 154:19]
  wire [31:0] csr_io_uop_pred_bpc; // @[Execution.scala 154:19]
  wire [63:0] csr_io_in1; // @[Execution.scala 154:19]
  wire  csr_io_ecp_jmp_valid; // @[Execution.scala 154:19]
  wire  csr_io_ecp_jmp; // @[Execution.scala 154:19]
  wire [31:0] csr_io_ecp_jmp_pc; // @[Execution.scala 154:19]
  wire  csr_io_ecp_mis; // @[Execution.scala 154:19]
  wire [63:0] csr_io_ecp_rd_data; // @[Execution.scala 154:19]
  wire  csr_mtip_0; // @[Execution.scala 154:19]
  wire [63:0] csr_intr_mcause_0; // @[Execution.scala 154:19]
  wire [63:0] csr_csr_minstret; // @[Execution.scala 154:19]
  wire [63:0] csr_intr_mstatus_0; // @[Execution.scala 154:19]
  wire [29:0] csr__T_6_0; // @[Execution.scala 154:19]
  wire  csr__T_5_0; // @[Execution.scala 154:19]
  wire  csr_intr_0; // @[Execution.scala 154:19]
  wire [63:0] csr_csr_mcycle; // @[Execution.scala 154:19]
  wire [63:0] csr_mstatus_0; // @[Execution.scala 154:19]
  wire [63:0] csr_intr_mepc_0; // @[Execution.scala 154:19]
  wire  csr_csr_mip_mtip; // @[Execution.scala 154:19]
  wire  fence_io_uop_valid; // @[Execution.scala 157:21]
  wire [31:0] fence_io_uop_npc; // @[Execution.scala 157:21]
  wire [2:0] fence_io_uop_fu_code; // @[Execution.scala 157:21]
  wire [2:0] fence_io_uop_sys_code; // @[Execution.scala 157:21]
  wire [31:0] fence_io_ecp_jmp_pc; // @[Execution.scala 157:21]
  wire  fence_fence_i_0; // @[Execution.scala 157:21]
  wire [31:0] _GEN_5 = io_uop_fu_code == 3'h3 & io_uop_sys_code != 3'h6 & io_uop_sys_code != 3'h7 ? io_uop_pred_bpc : 32'h0
    ; // @[Execution.scala 168:131 161:14 169:16]
  wire  _GEN_6 = io_uop_fu_code == 3'h3 & io_uop_sys_code != 3'h6 & io_uop_sys_code != 3'h7 & io_uop_pred_br; // @[Execution.scala 168:131 161:14 169:16]
  wire [2:0] _GEN_15 = io_uop_fu_code == 3'h3 & io_uop_sys_code != 3'h6 & io_uop_sys_code != 3'h7 ? io_uop_sys_code : 3'h0
    ; // @[Execution.scala 168:131 161:14 169:16]
  wire [31:0] _GEN_21 = io_uop_fu_code == 3'h3 & io_uop_sys_code != 3'h6 & io_uop_sys_code != 3'h7 ? io_uop_inst : 32'h0
    ; // @[Execution.scala 168:131 161:14 169:16]
  wire [31:0] _GEN_23 = io_uop_fu_code == 3'h3 & io_uop_sys_code != 3'h6 & io_uop_sys_code != 3'h7 ? io_uop_pc : 32'h0; // @[Execution.scala 168:131 161:14 169:16]
  wire [63:0] _GEN_25 = io_uop_fu_code == 3'h3 & io_uop_sys_code != 3'h6 & io_uop_sys_code != 3'h7 ? csr_io_ecp_rd_data
     : 64'h0; // @[Execution.scala 168:131 170:12 173:12]
  wire  _GEN_26 = io_uop_fu_code == 3'h3 & io_uop_sys_code != 3'h6 & io_uop_sys_code != 3'h7 ? csr_io_ecp_mis : 1'h1; // @[Execution.scala 168:131 170:12 173:12]
  wire [31:0] _GEN_27 = io_uop_fu_code == 3'h3 & io_uop_sys_code != 3'h6 & io_uop_sys_code != 3'h7 ? csr_io_ecp_jmp_pc
     : fence_io_ecp_jmp_pc; // @[Execution.scala 168:131 170:12 173:12]
  wire  _GEN_28 = io_uop_fu_code == 3'h3 & io_uop_sys_code != 3'h6 & io_uop_sys_code != 3'h7 ? csr_io_ecp_jmp : 1'h1; // @[Execution.scala 168:131 170:12 173:12]
  wire  _GEN_29 = io_uop_fu_code == 3'h3 & io_uop_sys_code != 3'h6 & io_uop_sys_code != 3'h7 ? csr_io_ecp_jmp_valid : 1'h1
    ; // @[Execution.scala 168:131 170:12 173:12]
  wire [2:0] _GEN_47 = io_uop_fu_code == 3'h3 & io_uop_sys_code != 3'h6 & io_uop_sys_code != 3'h7 ? 3'h0 :
    io_uop_sys_code; // @[Execution.scala 168:131 162:16 172:18]
  wire [2:0] _GEN_52 = io_uop_fu_code == 3'h3 & io_uop_sys_code != 3'h6 & io_uop_sys_code != 3'h7 ? 3'h0 :
    io_uop_fu_code; // @[Execution.scala 168:131 162:16 172:18]
  wire [31:0] _GEN_54 = io_uop_fu_code == 3'h3 & io_uop_sys_code != 3'h6 & io_uop_sys_code != 3'h7 ? 32'h0 : io_uop_npc; // @[Execution.scala 168:131 162:16 172:18]
  wire  _GEN_56 = io_uop_fu_code == 3'h3 & io_uop_sys_code != 3'h6 & io_uop_sys_code != 3'h7 ? 1'h0 : io_uop_valid; // @[Execution.scala 168:131 162:16 172:18]
  ysyx_210128_Alu alu ( // @[Execution.scala 150:19]
    .io_uop_pc(alu_io_uop_pc),
    .io_uop_npc(alu_io_uop_npc),
    .io_uop_fu_code(alu_io_uop_fu_code),
    .io_uop_alu_code(alu_io_uop_alu_code),
    .io_uop_jmp_code(alu_io_uop_jmp_code),
    .io_uop_w_type(alu_io_uop_w_type),
    .io_uop_imm(alu_io_uop_imm),
    .io_uop_pred_br(alu_io_uop_pred_br),
    .io_uop_pred_bpc(alu_io_uop_pred_bpc),
    .io_in1(alu_io_in1),
    .io_in2(alu_io_in2),
    .io_ecp_jmp_valid(alu_io_ecp_jmp_valid),
    .io_ecp_jmp(alu_io_ecp_jmp),
    .io_ecp_jmp_pc(alu_io_ecp_jmp_pc),
    .io_ecp_mis(alu_io_ecp_mis),
    .io_ecp_rd_data(alu_io_ecp_rd_data)
  );
  ysyx_210128_Csr csr ( // @[Execution.scala 154:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_uop_pc(csr_io_uop_pc),
    .io_uop_inst(csr_io_uop_inst),
    .io_uop_sys_code(csr_io_uop_sys_code),
    .io_uop_pred_br(csr_io_uop_pred_br),
    .io_uop_pred_bpc(csr_io_uop_pred_bpc),
    .io_in1(csr_io_in1),
    .io_ecp_jmp_valid(csr_io_ecp_jmp_valid),
    .io_ecp_jmp(csr_io_ecp_jmp),
    .io_ecp_jmp_pc(csr_io_ecp_jmp_pc),
    .io_ecp_mis(csr_io_ecp_mis),
    .io_ecp_rd_data(csr_io_ecp_rd_data),
    .mtip_0(csr_mtip_0),
    .intr_mcause_0(csr_intr_mcause_0),
    .csr_minstret(csr_csr_minstret),
    .intr_mstatus_0(csr_intr_mstatus_0),
    ._T_6_0(csr__T_6_0),
    ._T_5_0(csr__T_5_0),
    .intr_0(csr_intr_0),
    .csr_mcycle(csr_csr_mcycle),
    .mstatus_0(csr_mstatus_0),
    .intr_mepc_0(csr_intr_mepc_0),
    .csr_mip_mtip(csr_csr_mip_mtip)
  );
  ysyx_210128_Fence fence ( // @[Execution.scala 157:21]
    .io_uop_valid(fence_io_uop_valid),
    .io_uop_npc(fence_io_uop_npc),
    .io_uop_fu_code(fence_io_uop_fu_code),
    .io_uop_sys_code(fence_io_uop_sys_code),
    .io_ecp_jmp_pc(fence_io_ecp_jmp_pc),
    .fence_i_0(fence_fence_i_0)
  );
  assign io_ecp_jmp_valid = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? alu_io_ecp_jmp_valid : _GEN_29; // @[Execution.scala 165:79 167:12]
  assign io_ecp_jmp = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? alu_io_ecp_jmp : _GEN_28; // @[Execution.scala 165:79 167:12]
  assign io_ecp_jmp_pc = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? alu_io_ecp_jmp_pc : _GEN_27; // @[Execution.scala 165:79 167:12]
  assign io_ecp_mis = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? alu_io_ecp_mis : _GEN_26; // @[Execution.scala 165:79 167:12]
  assign io_ecp_rd_data = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? alu_io_ecp_rd_data : _GEN_25; // @[Execution.scala 165:79 167:12]
  assign mtip = csr_mtip_0;
  assign _T_6_0 = csr__T_6_0;
  assign _T_5_0 = csr__T_5_0;
  assign fence_i = fence_fence_i_0;
  assign mstatus = csr_mstatus_0;
  assign alu_io_uop_pc = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? io_uop_pc : 32'h0; // @[Execution.scala 160:14 165:79 166:16]
  assign alu_io_uop_npc = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? io_uop_npc : 32'h0; // @[Execution.scala 160:14 165:79 166:16]
  assign alu_io_uop_fu_code = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? io_uop_fu_code : 3'h0; // @[Execution.scala 160:14 165:79 166:16]
  assign alu_io_uop_alu_code = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? io_uop_alu_code : 4'h0; // @[Execution.scala 160:14 165:79 166:16]
  assign alu_io_uop_jmp_code = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? io_uop_jmp_code : 4'h0; // @[Execution.scala 160:14 165:79 166:16]
  assign alu_io_uop_w_type = (io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2) & io_uop_w_type; // @[Execution.scala 160:14 165:79 166:16]
  assign alu_io_uop_imm = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? io_uop_imm : 32'h0; // @[Execution.scala 160:14 165:79 166:16]
  assign alu_io_uop_pred_br = (io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2) & io_uop_pred_br; // @[Execution.scala 160:14 165:79 166:16]
  assign alu_io_uop_pred_bpc = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? io_uop_pred_bpc : 32'h0; // @[Execution.scala 160:14 165:79 166:16]
  assign alu_io_in1 = io_in1; // @[Execution.scala 151:14]
  assign alu_io_in2 = io_in2; // @[Execution.scala 152:14]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_uop_pc = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? 32'h0 : _GEN_23; // @[Execution.scala 161:14 165:79]
  assign csr_io_uop_inst = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? 32'h0 : _GEN_21; // @[Execution.scala 161:14 165:79]
  assign csr_io_uop_sys_code = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? 3'h0 : _GEN_15; // @[Execution.scala 161:14 165:79]
  assign csr_io_uop_pred_br = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? 1'h0 : _GEN_6; // @[Execution.scala 161:14 165:79]
  assign csr_io_uop_pred_bpc = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? 32'h0 : _GEN_5; // @[Execution.scala 161:14 165:79]
  assign csr_io_in1 = io_in1; // @[Execution.scala 155:14]
  assign csr_intr_mcause_0 = intr_mcause;
  assign csr_csr_minstret = instr_cnt;
  assign csr_intr_mstatus_0 = intr_mstatus;
  assign csr_intr_0 = intr;
  assign csr_csr_mcycle = cycle_cnt;
  assign csr_intr_mepc_0 = intr_mepc;
  assign csr_csr_mip_mtip = mtip_0;
  assign fence_io_uop_valid = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? 1'h0 : _GEN_56; // @[Execution.scala 162:16 165:79]
  assign fence_io_uop_npc = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? 32'h0 : _GEN_54; // @[Execution.scala 162:16 165:79]
  assign fence_io_uop_fu_code = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? 3'h0 : _GEN_52; // @[Execution.scala 162:16 165:79]
  assign fence_io_uop_sys_code = io_uop_fu_code == 3'h1 | io_uop_fu_code == 3'h2 ? 3'h0 : _GEN_47; // @[Execution.scala 162:16 165:79]
endmodule
module ysyx_210128_ExPipe1(
  input  [31:0] io_uop_pc,
  input  [31:0] io_uop_npc,
  input  [2:0]  io_uop_fu_code,
  input  [3:0]  io_uop_alu_code,
  input  [3:0]  io_uop_jmp_code,
  input         io_uop_w_type,
  input  [31:0] io_uop_imm,
  input         io_uop_pred_br,
  input  [31:0] io_uop_pred_bpc,
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output        io_ecp_jmp_valid,
  output        io_ecp_jmp,
  output [31:0] io_ecp_jmp_pc,
  output        io_ecp_mis,
  output [63:0] io_ecp_rd_data
);
  wire [31:0] alu_io_uop_pc; // @[Execution.scala 189:19]
  wire [31:0] alu_io_uop_npc; // @[Execution.scala 189:19]
  wire [2:0] alu_io_uop_fu_code; // @[Execution.scala 189:19]
  wire [3:0] alu_io_uop_alu_code; // @[Execution.scala 189:19]
  wire [3:0] alu_io_uop_jmp_code; // @[Execution.scala 189:19]
  wire  alu_io_uop_w_type; // @[Execution.scala 189:19]
  wire [31:0] alu_io_uop_imm; // @[Execution.scala 189:19]
  wire  alu_io_uop_pred_br; // @[Execution.scala 189:19]
  wire [31:0] alu_io_uop_pred_bpc; // @[Execution.scala 189:19]
  wire [63:0] alu_io_in1; // @[Execution.scala 189:19]
  wire [63:0] alu_io_in2; // @[Execution.scala 189:19]
  wire  alu_io_ecp_jmp_valid; // @[Execution.scala 189:19]
  wire  alu_io_ecp_jmp; // @[Execution.scala 189:19]
  wire [31:0] alu_io_ecp_jmp_pc; // @[Execution.scala 189:19]
  wire  alu_io_ecp_mis; // @[Execution.scala 189:19]
  wire [63:0] alu_io_ecp_rd_data; // @[Execution.scala 189:19]
  ysyx_210128_Alu alu ( // @[Execution.scala 189:19]
    .io_uop_pc(alu_io_uop_pc),
    .io_uop_npc(alu_io_uop_npc),
    .io_uop_fu_code(alu_io_uop_fu_code),
    .io_uop_alu_code(alu_io_uop_alu_code),
    .io_uop_jmp_code(alu_io_uop_jmp_code),
    .io_uop_w_type(alu_io_uop_w_type),
    .io_uop_imm(alu_io_uop_imm),
    .io_uop_pred_br(alu_io_uop_pred_br),
    .io_uop_pred_bpc(alu_io_uop_pred_bpc),
    .io_in1(alu_io_in1),
    .io_in2(alu_io_in2),
    .io_ecp_jmp_valid(alu_io_ecp_jmp_valid),
    .io_ecp_jmp(alu_io_ecp_jmp),
    .io_ecp_jmp_pc(alu_io_ecp_jmp_pc),
    .io_ecp_mis(alu_io_ecp_mis),
    .io_ecp_rd_data(alu_io_ecp_rd_data)
  );
  assign io_ecp_jmp_valid = alu_io_ecp_jmp_valid; // @[Execution.scala 194:10]
  assign io_ecp_jmp = alu_io_ecp_jmp; // @[Execution.scala 194:10]
  assign io_ecp_jmp_pc = alu_io_ecp_jmp_pc; // @[Execution.scala 194:10]
  assign io_ecp_mis = alu_io_ecp_mis; // @[Execution.scala 194:10]
  assign io_ecp_rd_data = alu_io_ecp_rd_data; // @[Execution.scala 194:10]
  assign alu_io_uop_pc = io_uop_pc; // @[Execution.scala 190:14]
  assign alu_io_uop_npc = io_uop_npc; // @[Execution.scala 190:14]
  assign alu_io_uop_fu_code = io_uop_fu_code; // @[Execution.scala 190:14]
  assign alu_io_uop_alu_code = io_uop_alu_code; // @[Execution.scala 190:14]
  assign alu_io_uop_jmp_code = io_uop_jmp_code; // @[Execution.scala 190:14]
  assign alu_io_uop_w_type = io_uop_w_type; // @[Execution.scala 190:14]
  assign alu_io_uop_imm = io_uop_imm; // @[Execution.scala 190:14]
  assign alu_io_uop_pred_br = io_uop_pred_br; // @[Execution.scala 190:14]
  assign alu_io_uop_pred_bpc = io_uop_pred_bpc; // @[Execution.scala 190:14]
  assign alu_io_in1 = io_in1; // @[Execution.scala 191:14]
  assign alu_io_in2 = io_in2; // @[Execution.scala 192:14]
endmodule
module ysyx_210128_Lsu(
  input         clock,
  input         reset,
  input         io_uop_valid,
  input  [2:0]  io_uop_fu_code,
  input  [1:0]  io_uop_mem_code,
  input  [1:0]  io_uop_mem_size,
  input  [31:0] io_uop_imm,
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output        io_ecp_store_valid,
  output [63:0] io_ecp_rd_data,
  output        io_busy,
  input         io_dmem_st_req_ready,
  output        io_dmem_st_req_valid,
  output [31:0] io_dmem_st_req_bits_addr,
  output [63:0] io_dmem_st_req_bits_wdata,
  output [7:0]  io_dmem_st_req_bits_wmask,
  output [1:0]  io_dmem_st_req_bits_size,
  output        io_dmem_st_resp_ready,
  input         io_dmem_st_resp_valid,
  input         io_dmem_ld_req_ready,
  output        io_dmem_ld_req_valid,
  output [31:0] io_dmem_ld_req_bits_addr,
  output [1:0]  io_dmem_ld_req_bits_size,
  output        io_dmem_ld_resp_ready,
  input         io_dmem_ld_resp_valid,
  input  [63:0] io_dmem_ld_resp_bits_rdata,
  input         io_flush,
  output        io_wakeup
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  _T_valid = io_flush ? 1'h0 : io_uop_valid; // @[Utils.scala 68:20]
  wire [2:0] _T_fu_code = io_flush ? 3'h0 : io_uop_fu_code; // @[Utils.scala 68:20]
  wire [1:0] _T_mem_code = io_flush ? 2'h0 : io_uop_mem_code; // @[Utils.scala 68:20]
  wire [1:0] _T_mem_size = io_flush ? 2'h0 : io_uop_mem_size; // @[Utils.scala 68:20]
  wire [31:0] _T_imm = io_flush ? 32'h0 : io_uop_imm; // @[Utils.scala 68:20]
  wire  _T_2 = io_uop_valid | io_flush; // @[Utils.scala 69:72]
  reg  r_valid; // @[Reg.scala 27:20]
  reg [2:0] r_fu_code; // @[Reg.scala 27:20]
  reg [1:0] r_mem_code; // @[Reg.scala 27:20]
  reg [1:0] r_mem_size; // @[Reg.scala 27:20]
  reg [31:0] r_imm; // @[Reg.scala 27:20]
  wire  uop_valid = io_uop_valid ? _T_valid : r_valid; // @[Utils.scala 69:8]
  wire [2:0] uop_fu_code = io_uop_valid ? _T_fu_code : r_fu_code; // @[Utils.scala 69:8]
  wire [1:0] uop_mem_code = io_uop_valid ? _T_mem_code : r_mem_code; // @[Utils.scala 69:8]
  wire [1:0] uop_mem_size = io_uop_valid ? _T_mem_size : r_mem_size; // @[Utils.scala 69:8]
  wire [31:0] uop_imm = io_uop_valid ? _T_imm : r_imm; // @[Utils.scala 69:8]
  wire [63:0] _T_3 = io_flush ? 64'h0 : io_in1; // @[Utils.scala 68:20]
  reg [63:0] r_1; // @[Reg.scala 27:20]
  wire [63:0] in1 = io_uop_valid ? _T_3 : r_1; // @[Utils.scala 69:8]
  wire [63:0] _T_6 = io_flush ? 64'h0 : io_in2; // @[Utils.scala 68:20]
  reg [63:0] r_2; // @[Reg.scala 27:20]
  wire [63:0] in2 = io_uop_valid ? _T_6 : r_2; // @[Utils.scala 69:8]
  reg  completed; // @[Lsu.scala 27:26]
  wire  _GEN_27 = io_uop_valid ? 1'h0 : completed; // @[Lsu.scala 28:21 29:15 27:26]
  wire  is_mem = uop_fu_code == 3'h4; // @[Lsu.scala 32:29]
  wire  _T_9 = uop_mem_code == 2'h1; // @[Lsu.scala 33:31]
  wire  _T_10 = uop_mem_code == 2'h2; // @[Lsu.scala 33:65]
  wire  is_load = uop_mem_code == 2'h1 | uop_mem_code == 2'h2; // @[Lsu.scala 33:49]
  wire  is_store = uop_mem_code == 2'h3; // @[Lsu.scala 34:32]
  reg [1:0] state; // @[Lsu.scala 37:22]
  wire [31:0] addr = in1[31:0] + uop_imm; // @[Lsu.scala 44:26]
  wire [2:0] addr_offset = addr[2:0]; // @[Lsu.scala 45:25]
  wire  mmio = ~addr[31]; // @[Lsu.scala 48:24]
  wire [14:0] _T_15 = 15'hff << addr_offset; // @[Lsu.scala 50:29]
  wire [7:0] mask = _T_15[7:0]; // @[Lsu.scala 50:44]
  wire [7:0] _T_17 = 2'h1 == uop_mem_size ? 8'h3 : 8'h1; // @[Mux.scala 80:57]
  wire [7:0] _T_19 = 2'h2 == uop_mem_size ? 8'hf : _T_17; // @[Mux.scala 80:57]
  wire [7:0] wmask = 2'h3 == uop_mem_size ? 8'hff : _T_19; // @[Mux.scala 80:57]
  wire  _T_22 = addr_offset == 3'h7; // @[Lsu.scala 64:40]
  wire  _T_23 = addr_offset > 3'h4; // @[Lsu.scala 65:49]
  wire  _T_24 = addr_offset != 3'h0; // @[Lsu.scala 66:40]
  wire  _T_28 = 2'h2 == uop_mem_size ? _T_23 : 2'h1 == uop_mem_size & _T_22; // @[Mux.scala 80:57]
  wire  _T_30 = 2'h3 == uop_mem_size ? _T_24 : _T_28; // @[Mux.scala 80:57]
  wire  addr_unaligned = is_mem & _T_30; // @[Lsu.scala 62:27]
  wire [31:0] _T_33 = {addr[31:3],3'h0}; // @[Cat.scala 30:58]
  wire [5:0] _T_35 = {addr_offset, 3'h0}; // @[Lsu.scala 72:47]
  wire [126:0] _GEN_0 = {{63'd0}, in2}; // @[Lsu.scala 72:31]
  wire [126:0] _T_36 = _GEN_0 << _T_35; // @[Lsu.scala 72:31]
  wire [14:0] _GEN_1 = {{7'd0}, wmask}; // @[Lsu.scala 73:39]
  wire [14:0] _T_38 = _GEN_1 << addr_offset; // @[Lsu.scala 73:39]
  wire  _T_45 = uop_valid & state == 2'h0 & ~addr_unaligned; // @[Lsu.scala 77:56]
  wire  _T_46 = uop_valid & state == 2'h0 & ~addr_unaligned & is_store; // @[Lsu.scala 77:75]
  wire  _T_48 = io_uop_valid | ~completed; // @[Lsu.scala 78:48]
  wire  _T_59 = _T_45 & is_load; // @[Lsu.scala 88:75]
  reg  store_valid; // @[Lsu.scala 94:28]
  wire  _T_64 = io_dmem_ld_req_ready & io_dmem_ld_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_65 = io_dmem_st_req_ready & io_dmem_st_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_28 = _T_65 ? 2'h2 : state; // @[Lsu.scala 103:35 104:15 37:22]
  wire  _GEN_29 = _T_65 | store_valid; // @[Lsu.scala 103:35 105:21 94:28]
  wire  _GEN_32 = addr_unaligned | _GEN_27; // @[Lsu.scala 107:29 108:19]
  wire  _T_67 = io_dmem_ld_resp_ready & io_dmem_ld_resp_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _T_69 = io_dmem_ld_resp_bits_rdata >> _T_35; // @[Lsu.scala 113:41]
  wire [63:0] _GEN_33 = _T_67 ? _T_69 : 64'h0; // @[Lsu.scala 112:29 113:19]
  wire  _GEN_35 = _T_67 | _GEN_27; // @[Lsu.scala 112:29 119:19]
  wire [1:0] _GEN_36 = _T_67 ? 2'h0 : state; // @[Lsu.scala 112:29 120:15 37:22]
  wire  _T_71 = io_dmem_st_resp_ready & io_dmem_st_resp_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_37 = _T_71 | _GEN_27; // @[Lsu.scala 124:29 129:19]
  wire [1:0] _GEN_38 = _T_71 ? 2'h0 : state; // @[Lsu.scala 124:29 130:15 37:22]
  wire  _GEN_39 = 2'h2 == state ? _GEN_37 : _GEN_27; // @[Lsu.scala 98:18]
  wire [1:0] _GEN_40 = 2'h2 == state ? _GEN_38 : state; // @[Lsu.scala 98:18 37:22]
  wire [63:0] _GEN_41 = 2'h1 == state ? _GEN_33 : 64'h0; // @[Lsu.scala 98:18]
  wire  _GEN_43 = 2'h1 == state ? _GEN_35 : _GEN_39; // @[Lsu.scala 98:18]
  wire  _GEN_47 = 2'h0 == state ? _GEN_32 : _GEN_43; // @[Lsu.scala 98:18]
  wire [63:0] load_data = 2'h0 == state ? 64'h0 : _GEN_41; // @[Lsu.scala 98:18]
  wire  _GEN_50 = io_flush | _GEN_47; // @[Lsu.scala 136:19 137:15]
  wire [55:0] _T_75 = load_data[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_77 = {_T_75,load_data[7:0]}; // @[Cat.scala 30:58]
  wire [47:0] _T_80 = load_data[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_82 = {_T_80,load_data[15:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_85 = load_data[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_87 = {_T_85,load_data[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_89 = 2'h1 == uop_mem_size ? _T_82 : _T_77; // @[Mux.scala 80:57]
  wire [63:0] _T_91 = 2'h2 == uop_mem_size ? _T_87 : _T_89; // @[Mux.scala 80:57]
  wire [63:0] _T_93 = 2'h3 == uop_mem_size ? load_data : _T_91; // @[Mux.scala 80:57]
  wire [63:0] ld_out = _T_9 ? _T_93 : 64'h0; // @[Lsu.scala 145:16]
  wire [63:0] _T_98 = {56'h0,load_data[7:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_101 = {48'h0,load_data[15:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_104 = {32'h0,load_data[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_106 = 2'h1 == uop_mem_size ? _T_101 : _T_98; // @[Mux.scala 80:57]
  wire [63:0] _T_108 = 2'h2 == uop_mem_size ? _T_104 : _T_106; // @[Mux.scala 80:57]
  wire [63:0] _T_110 = 2'h3 == uop_mem_size ? load_data : _T_108; // @[Mux.scala 80:57]
  wire [63:0] ldu_out = _T_10 ? _T_110 : 64'h0; // @[Lsu.scala 152:17]
  wire [63:0] _T_113 = 2'h1 == uop_mem_code ? ld_out : 64'h0; // @[Mux.scala 80:57]
  assign io_ecp_store_valid = store_valid; // @[Lsu.scala 165:22]
  assign io_ecp_rd_data = 2'h2 == uop_mem_code ? ldu_out : _T_113; // @[Mux.scala 80:57]
  assign io_busy = io_dmem_ld_req_valid | io_dmem_st_req_valid | state == 2'h1 & ~_T_67 | state == 2'h2 & ~_T_71; // @[Lsu.scala 168:86]
  assign io_dmem_st_req_valid = _T_46 & (io_uop_valid | ~completed); // @[Lsu.scala 78:33]
  assign io_dmem_st_req_bits_addr = mmio ? addr : _T_33; // @[Lsu.scala 71:27]
  assign io_dmem_st_req_bits_wdata = _T_36[63:0]; // @[Lsu.scala 72:53]
  assign io_dmem_st_req_bits_wmask = mask & _T_38[7:0]; // @[Lsu.scala 73:29]
  assign io_dmem_st_req_bits_size = mmio ? uop_mem_size : 2'h3; // @[Lsu.scala 75:27]
  assign io_dmem_st_resp_ready = io_dmem_st_resp_valid; // @[Lsu.scala 80:21]
  assign io_dmem_ld_req_valid = _T_59 & _T_48; // @[Lsu.scala 89:32]
  assign io_dmem_ld_req_bits_addr = mmio ? addr : _T_33; // @[Lsu.scala 82:27]
  assign io_dmem_ld_req_bits_size = mmio ? uop_mem_size : 2'h3; // @[Lsu.scala 86:27]
  assign io_dmem_ld_resp_ready = io_dmem_ld_resp_valid; // @[Lsu.scala 91:21]
  assign io_wakeup = 2'h0 == state ? 1'h0 : 2'h1 == state & _T_67; // @[Lsu.scala 96:13 98:18]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 27:20]
      r_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      if (io_flush) begin // @[Utils.scala 68:20]
        r_valid <= 1'h0;
      end else begin
        r_valid <= io_uop_valid;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_fu_code <= 3'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      if (io_flush) begin // @[Utils.scala 68:20]
        r_fu_code <= 3'h0;
      end else begin
        r_fu_code <= io_uop_fu_code;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_mem_code <= 2'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      if (io_flush) begin // @[Utils.scala 68:20]
        r_mem_code <= 2'h0;
      end else begin
        r_mem_code <= io_uop_mem_code;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_mem_size <= 2'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      if (io_flush) begin // @[Utils.scala 68:20]
        r_mem_size <= 2'h0;
      end else begin
        r_mem_size <= io_uop_mem_size;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_imm <= 32'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      if (io_flush) begin // @[Utils.scala 68:20]
        r_imm <= 32'h0;
      end else begin
        r_imm <= io_uop_imm;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1 <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      if (io_flush) begin // @[Utils.scala 68:20]
        r_1 <= 64'h0;
      end else begin
        r_1 <= io_in1;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_2 <= 64'h0; // @[Reg.scala 27:20]
    end else if (_T_2) begin // @[Reg.scala 28:19]
      if (io_flush) begin // @[Utils.scala 68:20]
        r_2 <= 64'h0;
      end else begin
        r_2 <= io_in2;
      end
    end
    completed <= reset | _GEN_50; // @[Lsu.scala 27:{26,26}]
    if (reset) begin // @[Lsu.scala 37:22]
      state <= 2'h0; // @[Lsu.scala 37:22]
    end else if (io_flush) begin // @[Lsu.scala 136:19]
      state <= 2'h0; // @[Lsu.scala 138:11]
    end else if (2'h0 == state) begin // @[Lsu.scala 98:18]
      if (_T_64) begin // @[Lsu.scala 100:28]
        state <= 2'h1; // @[Lsu.scala 101:15]
      end else begin
        state <= _GEN_28;
      end
    end else if (2'h1 == state) begin // @[Lsu.scala 98:18]
      state <= _GEN_36;
    end else begin
      state <= _GEN_40;
    end
    if (reset) begin // @[Lsu.scala 94:28]
      store_valid <= 1'h0; // @[Lsu.scala 94:28]
    end else if (2'h0 == state) begin // @[Lsu.scala 98:18]
      if (_T_64) begin // @[Lsu.scala 100:28]
        store_valid <= 1'h0; // @[Lsu.scala 102:21]
      end else begin
        store_valid <= _GEN_29;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_fu_code = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  r_mem_code = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  r_mem_size = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  r_imm = _RAND_4[31:0];
  _RAND_5 = {2{`RANDOM}};
  r_1 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  r_2 = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  completed = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  store_valid = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_ExPipe2(
  input         clock,
  input         reset,
  input         io_uop_valid,
  input  [2:0]  io_uop_fu_code,
  input  [1:0]  io_uop_mem_code,
  input  [1:0]  io_uop_mem_size,
  input  [31:0] io_uop_imm,
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output        io_ecp_store_valid,
  output [63:0] io_ecp_rd_data,
  output        io_ready,
  input         io_dmem_st_req_ready,
  output        io_dmem_st_req_valid,
  output [31:0] io_dmem_st_req_bits_addr,
  output [63:0] io_dmem_st_req_bits_wdata,
  output [7:0]  io_dmem_st_req_bits_wmask,
  output [1:0]  io_dmem_st_req_bits_size,
  output        io_dmem_st_resp_ready,
  input         io_dmem_st_resp_valid,
  input         io_dmem_ld_req_ready,
  output        io_dmem_ld_req_valid,
  output [31:0] io_dmem_ld_req_bits_addr,
  output [1:0]  io_dmem_ld_req_bits_size,
  output        io_dmem_ld_resp_ready,
  input         io_dmem_ld_resp_valid,
  input  [63:0] io_dmem_ld_resp_bits_rdata,
  input         io_flush,
  output        io_wakeup
);
  wire  lsu_clock; // @[Execution.scala 217:19]
  wire  lsu_reset; // @[Execution.scala 217:19]
  wire  lsu_io_uop_valid; // @[Execution.scala 217:19]
  wire [2:0] lsu_io_uop_fu_code; // @[Execution.scala 217:19]
  wire [1:0] lsu_io_uop_mem_code; // @[Execution.scala 217:19]
  wire [1:0] lsu_io_uop_mem_size; // @[Execution.scala 217:19]
  wire [31:0] lsu_io_uop_imm; // @[Execution.scala 217:19]
  wire [63:0] lsu_io_in1; // @[Execution.scala 217:19]
  wire [63:0] lsu_io_in2; // @[Execution.scala 217:19]
  wire  lsu_io_ecp_store_valid; // @[Execution.scala 217:19]
  wire [63:0] lsu_io_ecp_rd_data; // @[Execution.scala 217:19]
  wire  lsu_io_busy; // @[Execution.scala 217:19]
  wire  lsu_io_dmem_st_req_ready; // @[Execution.scala 217:19]
  wire  lsu_io_dmem_st_req_valid; // @[Execution.scala 217:19]
  wire [31:0] lsu_io_dmem_st_req_bits_addr; // @[Execution.scala 217:19]
  wire [63:0] lsu_io_dmem_st_req_bits_wdata; // @[Execution.scala 217:19]
  wire [7:0] lsu_io_dmem_st_req_bits_wmask; // @[Execution.scala 217:19]
  wire [1:0] lsu_io_dmem_st_req_bits_size; // @[Execution.scala 217:19]
  wire  lsu_io_dmem_st_resp_ready; // @[Execution.scala 217:19]
  wire  lsu_io_dmem_st_resp_valid; // @[Execution.scala 217:19]
  wire  lsu_io_dmem_ld_req_ready; // @[Execution.scala 217:19]
  wire  lsu_io_dmem_ld_req_valid; // @[Execution.scala 217:19]
  wire [31:0] lsu_io_dmem_ld_req_bits_addr; // @[Execution.scala 217:19]
  wire [1:0] lsu_io_dmem_ld_req_bits_size; // @[Execution.scala 217:19]
  wire  lsu_io_dmem_ld_resp_ready; // @[Execution.scala 217:19]
  wire  lsu_io_dmem_ld_resp_valid; // @[Execution.scala 217:19]
  wire [63:0] lsu_io_dmem_ld_resp_bits_rdata; // @[Execution.scala 217:19]
  wire  lsu_io_flush; // @[Execution.scala 217:19]
  wire  lsu_io_wakeup; // @[Execution.scala 217:19]
  ysyx_210128_Lsu lsu ( // @[Execution.scala 217:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io_uop_valid(lsu_io_uop_valid),
    .io_uop_fu_code(lsu_io_uop_fu_code),
    .io_uop_mem_code(lsu_io_uop_mem_code),
    .io_uop_mem_size(lsu_io_uop_mem_size),
    .io_uop_imm(lsu_io_uop_imm),
    .io_in1(lsu_io_in1),
    .io_in2(lsu_io_in2),
    .io_ecp_store_valid(lsu_io_ecp_store_valid),
    .io_ecp_rd_data(lsu_io_ecp_rd_data),
    .io_busy(lsu_io_busy),
    .io_dmem_st_req_ready(lsu_io_dmem_st_req_ready),
    .io_dmem_st_req_valid(lsu_io_dmem_st_req_valid),
    .io_dmem_st_req_bits_addr(lsu_io_dmem_st_req_bits_addr),
    .io_dmem_st_req_bits_wdata(lsu_io_dmem_st_req_bits_wdata),
    .io_dmem_st_req_bits_wmask(lsu_io_dmem_st_req_bits_wmask),
    .io_dmem_st_req_bits_size(lsu_io_dmem_st_req_bits_size),
    .io_dmem_st_resp_ready(lsu_io_dmem_st_resp_ready),
    .io_dmem_st_resp_valid(lsu_io_dmem_st_resp_valid),
    .io_dmem_ld_req_ready(lsu_io_dmem_ld_req_ready),
    .io_dmem_ld_req_valid(lsu_io_dmem_ld_req_valid),
    .io_dmem_ld_req_bits_addr(lsu_io_dmem_ld_req_bits_addr),
    .io_dmem_ld_req_bits_size(lsu_io_dmem_ld_req_bits_size),
    .io_dmem_ld_resp_ready(lsu_io_dmem_ld_resp_ready),
    .io_dmem_ld_resp_valid(lsu_io_dmem_ld_resp_valid),
    .io_dmem_ld_resp_bits_rdata(lsu_io_dmem_ld_resp_bits_rdata),
    .io_flush(lsu_io_flush),
    .io_wakeup(lsu_io_wakeup)
  );
  assign io_ecp_store_valid = lsu_io_ecp_store_valid; // @[Execution.scala 225:10]
  assign io_ecp_rd_data = lsu_io_ecp_rd_data; // @[Execution.scala 225:10]
  assign io_ready = ~lsu_io_busy; // @[Execution.scala 226:15]
  assign io_dmem_st_req_valid = lsu_io_dmem_st_req_valid; // @[Execution.scala 221:18]
  assign io_dmem_st_req_bits_addr = lsu_io_dmem_st_req_bits_addr; // @[Execution.scala 221:18]
  assign io_dmem_st_req_bits_wdata = lsu_io_dmem_st_req_bits_wdata; // @[Execution.scala 221:18]
  assign io_dmem_st_req_bits_wmask = lsu_io_dmem_st_req_bits_wmask; // @[Execution.scala 221:18]
  assign io_dmem_st_req_bits_size = lsu_io_dmem_st_req_bits_size; // @[Execution.scala 221:18]
  assign io_dmem_st_resp_ready = lsu_io_dmem_st_resp_ready; // @[Execution.scala 221:18]
  assign io_dmem_ld_req_valid = lsu_io_dmem_ld_req_valid; // @[Execution.scala 222:18]
  assign io_dmem_ld_req_bits_addr = lsu_io_dmem_ld_req_bits_addr; // @[Execution.scala 222:18]
  assign io_dmem_ld_req_bits_size = lsu_io_dmem_ld_req_bits_size; // @[Execution.scala 222:18]
  assign io_dmem_ld_resp_ready = lsu_io_dmem_ld_resp_ready; // @[Execution.scala 222:18]
  assign io_wakeup = lsu_io_wakeup; // @[Execution.scala 227:13]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io_uop_valid = io_uop_valid; // @[Execution.scala 218:14]
  assign lsu_io_uop_fu_code = io_uop_fu_code; // @[Execution.scala 218:14]
  assign lsu_io_uop_mem_code = io_uop_mem_code; // @[Execution.scala 218:14]
  assign lsu_io_uop_mem_size = io_uop_mem_size; // @[Execution.scala 218:14]
  assign lsu_io_uop_imm = io_uop_imm; // @[Execution.scala 218:14]
  assign lsu_io_in1 = io_in1; // @[Execution.scala 219:14]
  assign lsu_io_in2 = io_in2; // @[Execution.scala 220:14]
  assign lsu_io_dmem_st_req_ready = io_dmem_st_req_ready; // @[Execution.scala 221:18]
  assign lsu_io_dmem_st_resp_valid = io_dmem_st_resp_valid; // @[Execution.scala 221:18]
  assign lsu_io_dmem_ld_req_ready = io_dmem_ld_req_ready; // @[Execution.scala 222:18]
  assign lsu_io_dmem_ld_resp_valid = io_dmem_ld_resp_valid; // @[Execution.scala 222:18]
  assign lsu_io_dmem_ld_resp_bits_rdata = io_dmem_ld_resp_bits_rdata; // @[Execution.scala 222:18]
  assign lsu_io_flush = io_flush; // @[Execution.scala 223:16]
endmodule
module ysyx_210128_Execution(
  input         clock,
  input         reset,
  input         io_in_0_valid,
  input  [31:0] io_in_0_pc,
  input  [31:0] io_in_0_npc,
  input  [31:0] io_in_0_inst,
  input  [2:0]  io_in_0_fu_code,
  input  [3:0]  io_in_0_alu_code,
  input  [3:0]  io_in_0_jmp_code,
  input  [2:0]  io_in_0_sys_code,
  input         io_in_0_w_type,
  input  [1:0]  io_in_0_rs1_src,
  input  [1:0]  io_in_0_rs2_src,
  input         io_in_0_rd_en,
  input  [31:0] io_in_0_imm,
  input         io_in_0_pred_br,
  input  [31:0] io_in_0_pred_bpc,
  input  [5:0]  io_in_0_rd_paddr,
  input  [3:0]  io_in_0_rob_addr,
  input         io_in_1_valid,
  input  [31:0] io_in_1_pc,
  input  [31:0] io_in_1_npc,
  input  [2:0]  io_in_1_fu_code,
  input  [3:0]  io_in_1_alu_code,
  input  [3:0]  io_in_1_jmp_code,
  input         io_in_1_w_type,
  input  [1:0]  io_in_1_rs1_src,
  input  [1:0]  io_in_1_rs2_src,
  input         io_in_1_rd_en,
  input  [31:0] io_in_1_imm,
  input         io_in_1_pred_br,
  input  [31:0] io_in_1_pred_bpc,
  input  [5:0]  io_in_1_rd_paddr,
  input  [3:0]  io_in_1_rob_addr,
  input         io_in_2_valid,
  input  [31:0] io_in_2_pc,
  input  [2:0]  io_in_2_fu_code,
  input  [3:0]  io_in_2_alu_code,
  input  [1:0]  io_in_2_mem_code,
  input  [1:0]  io_in_2_mem_size,
  input         io_in_2_w_type,
  input  [1:0]  io_in_2_rs1_src,
  input  [1:0]  io_in_2_rs2_src,
  input         io_in_2_rd_en,
  input  [31:0] io_in_2_imm,
  input  [5:0]  io_in_2_rd_paddr,
  input  [3:0]  io_in_2_rob_addr,
  input  [63:0] io_rs1_data_0,
  input  [63:0] io_rs1_data_1,
  input  [63:0] io_rs1_data_2,
  input  [63:0] io_rs2_data_0,
  input  [63:0] io_rs2_data_1,
  input  [63:0] io_rs2_data_2,
  output        io_out_0_valid,
  output [3:0]  io_out_0_rob_addr,
  output        io_out_1_valid,
  output [3:0]  io_out_1_rob_addr,
  output        io_out_2_valid,
  output [3:0]  io_out_2_rob_addr,
  output        io_out_ecp_0_jmp_valid,
  output        io_out_ecp_0_jmp,
  output [31:0] io_out_ecp_0_jmp_pc,
  output        io_out_ecp_0_mis,
  output        io_out_ecp_1_jmp_valid,
  output        io_out_ecp_1_jmp,
  output [31:0] io_out_ecp_1_jmp_pc,
  output        io_out_ecp_1_mis,
  output        io_out_ecp_2_store_valid,
  output        io_rd_en_0,
  output        io_rd_en_1,
  output        io_rd_en_2,
  output [5:0]  io_rd_paddr_0,
  output [5:0]  io_rd_paddr_1,
  output [5:0]  io_rd_paddr_2,
  output [63:0] io_rd_data_0,
  output [63:0] io_rd_data_1,
  output [63:0] io_rd_data_2,
  input         io_flush,
  output        io_lsu_ready,
  input         io_dmem_st_req_ready,
  output        io_dmem_st_req_valid,
  output [31:0] io_dmem_st_req_bits_addr,
  output [63:0] io_dmem_st_req_bits_wdata,
  output [7:0]  io_dmem_st_req_bits_wmask,
  output [1:0]  io_dmem_st_req_bits_size,
  output        io_dmem_st_resp_ready,
  input         io_dmem_st_resp_valid,
  input         io_dmem_ld_req_ready,
  output        io_dmem_ld_req_valid,
  output [31:0] io_dmem_ld_req_bits_addr,
  output [1:0]  io_dmem_ld_req_bits_size,
  output        io_dmem_ld_resp_ready,
  input         io_dmem_ld_resp_valid,
  input  [63:0] io_dmem_ld_resp_bits_rdata,
  output        io_lsu_wakeup_uop_valid,
  output        io_lsu_wakeup_uop_rd_en,
  output [5:0]  io_lsu_wakeup_uop_rd_paddr,
  output        mtip,
  input  [63:0] intr_mcause,
  input  [63:0] instr_cnt,
  input  [63:0] intr_mstatus,
  output [29:0] _T_6_0,
  output        _T_5_0,
  input         intr,
  output        fence_i,
  input  [63:0] cycle_cnt,
  output [63:0] mstatus,
  input  [63:0] intr_mepc,
  input         mtip_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  wire  pipe0_clock; // @[Execution.scala 65:21]
  wire  pipe0_reset; // @[Execution.scala 65:21]
  wire  pipe0_io_uop_valid; // @[Execution.scala 65:21]
  wire [31:0] pipe0_io_uop_pc; // @[Execution.scala 65:21]
  wire [31:0] pipe0_io_uop_npc; // @[Execution.scala 65:21]
  wire [31:0] pipe0_io_uop_inst; // @[Execution.scala 65:21]
  wire [2:0] pipe0_io_uop_fu_code; // @[Execution.scala 65:21]
  wire [3:0] pipe0_io_uop_alu_code; // @[Execution.scala 65:21]
  wire [3:0] pipe0_io_uop_jmp_code; // @[Execution.scala 65:21]
  wire [2:0] pipe0_io_uop_sys_code; // @[Execution.scala 65:21]
  wire  pipe0_io_uop_w_type; // @[Execution.scala 65:21]
  wire [31:0] pipe0_io_uop_imm; // @[Execution.scala 65:21]
  wire  pipe0_io_uop_pred_br; // @[Execution.scala 65:21]
  wire [31:0] pipe0_io_uop_pred_bpc; // @[Execution.scala 65:21]
  wire [63:0] pipe0_io_in1; // @[Execution.scala 65:21]
  wire [63:0] pipe0_io_in2; // @[Execution.scala 65:21]
  wire  pipe0_io_ecp_jmp_valid; // @[Execution.scala 65:21]
  wire  pipe0_io_ecp_jmp; // @[Execution.scala 65:21]
  wire [31:0] pipe0_io_ecp_jmp_pc; // @[Execution.scala 65:21]
  wire  pipe0_io_ecp_mis; // @[Execution.scala 65:21]
  wire [63:0] pipe0_io_ecp_rd_data; // @[Execution.scala 65:21]
  wire  pipe0_mtip; // @[Execution.scala 65:21]
  wire [63:0] pipe0_intr_mcause; // @[Execution.scala 65:21]
  wire [63:0] pipe0_instr_cnt; // @[Execution.scala 65:21]
  wire [63:0] pipe0_intr_mstatus; // @[Execution.scala 65:21]
  wire [29:0] pipe0__T_6_0; // @[Execution.scala 65:21]
  wire  pipe0__T_5_0; // @[Execution.scala 65:21]
  wire  pipe0_intr; // @[Execution.scala 65:21]
  wire  pipe0_fence_i; // @[Execution.scala 65:21]
  wire [63:0] pipe0_cycle_cnt; // @[Execution.scala 65:21]
  wire [63:0] pipe0_mstatus; // @[Execution.scala 65:21]
  wire [63:0] pipe0_intr_mepc; // @[Execution.scala 65:21]
  wire  pipe0_mtip_0; // @[Execution.scala 65:21]
  wire [31:0] pipe1_io_uop_pc; // @[Execution.scala 70:21]
  wire [31:0] pipe1_io_uop_npc; // @[Execution.scala 70:21]
  wire [2:0] pipe1_io_uop_fu_code; // @[Execution.scala 70:21]
  wire [3:0] pipe1_io_uop_alu_code; // @[Execution.scala 70:21]
  wire [3:0] pipe1_io_uop_jmp_code; // @[Execution.scala 70:21]
  wire  pipe1_io_uop_w_type; // @[Execution.scala 70:21]
  wire [31:0] pipe1_io_uop_imm; // @[Execution.scala 70:21]
  wire  pipe1_io_uop_pred_br; // @[Execution.scala 70:21]
  wire [31:0] pipe1_io_uop_pred_bpc; // @[Execution.scala 70:21]
  wire [63:0] pipe1_io_in1; // @[Execution.scala 70:21]
  wire [63:0] pipe1_io_in2; // @[Execution.scala 70:21]
  wire  pipe1_io_ecp_jmp_valid; // @[Execution.scala 70:21]
  wire  pipe1_io_ecp_jmp; // @[Execution.scala 70:21]
  wire [31:0] pipe1_io_ecp_jmp_pc; // @[Execution.scala 70:21]
  wire  pipe1_io_ecp_mis; // @[Execution.scala 70:21]
  wire [63:0] pipe1_io_ecp_rd_data; // @[Execution.scala 70:21]
  wire  pipe2_clock; // @[Execution.scala 75:21]
  wire  pipe2_reset; // @[Execution.scala 75:21]
  wire  pipe2_io_uop_valid; // @[Execution.scala 75:21]
  wire [2:0] pipe2_io_uop_fu_code; // @[Execution.scala 75:21]
  wire [1:0] pipe2_io_uop_mem_code; // @[Execution.scala 75:21]
  wire [1:0] pipe2_io_uop_mem_size; // @[Execution.scala 75:21]
  wire [31:0] pipe2_io_uop_imm; // @[Execution.scala 75:21]
  wire [63:0] pipe2_io_in1; // @[Execution.scala 75:21]
  wire [63:0] pipe2_io_in2; // @[Execution.scala 75:21]
  wire  pipe2_io_ecp_store_valid; // @[Execution.scala 75:21]
  wire [63:0] pipe2_io_ecp_rd_data; // @[Execution.scala 75:21]
  wire  pipe2_io_ready; // @[Execution.scala 75:21]
  wire  pipe2_io_dmem_st_req_ready; // @[Execution.scala 75:21]
  wire  pipe2_io_dmem_st_req_valid; // @[Execution.scala 75:21]
  wire [31:0] pipe2_io_dmem_st_req_bits_addr; // @[Execution.scala 75:21]
  wire [63:0] pipe2_io_dmem_st_req_bits_wdata; // @[Execution.scala 75:21]
  wire [7:0] pipe2_io_dmem_st_req_bits_wmask; // @[Execution.scala 75:21]
  wire [1:0] pipe2_io_dmem_st_req_bits_size; // @[Execution.scala 75:21]
  wire  pipe2_io_dmem_st_resp_ready; // @[Execution.scala 75:21]
  wire  pipe2_io_dmem_st_resp_valid; // @[Execution.scala 75:21]
  wire  pipe2_io_dmem_ld_req_ready; // @[Execution.scala 75:21]
  wire  pipe2_io_dmem_ld_req_valid; // @[Execution.scala 75:21]
  wire [31:0] pipe2_io_dmem_ld_req_bits_addr; // @[Execution.scala 75:21]
  wire [1:0] pipe2_io_dmem_ld_req_bits_size; // @[Execution.scala 75:21]
  wire  pipe2_io_dmem_ld_resp_ready; // @[Execution.scala 75:21]
  wire  pipe2_io_dmem_ld_resp_valid; // @[Execution.scala 75:21]
  wire [63:0] pipe2_io_dmem_ld_resp_bits_rdata; // @[Execution.scala 75:21]
  wire  pipe2_io_flush; // @[Execution.scala 75:21]
  wire  pipe2_io_wakeup; // @[Execution.scala 75:21]
  reg  reg_uop_lsu_valid; // @[Execution.scala 32:28]
  reg  reg_uop_lsu_rd_en; // @[Execution.scala 32:28]
  reg [5:0] reg_uop_lsu_rd_paddr; // @[Execution.scala 32:28]
  reg [3:0] reg_uop_lsu_rob_addr; // @[Execution.scala 32:28]
  reg  REG; // @[Execution.scala 33:26]
  wire  reg_valid = REG & io_lsu_ready; // @[Execution.scala 33:42]
  wire [31:0] _T_3 = io_in_0_imm[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_4 = {_T_3,io_in_0_imm}; // @[Cat.scala 30:58]
  wire [63:0] _T_6 = {32'h0,io_in_0_pc}; // @[Cat.scala 30:58]
  wire [63:0] _T_8 = 2'h1 == io_in_0_rs1_src ? io_rs1_data_0 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _T_10 = 2'h2 == io_in_0_rs1_src ? _T_4 : _T_8; // @[Mux.scala 80:57]
  wire [63:0] in1_0_0 = 2'h3 == io_in_0_rs1_src ? _T_6 : _T_10; // @[Mux.scala 80:57]
  wire [63:0] _T_21 = 2'h1 == io_in_0_rs2_src ? io_rs2_data_0 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _T_23 = 2'h2 == io_in_0_rs2_src ? _T_4 : _T_21; // @[Mux.scala 80:57]
  wire [63:0] in2_0_0 = 2'h3 == io_in_0_rs2_src ? _T_6 : _T_23; // @[Mux.scala 80:57]
  wire [63:0] _T_30 = {32'h0,in1_0_0[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_34 = in1_0_0[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_35 = {_T_34,in1_0_0[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_36 = io_in_0_alu_code == 4'h9 ? _T_30 : _T_35; // @[Execution.scala 58:22]
  wire [31:0] _T_41 = in2_0_0[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_42 = {_T_41,in2_0_0[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_46 = io_in_1_imm[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_47 = {_T_46,io_in_1_imm}; // @[Cat.scala 30:58]
  wire [63:0] _T_49 = {32'h0,io_in_1_pc}; // @[Cat.scala 30:58]
  wire [63:0] _T_51 = 2'h1 == io_in_1_rs1_src ? io_rs1_data_1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _T_53 = 2'h2 == io_in_1_rs1_src ? _T_47 : _T_51; // @[Mux.scala 80:57]
  wire [63:0] in1_0_1 = 2'h3 == io_in_1_rs1_src ? _T_49 : _T_53; // @[Mux.scala 80:57]
  wire [63:0] _T_64 = 2'h1 == io_in_1_rs2_src ? io_rs2_data_1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _T_66 = 2'h2 == io_in_1_rs2_src ? _T_47 : _T_64; // @[Mux.scala 80:57]
  wire [63:0] in2_0_1 = 2'h3 == io_in_1_rs2_src ? _T_49 : _T_66; // @[Mux.scala 80:57]
  wire [63:0] _T_73 = {32'h0,in1_0_1[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_77 = in1_0_1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_78 = {_T_77,in1_0_1[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_79 = io_in_1_alu_code == 4'h9 ? _T_73 : _T_78; // @[Execution.scala 58:22]
  wire [31:0] _T_84 = in2_0_1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_85 = {_T_84,in2_0_1[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_89 = io_in_2_imm[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_90 = {_T_89,io_in_2_imm}; // @[Cat.scala 30:58]
  wire [63:0] _T_92 = {32'h0,io_in_2_pc}; // @[Cat.scala 30:58]
  wire [63:0] _T_94 = 2'h1 == io_in_2_rs1_src ? io_rs1_data_2 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _T_96 = 2'h2 == io_in_2_rs1_src ? _T_90 : _T_94; // @[Mux.scala 80:57]
  wire [63:0] in1_0_2 = 2'h3 == io_in_2_rs1_src ? _T_92 : _T_96; // @[Mux.scala 80:57]
  wire [63:0] _T_107 = 2'h1 == io_in_2_rs2_src ? io_rs2_data_2 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _T_109 = 2'h2 == io_in_2_rs2_src ? _T_90 : _T_107; // @[Mux.scala 80:57]
  wire [63:0] in2_0_2 = 2'h3 == io_in_2_rs2_src ? _T_92 : _T_109; // @[Mux.scala 80:57]
  wire [63:0] _T_116 = {32'h0,in1_0_2[31:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_120 = in1_0_2[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_121 = {_T_120,in1_0_2[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_122 = io_in_2_alu_code == 4'h9 ? _T_116 : _T_121; // @[Execution.scala 58:22]
  wire [31:0] _T_127 = in2_0_2[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_128 = {_T_127,in2_0_2[31:0]}; // @[Cat.scala 30:58]
  reg  out_uop_0_valid; // @[Execution.scala 92:24]
  reg [3:0] out_uop_0_rob_addr; // @[Execution.scala 92:24]
  reg  out_uop_1_valid; // @[Execution.scala 92:24]
  reg [3:0] out_uop_1_rob_addr; // @[Execution.scala 92:24]
  reg  out_uop_2_valid; // @[Execution.scala 92:24]
  reg [3:0] out_uop_2_rob_addr; // @[Execution.scala 92:24]
  reg  out_ecp_0_jmp_valid; // @[Execution.scala 93:24]
  reg  out_ecp_0_jmp; // @[Execution.scala 93:24]
  reg [31:0] out_ecp_0_jmp_pc; // @[Execution.scala 93:24]
  reg  out_ecp_0_mis; // @[Execution.scala 93:24]
  reg  out_ecp_1_jmp_valid; // @[Execution.scala 93:24]
  reg  out_ecp_1_jmp; // @[Execution.scala 93:24]
  reg [31:0] out_ecp_1_jmp_pc; // @[Execution.scala 93:24]
  reg  out_ecp_1_mis; // @[Execution.scala 93:24]
  reg  out_ecp_2_store_valid; // @[Execution.scala 93:24]
  wire  _T_130_rd_en = reg_valid & reg_uop_lsu_rd_en; // @[Execution.scala 123:27]
  ysyx_210128_ExPipe0 pipe0 ( // @[Execution.scala 65:21]
    .clock(pipe0_clock),
    .reset(pipe0_reset),
    .io_uop_valid(pipe0_io_uop_valid),
    .io_uop_pc(pipe0_io_uop_pc),
    .io_uop_npc(pipe0_io_uop_npc),
    .io_uop_inst(pipe0_io_uop_inst),
    .io_uop_fu_code(pipe0_io_uop_fu_code),
    .io_uop_alu_code(pipe0_io_uop_alu_code),
    .io_uop_jmp_code(pipe0_io_uop_jmp_code),
    .io_uop_sys_code(pipe0_io_uop_sys_code),
    .io_uop_w_type(pipe0_io_uop_w_type),
    .io_uop_imm(pipe0_io_uop_imm),
    .io_uop_pred_br(pipe0_io_uop_pred_br),
    .io_uop_pred_bpc(pipe0_io_uop_pred_bpc),
    .io_in1(pipe0_io_in1),
    .io_in2(pipe0_io_in2),
    .io_ecp_jmp_valid(pipe0_io_ecp_jmp_valid),
    .io_ecp_jmp(pipe0_io_ecp_jmp),
    .io_ecp_jmp_pc(pipe0_io_ecp_jmp_pc),
    .io_ecp_mis(pipe0_io_ecp_mis),
    .io_ecp_rd_data(pipe0_io_ecp_rd_data),
    .mtip(pipe0_mtip),
    .intr_mcause(pipe0_intr_mcause),
    .instr_cnt(pipe0_instr_cnt),
    .intr_mstatus(pipe0_intr_mstatus),
    ._T_6_0(pipe0__T_6_0),
    ._T_5_0(pipe0__T_5_0),
    .intr(pipe0_intr),
    .fence_i(pipe0_fence_i),
    .cycle_cnt(pipe0_cycle_cnt),
    .mstatus(pipe0_mstatus),
    .intr_mepc(pipe0_intr_mepc),
    .mtip_0(pipe0_mtip_0)
  );
  ysyx_210128_ExPipe1 pipe1 ( // @[Execution.scala 70:21]
    .io_uop_pc(pipe1_io_uop_pc),
    .io_uop_npc(pipe1_io_uop_npc),
    .io_uop_fu_code(pipe1_io_uop_fu_code),
    .io_uop_alu_code(pipe1_io_uop_alu_code),
    .io_uop_jmp_code(pipe1_io_uop_jmp_code),
    .io_uop_w_type(pipe1_io_uop_w_type),
    .io_uop_imm(pipe1_io_uop_imm),
    .io_uop_pred_br(pipe1_io_uop_pred_br),
    .io_uop_pred_bpc(pipe1_io_uop_pred_bpc),
    .io_in1(pipe1_io_in1),
    .io_in2(pipe1_io_in2),
    .io_ecp_jmp_valid(pipe1_io_ecp_jmp_valid),
    .io_ecp_jmp(pipe1_io_ecp_jmp),
    .io_ecp_jmp_pc(pipe1_io_ecp_jmp_pc),
    .io_ecp_mis(pipe1_io_ecp_mis),
    .io_ecp_rd_data(pipe1_io_ecp_rd_data)
  );
  ysyx_210128_ExPipe2 pipe2 ( // @[Execution.scala 75:21]
    .clock(pipe2_clock),
    .reset(pipe2_reset),
    .io_uop_valid(pipe2_io_uop_valid),
    .io_uop_fu_code(pipe2_io_uop_fu_code),
    .io_uop_mem_code(pipe2_io_uop_mem_code),
    .io_uop_mem_size(pipe2_io_uop_mem_size),
    .io_uop_imm(pipe2_io_uop_imm),
    .io_in1(pipe2_io_in1),
    .io_in2(pipe2_io_in2),
    .io_ecp_store_valid(pipe2_io_ecp_store_valid),
    .io_ecp_rd_data(pipe2_io_ecp_rd_data),
    .io_ready(pipe2_io_ready),
    .io_dmem_st_req_ready(pipe2_io_dmem_st_req_ready),
    .io_dmem_st_req_valid(pipe2_io_dmem_st_req_valid),
    .io_dmem_st_req_bits_addr(pipe2_io_dmem_st_req_bits_addr),
    .io_dmem_st_req_bits_wdata(pipe2_io_dmem_st_req_bits_wdata),
    .io_dmem_st_req_bits_wmask(pipe2_io_dmem_st_req_bits_wmask),
    .io_dmem_st_req_bits_size(pipe2_io_dmem_st_req_bits_size),
    .io_dmem_st_resp_ready(pipe2_io_dmem_st_resp_ready),
    .io_dmem_st_resp_valid(pipe2_io_dmem_st_resp_valid),
    .io_dmem_ld_req_ready(pipe2_io_dmem_ld_req_ready),
    .io_dmem_ld_req_valid(pipe2_io_dmem_ld_req_valid),
    .io_dmem_ld_req_bits_addr(pipe2_io_dmem_ld_req_bits_addr),
    .io_dmem_ld_req_bits_size(pipe2_io_dmem_ld_req_bits_size),
    .io_dmem_ld_resp_ready(pipe2_io_dmem_ld_resp_ready),
    .io_dmem_ld_resp_valid(pipe2_io_dmem_ld_resp_valid),
    .io_dmem_ld_resp_bits_rdata(pipe2_io_dmem_ld_resp_bits_rdata),
    .io_flush(pipe2_io_flush),
    .io_wakeup(pipe2_io_wakeup)
  );
  assign io_out_0_valid = out_uop_0_valid; // @[Execution.scala 130:15]
  assign io_out_0_rob_addr = out_uop_0_rob_addr; // @[Execution.scala 130:15]
  assign io_out_1_valid = out_uop_1_valid; // @[Execution.scala 130:15]
  assign io_out_1_rob_addr = out_uop_1_rob_addr; // @[Execution.scala 130:15]
  assign io_out_2_valid = out_uop_2_valid; // @[Execution.scala 130:15]
  assign io_out_2_rob_addr = out_uop_2_rob_addr; // @[Execution.scala 130:15]
  assign io_out_ecp_0_jmp_valid = out_ecp_0_jmp_valid; // @[Execution.scala 131:15]
  assign io_out_ecp_0_jmp = out_ecp_0_jmp; // @[Execution.scala 131:15]
  assign io_out_ecp_0_jmp_pc = out_ecp_0_jmp_pc; // @[Execution.scala 131:15]
  assign io_out_ecp_0_mis = out_ecp_0_mis; // @[Execution.scala 131:15]
  assign io_out_ecp_1_jmp_valid = out_ecp_1_jmp_valid; // @[Execution.scala 131:15]
  assign io_out_ecp_1_jmp = out_ecp_1_jmp; // @[Execution.scala 131:15]
  assign io_out_ecp_1_jmp_pc = out_ecp_1_jmp_pc; // @[Execution.scala 131:15]
  assign io_out_ecp_1_mis = out_ecp_1_mis; // @[Execution.scala 131:15]
  assign io_out_ecp_2_store_valid = out_ecp_2_store_valid; // @[Execution.scala 131:15]
  assign io_rd_en_0 = io_flush ? 1'h0 : io_in_0_rd_en; // @[Execution.scala 98:19 102:20 111:21]
  assign io_rd_en_1 = io_flush ? 1'h0 : io_in_1_rd_en; // @[Execution.scala 98:19 102:20 118:21]
  assign io_rd_en_2 = io_flush ? 1'h0 : _T_130_rd_en; // @[Execution.scala 98:19 102:20 125:21]
  assign io_rd_paddr_0 = io_flush ? 6'h0 : io_in_0_rd_paddr; // @[Execution.scala 98:19 103:23 112:21]
  assign io_rd_paddr_1 = io_flush ? 6'h0 : io_in_1_rd_paddr; // @[Execution.scala 98:19 103:23 119:21]
  assign io_rd_paddr_2 = io_flush ? 6'h0 : reg_uop_lsu_rd_paddr; // @[Execution.scala 98:19 103:23 126:21]
  assign io_rd_data_0 = io_flush ? 64'h0 : pipe0_io_ecp_rd_data; // @[Execution.scala 98:19 104:22 113:21]
  assign io_rd_data_1 = io_flush ? 64'h0 : pipe1_io_ecp_rd_data; // @[Execution.scala 98:19 104:22 120:21]
  assign io_rd_data_2 = io_flush ? 64'h0 : pipe2_io_ecp_rd_data; // @[Execution.scala 98:19 104:22 127:21]
  assign io_lsu_ready = pipe2_io_ready; // @[Execution.scala 79:16]
  assign io_dmem_st_req_valid = pipe2_io_dmem_st_req_valid; // @[Execution.scala 80:20]
  assign io_dmem_st_req_bits_addr = pipe2_io_dmem_st_req_bits_addr; // @[Execution.scala 80:20]
  assign io_dmem_st_req_bits_wdata = pipe2_io_dmem_st_req_bits_wdata; // @[Execution.scala 80:20]
  assign io_dmem_st_req_bits_wmask = pipe2_io_dmem_st_req_bits_wmask; // @[Execution.scala 80:20]
  assign io_dmem_st_req_bits_size = pipe2_io_dmem_st_req_bits_size; // @[Execution.scala 80:20]
  assign io_dmem_st_resp_ready = pipe2_io_dmem_st_resp_ready; // @[Execution.scala 80:20]
  assign io_dmem_ld_req_valid = pipe2_io_dmem_ld_req_valid; // @[Execution.scala 81:20]
  assign io_dmem_ld_req_bits_addr = pipe2_io_dmem_ld_req_bits_addr; // @[Execution.scala 81:20]
  assign io_dmem_ld_req_bits_size = pipe2_io_dmem_ld_req_bits_size; // @[Execution.scala 81:20]
  assign io_dmem_ld_resp_ready = pipe2_io_dmem_ld_resp_ready; // @[Execution.scala 81:20]
  assign io_lsu_wakeup_uop_valid = pipe2_io_wakeup & reg_uop_lsu_valid; // @[Execution.scala 85:21 86:26 87:23]
  assign io_lsu_wakeup_uop_rd_en = pipe2_io_wakeup & reg_uop_lsu_rd_en; // @[Execution.scala 85:21 86:26 87:23]
  assign io_lsu_wakeup_uop_rd_paddr = pipe2_io_wakeup ? reg_uop_lsu_rd_paddr : 6'h0; // @[Execution.scala 85:21 86:26 87:23]
  assign mtip = pipe0_mtip;
  assign _T_6_0 = pipe0__T_6_0;
  assign _T_5_0 = pipe0__T_5_0;
  assign fence_i = pipe0_fence_i;
  assign mstatus = pipe0_mstatus;
  assign pipe0_clock = clock;
  assign pipe0_reset = reset;
  assign pipe0_io_uop_valid = io_in_0_valid; // @[Execution.scala 66:16]
  assign pipe0_io_uop_pc = io_in_0_pc; // @[Execution.scala 66:16]
  assign pipe0_io_uop_npc = io_in_0_npc; // @[Execution.scala 66:16]
  assign pipe0_io_uop_inst = io_in_0_inst; // @[Execution.scala 66:16]
  assign pipe0_io_uop_fu_code = io_in_0_fu_code; // @[Execution.scala 66:16]
  assign pipe0_io_uop_alu_code = io_in_0_alu_code; // @[Execution.scala 66:16]
  assign pipe0_io_uop_jmp_code = io_in_0_jmp_code; // @[Execution.scala 66:16]
  assign pipe0_io_uop_sys_code = io_in_0_sys_code; // @[Execution.scala 66:16]
  assign pipe0_io_uop_w_type = io_in_0_w_type; // @[Execution.scala 66:16]
  assign pipe0_io_uop_imm = io_in_0_imm; // @[Execution.scala 66:16]
  assign pipe0_io_uop_pred_br = io_in_0_pred_br; // @[Execution.scala 66:16]
  assign pipe0_io_uop_pred_bpc = io_in_0_pred_bpc; // @[Execution.scala 66:16]
  assign pipe0_io_in1 = io_in_0_w_type ? _T_36 : in1_0_0; // @[Execution.scala 57:18]
  assign pipe0_io_in2 = io_in_0_w_type ? _T_42 : in2_0_0; // @[Execution.scala 62:18]
  assign pipe0_intr_mcause = intr_mcause;
  assign pipe0_instr_cnt = instr_cnt;
  assign pipe0_intr_mstatus = intr_mstatus;
  assign pipe0_intr = intr;
  assign pipe0_cycle_cnt = cycle_cnt;
  assign pipe0_intr_mepc = intr_mepc;
  assign pipe0_mtip_0 = mtip_0;
  assign pipe1_io_uop_pc = io_in_1_pc; // @[Execution.scala 71:16]
  assign pipe1_io_uop_npc = io_in_1_npc; // @[Execution.scala 71:16]
  assign pipe1_io_uop_fu_code = io_in_1_fu_code; // @[Execution.scala 71:16]
  assign pipe1_io_uop_alu_code = io_in_1_alu_code; // @[Execution.scala 71:16]
  assign pipe1_io_uop_jmp_code = io_in_1_jmp_code; // @[Execution.scala 71:16]
  assign pipe1_io_uop_w_type = io_in_1_w_type; // @[Execution.scala 71:16]
  assign pipe1_io_uop_imm = io_in_1_imm; // @[Execution.scala 71:16]
  assign pipe1_io_uop_pred_br = io_in_1_pred_br; // @[Execution.scala 71:16]
  assign pipe1_io_uop_pred_bpc = io_in_1_pred_bpc; // @[Execution.scala 71:16]
  assign pipe1_io_in1 = io_in_1_w_type ? _T_79 : in1_0_1; // @[Execution.scala 57:18]
  assign pipe1_io_in2 = io_in_1_w_type ? _T_85 : in2_0_1; // @[Execution.scala 62:18]
  assign pipe2_clock = clock;
  assign pipe2_reset = reset;
  assign pipe2_io_uop_valid = io_in_2_valid; // @[Execution.scala 76:16]
  assign pipe2_io_uop_fu_code = io_in_2_fu_code; // @[Execution.scala 76:16]
  assign pipe2_io_uop_mem_code = io_in_2_mem_code; // @[Execution.scala 76:16]
  assign pipe2_io_uop_mem_size = io_in_2_mem_size; // @[Execution.scala 76:16]
  assign pipe2_io_uop_imm = io_in_2_imm; // @[Execution.scala 76:16]
  assign pipe2_io_in1 = io_in_2_w_type ? _T_122 : in1_0_2; // @[Execution.scala 57:18]
  assign pipe2_io_in2 = io_in_2_w_type ? _T_128 : in2_0_2; // @[Execution.scala 62:18]
  assign pipe2_io_dmem_st_req_ready = io_dmem_st_req_ready; // @[Execution.scala 80:20]
  assign pipe2_io_dmem_st_resp_valid = io_dmem_st_resp_valid; // @[Execution.scala 80:20]
  assign pipe2_io_dmem_ld_req_ready = io_dmem_ld_req_ready; // @[Execution.scala 81:20]
  assign pipe2_io_dmem_ld_resp_valid = io_dmem_ld_resp_valid; // @[Execution.scala 81:20]
  assign pipe2_io_dmem_ld_resp_bits_rdata = io_dmem_ld_resp_bits_rdata; // @[Execution.scala 81:20]
  assign pipe2_io_flush = io_flush; // @[Execution.scala 82:18]
  always @(posedge clock) begin
    if (reset) begin // @[Execution.scala 32:28]
      reg_uop_lsu_valid <= 1'h0; // @[Execution.scala 32:28]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      reg_uop_lsu_valid <= 1'h0; // @[Execution.scala 106:17]
    end else if (io_in_2_valid) begin // @[Execution.scala 35:36]
      reg_uop_lsu_valid <= io_in_2_valid; // @[Execution.scala 36:17]
    end
    if (reset) begin // @[Execution.scala 32:28]
      reg_uop_lsu_rd_en <= 1'h0; // @[Execution.scala 32:28]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      reg_uop_lsu_rd_en <= 1'h0; // @[Execution.scala 106:17]
    end else if (io_in_2_valid) begin // @[Execution.scala 35:36]
      reg_uop_lsu_rd_en <= io_in_2_rd_en; // @[Execution.scala 36:17]
    end
    if (reset) begin // @[Execution.scala 32:28]
      reg_uop_lsu_rd_paddr <= 6'h0; // @[Execution.scala 32:28]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      reg_uop_lsu_rd_paddr <= 6'h0; // @[Execution.scala 106:17]
    end else if (io_in_2_valid) begin // @[Execution.scala 35:36]
      reg_uop_lsu_rd_paddr <= io_in_2_rd_paddr; // @[Execution.scala 36:17]
    end
    if (reset) begin // @[Execution.scala 32:28]
      reg_uop_lsu_rob_addr <= 4'h0; // @[Execution.scala 32:28]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      reg_uop_lsu_rob_addr <= 4'h0; // @[Execution.scala 106:17]
    end else if (io_in_2_valid) begin // @[Execution.scala 35:36]
      reg_uop_lsu_rob_addr <= io_in_2_rob_addr; // @[Execution.scala 36:17]
    end
    REG <= ~io_lsu_ready; // @[Execution.scala 33:27]
    if (reset) begin // @[Execution.scala 92:24]
      out_uop_0_valid <= 1'h0; // @[Execution.scala 92:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_uop_0_valid <= 1'h0; // @[Execution.scala 100:18]
    end else begin
      out_uop_0_valid <= io_in_0_valid; // @[Execution.scala 109:21]
    end
    if (reset) begin // @[Execution.scala 92:24]
      out_uop_0_rob_addr <= 4'h0; // @[Execution.scala 92:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_uop_0_rob_addr <= 4'h0; // @[Execution.scala 100:18]
    end else begin
      out_uop_0_rob_addr <= io_in_0_rob_addr; // @[Execution.scala 109:21]
    end
    if (reset) begin // @[Execution.scala 92:24]
      out_uop_1_valid <= 1'h0; // @[Execution.scala 92:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_uop_1_valid <= 1'h0; // @[Execution.scala 100:18]
    end else begin
      out_uop_1_valid <= io_in_1_valid; // @[Execution.scala 116:21]
    end
    if (reset) begin // @[Execution.scala 92:24]
      out_uop_1_rob_addr <= 4'h0; // @[Execution.scala 92:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_uop_1_rob_addr <= 4'h0; // @[Execution.scala 100:18]
    end else begin
      out_uop_1_rob_addr <= io_in_1_rob_addr; // @[Execution.scala 116:21]
    end
    if (reset) begin // @[Execution.scala 92:24]
      out_uop_2_valid <= 1'h0; // @[Execution.scala 92:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_uop_2_valid <= 1'h0; // @[Execution.scala 100:18]
    end else begin
      out_uop_2_valid <= reg_valid & reg_uop_lsu_valid; // @[Execution.scala 123:21]
    end
    if (reset) begin // @[Execution.scala 92:24]
      out_uop_2_rob_addr <= 4'h0; // @[Execution.scala 92:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_uop_2_rob_addr <= 4'h0; // @[Execution.scala 100:18]
    end else if (reg_valid) begin // @[Execution.scala 123:27]
      out_uop_2_rob_addr <= reg_uop_lsu_rob_addr;
    end else begin
      out_uop_2_rob_addr <= 4'h0;
    end
    if (reset) begin // @[Execution.scala 93:24]
      out_ecp_0_jmp_valid <= 1'h0; // @[Execution.scala 93:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_ecp_0_jmp_valid <= 1'h0; // @[Execution.scala 101:18]
    end else begin
      out_ecp_0_jmp_valid <= pipe0_io_ecp_jmp_valid; // @[Execution.scala 110:21]
    end
    if (reset) begin // @[Execution.scala 93:24]
      out_ecp_0_jmp <= 1'h0; // @[Execution.scala 93:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_ecp_0_jmp <= 1'h0; // @[Execution.scala 101:18]
    end else begin
      out_ecp_0_jmp <= pipe0_io_ecp_jmp; // @[Execution.scala 110:21]
    end
    if (reset) begin // @[Execution.scala 93:24]
      out_ecp_0_jmp_pc <= 32'h0; // @[Execution.scala 93:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_ecp_0_jmp_pc <= 32'h0; // @[Execution.scala 101:18]
    end else begin
      out_ecp_0_jmp_pc <= pipe0_io_ecp_jmp_pc; // @[Execution.scala 110:21]
    end
    if (reset) begin // @[Execution.scala 93:24]
      out_ecp_0_mis <= 1'h0; // @[Execution.scala 93:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_ecp_0_mis <= 1'h0; // @[Execution.scala 101:18]
    end else begin
      out_ecp_0_mis <= pipe0_io_ecp_mis; // @[Execution.scala 110:21]
    end
    if (reset) begin // @[Execution.scala 93:24]
      out_ecp_1_jmp_valid <= 1'h0; // @[Execution.scala 93:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_ecp_1_jmp_valid <= 1'h0; // @[Execution.scala 101:18]
    end else begin
      out_ecp_1_jmp_valid <= pipe1_io_ecp_jmp_valid; // @[Execution.scala 117:21]
    end
    if (reset) begin // @[Execution.scala 93:24]
      out_ecp_1_jmp <= 1'h0; // @[Execution.scala 93:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_ecp_1_jmp <= 1'h0; // @[Execution.scala 101:18]
    end else begin
      out_ecp_1_jmp <= pipe1_io_ecp_jmp; // @[Execution.scala 117:21]
    end
    if (reset) begin // @[Execution.scala 93:24]
      out_ecp_1_jmp_pc <= 32'h0; // @[Execution.scala 93:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_ecp_1_jmp_pc <= 32'h0; // @[Execution.scala 101:18]
    end else begin
      out_ecp_1_jmp_pc <= pipe1_io_ecp_jmp_pc; // @[Execution.scala 117:21]
    end
    if (reset) begin // @[Execution.scala 93:24]
      out_ecp_1_mis <= 1'h0; // @[Execution.scala 93:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_ecp_1_mis <= 1'h0; // @[Execution.scala 101:18]
    end else begin
      out_ecp_1_mis <= pipe1_io_ecp_mis; // @[Execution.scala 117:21]
    end
    if (reset) begin // @[Execution.scala 93:24]
      out_ecp_2_store_valid <= 1'h0; // @[Execution.scala 93:24]
    end else if (io_flush) begin // @[Execution.scala 98:19]
      out_ecp_2_store_valid <= 1'h0; // @[Execution.scala 101:18]
    end else begin
      out_ecp_2_store_valid <= pipe2_io_ecp_store_valid; // @[Execution.scala 124:21]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_uop_lsu_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_uop_lsu_rd_en = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  reg_uop_lsu_rd_paddr = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  reg_uop_lsu_rob_addr = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_uop_0_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  out_uop_0_rob_addr = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  out_uop_1_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  out_uop_1_rob_addr = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  out_uop_2_valid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  out_uop_2_rob_addr = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  out_ecp_0_jmp_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  out_ecp_0_jmp = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  out_ecp_0_jmp_pc = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  out_ecp_0_mis = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  out_ecp_1_jmp_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  out_ecp_1_jmp = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  out_ecp_1_jmp_pc = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  out_ecp_1_mis = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  out_ecp_2_store_valid = _RAND_19[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_StoreQueue(
  input         clock,
  input         reset,
  input         io_flush,
  output        io_in_st_req_ready,
  input         io_in_st_req_valid,
  input  [31:0] io_in_st_req_bits_addr,
  input  [63:0] io_in_st_req_bits_wdata,
  input  [7:0]  io_in_st_req_bits_wmask,
  input  [1:0]  io_in_st_req_bits_size,
  input         io_in_st_resp_ready,
  output        io_in_st_resp_valid,
  output        io_in_ld_req_ready,
  input         io_in_ld_req_valid,
  input  [31:0] io_in_ld_req_bits_addr,
  input  [1:0]  io_in_ld_req_bits_size,
  input         io_in_ld_resp_ready,
  output        io_in_ld_resp_valid,
  output [63:0] io_in_ld_resp_bits_rdata,
  input         io_out_st_req_ready,
  output        io_out_st_req_valid,
  output [31:0] io_out_st_req_bits_addr,
  output [63:0] io_out_st_req_bits_wdata,
  output [7:0]  io_out_st_req_bits_wmask,
  output [1:0]  io_out_st_req_bits_size,
  output        io_out_st_resp_ready,
  input         io_out_st_resp_valid,
  input         io_out_ld_req_ready,
  output        io_out_ld_req_valid,
  output [31:0] io_out_ld_req_bits_addr,
  output [1:0]  io_out_ld_req_bits_size,
  output        io_out_ld_resp_ready,
  input         io_out_ld_resp_valid,
  input  [63:0] io_out_ld_resp_bits_rdata,
  input         io_deq_req,
  output        empty_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] sq_0_addr; // @[StoreQueue.scala 31:19]
  reg [63:0] sq_0_wdata; // @[StoreQueue.scala 31:19]
  reg [7:0] sq_0_wmask; // @[StoreQueue.scala 31:19]
  reg [1:0] sq_0_wsize; // @[StoreQueue.scala 31:19]
  reg  sq_0_valid; // @[StoreQueue.scala 31:19]
  reg [31:0] sq_1_addr; // @[StoreQueue.scala 31:19]
  reg [63:0] sq_1_wdata; // @[StoreQueue.scala 31:19]
  reg [7:0] sq_1_wmask; // @[StoreQueue.scala 31:19]
  reg [1:0] sq_1_wsize; // @[StoreQueue.scala 31:19]
  reg  sq_1_valid; // @[StoreQueue.scala 31:19]
  reg [31:0] sq_2_addr; // @[StoreQueue.scala 31:19]
  reg [63:0] sq_2_wdata; // @[StoreQueue.scala 31:19]
  reg [7:0] sq_2_wmask; // @[StoreQueue.scala 31:19]
  reg [1:0] sq_2_wsize; // @[StoreQueue.scala 31:19]
  reg  sq_2_valid; // @[StoreQueue.scala 31:19]
  reg [31:0] sq_3_addr; // @[StoreQueue.scala 31:19]
  reg [63:0] sq_3_wdata; // @[StoreQueue.scala 31:19]
  reg [7:0] sq_3_wmask; // @[StoreQueue.scala 31:19]
  reg [1:0] sq_3_wsize; // @[StoreQueue.scala 31:19]
  reg  sq_3_valid; // @[StoreQueue.scala 31:19]
  reg [1:0] value; // @[Counter.scala 60:40]
  reg [1:0] value_1; // @[Counter.scala 60:40]
  reg  maybe_full; // @[StoreQueue.scala 34:27]
  wire  _T = value == value_1; // @[StoreQueue.scala 35:30]
  wire  empty = value == value_1 & ~maybe_full; // @[StoreQueue.scala 35:49]
  wire  full = _T & maybe_full; // @[StoreQueue.scala 36:48]
  reg  deq_state; // @[StoreQueue.scala 43:26]
  reg  enq_state; // @[StoreQueue.scala 46:26]
  reg  flush_state; // @[StoreQueue.scala 49:28]
  reg [2:0] deq_req_counter; // @[StoreQueue.scala 55:32]
  wire  deq_req_empty = deq_req_counter == 3'h0; // @[StoreQueue.scala 56:40]
  wire  deq_valid = ~empty & ~deq_req_empty; // @[StoreQueue.scala 59:26]
  wire  _T_5 = ~deq_state; // @[StoreQueue.scala 60:53]
  wire  deq_ready = io_out_st_req_ready & ~deq_state; // @[StoreQueue.scala 60:39]
  wire  deq_fire = deq_valid & deq_ready; // @[StoreQueue.scala 61:25]
  wire [2:0] _T_10 = deq_req_counter + 3'h1; // @[StoreQueue.scala 64:40]
  wire  _T_11 = ~io_deq_req; // @[StoreQueue.scala 65:16]
  wire [2:0] _T_14 = deq_req_counter - 3'h1; // @[StoreQueue.scala 66:40]
  wire  _GEN_2 = 2'h0 == value_1 ? 1'h0 : sq_0_valid; // @[StoreQueue.scala 31:19 70:{29,29}]
  wire  _GEN_3 = 2'h1 == value_1 ? 1'h0 : sq_1_valid; // @[StoreQueue.scala 31:19 70:{29,29}]
  wire  _GEN_4 = 2'h2 == value_1 ? 1'h0 : sq_2_valid; // @[StoreQueue.scala 31:19 70:{29,29}]
  wire  _GEN_5 = 2'h3 == value_1 ? 1'h0 : sq_3_valid; // @[StoreQueue.scala 31:19 70:{29,29}]
  wire [1:0] _value_T_1 = value_1 + 2'h1; // @[Counter.scala 76:24]
  wire  _GEN_6 = deq_fire ? _GEN_2 : sq_0_valid; // @[StoreQueue.scala 31:19 69:19]
  wire  _GEN_7 = deq_fire ? _GEN_3 : sq_1_valid; // @[StoreQueue.scala 31:19 69:19]
  wire  _GEN_8 = deq_fire ? _GEN_4 : sq_2_valid; // @[StoreQueue.scala 31:19 69:19]
  wire  _GEN_9 = deq_fire ? _GEN_5 : sq_3_valid; // @[StoreQueue.scala 31:19 69:19]
  wire [1:0] _GEN_10 = deq_fire ? _value_T_1 : value_1; // @[StoreQueue.scala 69:19 Counter.scala 76:15 60:40]
  wire  _GEN_11 = deq_fire | deq_state; // @[StoreQueue.scala 81:23 82:19 43:26]
  wire  _T_17 = io_out_st_resp_ready & io_out_st_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_20 = ~enq_state; // @[StoreQueue.scala 95:53]
  wire  _T_22 = ~flush_state; // @[StoreQueue.scala 95:83]
  wire  enq_ready = (~full | deq_fire) & ~enq_state & ~flush_state; // @[StoreQueue.scala 95:67]
  wire  enq_fire = io_in_st_req_valid & enq_ready; // @[StoreQueue.scala 96:28]
  wire  _GEN_15 = 2'h0 == value | _GEN_6; // @[StoreQueue.scala 105:{23,23}]
  wire  _GEN_16 = 2'h1 == value | _GEN_7; // @[StoreQueue.scala 105:{23,23}]
  wire  _GEN_17 = 2'h2 == value | _GEN_8; // @[StoreQueue.scala 105:{23,23}]
  wire  _GEN_18 = 2'h3 == value | _GEN_9; // @[StoreQueue.scala 105:{23,23}]
  wire [1:0] _value_T_3 = value + 2'h1; // @[Counter.scala 76:24]
  wire  _GEN_35 = enq_fire ? _GEN_15 : _GEN_6; // @[StoreQueue.scala 98:19]
  wire  _GEN_36 = enq_fire ? _GEN_16 : _GEN_7; // @[StoreQueue.scala 98:19]
  wire  _GEN_37 = enq_fire ? _GEN_17 : _GEN_8; // @[StoreQueue.scala 98:19]
  wire  _GEN_38 = enq_fire ? _GEN_18 : _GEN_9; // @[StoreQueue.scala 98:19]
  wire [1:0] _GEN_55 = enq_fire ? _value_T_3 : value; // @[Counter.scala 76:15 StoreQueue.scala 98:19 Counter.scala 60:40]
  wire  _GEN_56 = enq_fire | enq_state; // @[StoreQueue.scala 116:23 117:19 46:26]
  wire  _T_25 = io_in_st_resp_ready & io_in_st_resp_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_60 = enq_fire != deq_fire ? enq_fire : maybe_full; // @[StoreQueue.scala 127:32 128:16 34:27]
  wire  load_addr_match_0 = sq_0_valid & sq_0_addr == io_in_ld_req_bits_addr; // @[StoreQueue.scala 136:39]
  wire  load_addr_match_1 = sq_1_valid & sq_1_addr == io_in_ld_req_bits_addr; // @[StoreQueue.scala 136:39]
  wire  load_addr_match_2 = sq_2_valid & sq_2_addr == io_in_ld_req_bits_addr; // @[StoreQueue.scala 136:39]
  wire  load_addr_match_3 = sq_3_valid & sq_3_addr == io_in_ld_req_bits_addr; // @[StoreQueue.scala 136:39]
  wire [3:0] _T_35 = {load_addr_match_3,load_addr_match_2,load_addr_match_1,load_addr_match_0}; // @[Cat.scala 30:58]
  wire  load_hit = |_T_35; // @[StoreQueue.scala 139:47]
  wire  _T_40 = ~load_hit; // @[StoreQueue.scala 185:54]
  wire [31:0] _GEN_102 = 2'h1 == value_1 ? sq_1_addr : sq_0_addr; // @[StoreQueue.scala 196:{28,28}]
  wire [31:0] _GEN_103 = 2'h2 == value_1 ? sq_2_addr : _GEN_102; // @[StoreQueue.scala 196:{28,28}]
  wire [63:0] _GEN_106 = 2'h1 == value_1 ? sq_1_wdata : sq_0_wdata; // @[StoreQueue.scala 197:{28,28}]
  wire [63:0] _GEN_107 = 2'h2 == value_1 ? sq_2_wdata : _GEN_106; // @[StoreQueue.scala 197:{28,28}]
  wire [7:0] _GEN_110 = 2'h1 == value_1 ? sq_1_wmask : sq_0_wmask; // @[StoreQueue.scala 198:{28,28}]
  wire [7:0] _GEN_111 = 2'h2 == value_1 ? sq_2_wmask : _GEN_110; // @[StoreQueue.scala 198:{28,28}]
  wire [1:0] _GEN_114 = 2'h1 == value_1 ? sq_1_wsize : sq_0_wsize; // @[StoreQueue.scala 200:{28,28}]
  wire [1:0] _GEN_115 = 2'h2 == value_1 ? sq_2_wsize : _GEN_114; // @[StoreQueue.scala 200:{28,28}]
  assign io_in_st_req_ready = (~full | deq_fire) & ~enq_state & ~flush_state; // @[StoreQueue.scala 95:67]
  assign io_in_st_resp_valid = enq_state; // @[StoreQueue.scala 187:42]
  assign io_in_ld_req_ready = io_out_ld_req_ready & ~load_hit & _T_22; // @[StoreQueue.scala 185:64]
  assign io_in_ld_resp_valid = io_out_ld_resp_valid; // @[StoreQueue.scala 191:28]
  assign io_in_ld_resp_bits_rdata = io_out_ld_resp_bits_rdata; // @[StoreQueue.scala 192:28]
  assign io_out_st_req_valid = deq_valid & _T_5; // @[StoreQueue.scala 195:41]
  assign io_out_st_req_bits_addr = 2'h3 == value_1 ? sq_3_addr : _GEN_103; // @[StoreQueue.scala 196:{28,28}]
  assign io_out_st_req_bits_wdata = 2'h3 == value_1 ? sq_3_wdata : _GEN_107; // @[StoreQueue.scala 197:{28,28}]
  assign io_out_st_req_bits_wmask = 2'h3 == value_1 ? sq_3_wmask : _GEN_111; // @[StoreQueue.scala 198:{28,28}]
  assign io_out_st_req_bits_size = 2'h3 == value_1 ? sq_3_wsize : _GEN_115; // @[StoreQueue.scala 200:{28,28}]
  assign io_out_st_resp_ready = deq_state; // @[StoreQueue.scala 203:42]
  assign io_out_ld_req_valid = io_in_ld_req_valid & _T_40 & _T_22; // @[StoreQueue.scala 205:89]
  assign io_out_ld_req_bits_addr = io_in_ld_req_bits_addr; // @[StoreQueue.scala 206:28]
  assign io_out_ld_req_bits_size = io_in_ld_req_bits_size; // @[StoreQueue.scala 210:28]
  assign io_out_ld_resp_ready = io_in_ld_resp_ready; // @[StoreQueue.scala 213:28]
  assign empty_0 = empty;
  always @(posedge clock) begin
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_0_addr <= 32'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h0 == value) begin // @[StoreQueue.scala 105:23]
        sq_0_addr <= io_in_st_req_bits_addr; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_0_wdata <= 64'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h0 == value) begin // @[StoreQueue.scala 105:23]
        sq_0_wdata <= io_in_st_req_bits_wdata; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_0_wmask <= 8'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h0 == value) begin // @[StoreQueue.scala 105:23]
        sq_0_wmask <= io_in_st_req_bits_wmask; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_0_wsize <= 2'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h0 == value) begin // @[StoreQueue.scala 105:23]
        sq_0_wsize <= io_in_st_req_bits_size; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_0_valid <= 1'h0; // @[StoreQueue.scala 31:19]
    end else if (_T_22) begin // @[StoreQueue.scala 153:24]
      if (io_flush) begin // @[StoreQueue.scala 156:23]
        if (deq_req_empty & _T_11) begin // @[StoreQueue.scala 157:45]
          sq_0_valid <= 1'h0; // @[StoreQueue.scala 149:19]
        end else begin
          sq_0_valid <= _GEN_35;
        end
      end else begin
        sq_0_valid <= _GEN_35;
      end
    end else if (flush_state) begin // @[StoreQueue.scala 153:24]
      if (deq_req_empty) begin // @[StoreQueue.scala 172:28]
        sq_0_valid <= 1'h0; // @[StoreQueue.scala 149:19]
      end else begin
        sq_0_valid <= _GEN_35;
      end
    end else begin
      sq_0_valid <= _GEN_35;
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_1_addr <= 32'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h1 == value) begin // @[StoreQueue.scala 105:23]
        sq_1_addr <= io_in_st_req_bits_addr; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_1_wdata <= 64'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h1 == value) begin // @[StoreQueue.scala 105:23]
        sq_1_wdata <= io_in_st_req_bits_wdata; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_1_wmask <= 8'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h1 == value) begin // @[StoreQueue.scala 105:23]
        sq_1_wmask <= io_in_st_req_bits_wmask; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_1_wsize <= 2'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h1 == value) begin // @[StoreQueue.scala 105:23]
        sq_1_wsize <= io_in_st_req_bits_size; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_1_valid <= 1'h0; // @[StoreQueue.scala 31:19]
    end else if (_T_22) begin // @[StoreQueue.scala 153:24]
      if (io_flush) begin // @[StoreQueue.scala 156:23]
        if (deq_req_empty & _T_11) begin // @[StoreQueue.scala 157:45]
          sq_1_valid <= 1'h0; // @[StoreQueue.scala 149:19]
        end else begin
          sq_1_valid <= _GEN_36;
        end
      end else begin
        sq_1_valid <= _GEN_36;
      end
    end else if (flush_state) begin // @[StoreQueue.scala 153:24]
      if (deq_req_empty) begin // @[StoreQueue.scala 172:28]
        sq_1_valid <= 1'h0; // @[StoreQueue.scala 149:19]
      end else begin
        sq_1_valid <= _GEN_36;
      end
    end else begin
      sq_1_valid <= _GEN_36;
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_2_addr <= 32'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h2 == value) begin // @[StoreQueue.scala 105:23]
        sq_2_addr <= io_in_st_req_bits_addr; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_2_wdata <= 64'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h2 == value) begin // @[StoreQueue.scala 105:23]
        sq_2_wdata <= io_in_st_req_bits_wdata; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_2_wmask <= 8'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h2 == value) begin // @[StoreQueue.scala 105:23]
        sq_2_wmask <= io_in_st_req_bits_wmask; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_2_wsize <= 2'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h2 == value) begin // @[StoreQueue.scala 105:23]
        sq_2_wsize <= io_in_st_req_bits_size; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_2_valid <= 1'h0; // @[StoreQueue.scala 31:19]
    end else if (_T_22) begin // @[StoreQueue.scala 153:24]
      if (io_flush) begin // @[StoreQueue.scala 156:23]
        if (deq_req_empty & _T_11) begin // @[StoreQueue.scala 157:45]
          sq_2_valid <= 1'h0; // @[StoreQueue.scala 149:19]
        end else begin
          sq_2_valid <= _GEN_37;
        end
      end else begin
        sq_2_valid <= _GEN_37;
      end
    end else if (flush_state) begin // @[StoreQueue.scala 153:24]
      if (deq_req_empty) begin // @[StoreQueue.scala 172:28]
        sq_2_valid <= 1'h0; // @[StoreQueue.scala 149:19]
      end else begin
        sq_2_valid <= _GEN_37;
      end
    end else begin
      sq_2_valid <= _GEN_37;
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_3_addr <= 32'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h3 == value) begin // @[StoreQueue.scala 105:23]
        sq_3_addr <= io_in_st_req_bits_addr; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_3_wdata <= 64'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h3 == value) begin // @[StoreQueue.scala 105:23]
        sq_3_wdata <= io_in_st_req_bits_wdata; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_3_wmask <= 8'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h3 == value) begin // @[StoreQueue.scala 105:23]
        sq_3_wmask <= io_in_st_req_bits_wmask; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_3_wsize <= 2'h0; // @[StoreQueue.scala 31:19]
    end else if (enq_fire) begin // @[StoreQueue.scala 98:19]
      if (2'h3 == value) begin // @[StoreQueue.scala 105:23]
        sq_3_wsize <= io_in_st_req_bits_size; // @[StoreQueue.scala 105:23]
      end
    end
    if (reset) begin // @[StoreQueue.scala 31:19]
      sq_3_valid <= 1'h0; // @[StoreQueue.scala 31:19]
    end else if (_T_22) begin // @[StoreQueue.scala 153:24]
      if (io_flush) begin // @[StoreQueue.scala 156:23]
        if (deq_req_empty & _T_11) begin // @[StoreQueue.scala 157:45]
          sq_3_valid <= 1'h0; // @[StoreQueue.scala 149:19]
        end else begin
          sq_3_valid <= _GEN_38;
        end
      end else begin
        sq_3_valid <= _GEN_38;
      end
    end else if (flush_state) begin // @[StoreQueue.scala 153:24]
      if (deq_req_empty) begin // @[StoreQueue.scala 172:28]
        sq_3_valid <= 1'h0; // @[StoreQueue.scala 149:19]
      end else begin
        sq_3_valid <= _GEN_38;
      end
    end else begin
      sq_3_valid <= _GEN_38;
    end
    if (reset) begin // @[Counter.scala 60:40]
      value <= 2'h0; // @[Counter.scala 60:40]
    end else if (_T_22) begin // @[StoreQueue.scala 153:24]
      if (io_flush) begin // @[StoreQueue.scala 156:23]
        if (deq_req_empty & _T_11) begin // @[StoreQueue.scala 157:45]
          value <= 2'h0; // @[Counter.scala 97:11]
        end else begin
          value <= _GEN_55;
        end
      end else begin
        value <= _GEN_55;
      end
    end else if (flush_state) begin // @[StoreQueue.scala 153:24]
      if (deq_req_empty) begin // @[StoreQueue.scala 172:28]
        value <= 2'h0; // @[Counter.scala 97:11]
      end else begin
        value <= _GEN_55;
      end
    end else begin
      value <= _GEN_55;
    end
    if (reset) begin // @[Counter.scala 60:40]
      value_1 <= 2'h0; // @[Counter.scala 60:40]
    end else if (_T_22) begin // @[StoreQueue.scala 153:24]
      if (io_flush) begin // @[StoreQueue.scala 156:23]
        if (deq_req_empty & _T_11) begin // @[StoreQueue.scala 157:45]
          value_1 <= 2'h0; // @[Counter.scala 97:11]
        end else begin
          value_1 <= _GEN_10;
        end
      end else begin
        value_1 <= _GEN_10;
      end
    end else if (flush_state) begin // @[StoreQueue.scala 153:24]
      if (deq_req_empty) begin // @[StoreQueue.scala 172:28]
        value_1 <= 2'h0; // @[Counter.scala 97:11]
      end else begin
        value_1 <= _GEN_10;
      end
    end else begin
      value_1 <= _GEN_10;
    end
    if (reset) begin // @[StoreQueue.scala 34:27]
      maybe_full <= 1'h0; // @[StoreQueue.scala 34:27]
    end else if (_T_22) begin // @[StoreQueue.scala 153:24]
      if (io_flush) begin // @[StoreQueue.scala 156:23]
        if (deq_req_empty & _T_11) begin // @[StoreQueue.scala 157:45]
          maybe_full <= 1'h0; // @[StoreQueue.scala 147:16]
        end else begin
          maybe_full <= _GEN_60;
        end
      end else begin
        maybe_full <= _GEN_60;
      end
    end else if (flush_state) begin // @[StoreQueue.scala 153:24]
      if (deq_req_empty) begin // @[StoreQueue.scala 172:28]
        maybe_full <= 1'h0; // @[StoreQueue.scala 147:16]
      end else begin
        maybe_full <= _GEN_60;
      end
    end else begin
      maybe_full <= _GEN_60;
    end
    if (reset) begin // @[StoreQueue.scala 43:26]
      deq_state <= 1'h0; // @[StoreQueue.scala 43:26]
    end else if (_T_5) begin // @[StoreQueue.scala 79:22]
      deq_state <= _GEN_11;
    end else if (deq_state) begin // @[StoreQueue.scala 79:22]
      if (_T_17) begin // @[StoreQueue.scala 86:36]
        deq_state <= 1'h0; // @[StoreQueue.scala 87:19]
      end
    end
    if (reset) begin // @[StoreQueue.scala 46:26]
      enq_state <= 1'h0; // @[StoreQueue.scala 46:26]
    end else if (_T_20) begin // @[StoreQueue.scala 114:22]
      enq_state <= _GEN_56;
    end else if (enq_state) begin // @[StoreQueue.scala 114:22]
      if (_T_25) begin // @[StoreQueue.scala 121:35]
        enq_state <= 1'h0; // @[StoreQueue.scala 122:19]
      end
    end
    if (reset) begin // @[StoreQueue.scala 49:28]
      flush_state <= 1'h0; // @[StoreQueue.scala 49:28]
    end else if (_T_22) begin // @[StoreQueue.scala 153:24]
      if (io_flush) begin // @[StoreQueue.scala 156:23]
        if (!(deq_req_empty & _T_11)) begin // @[StoreQueue.scala 157:45]
          flush_state <= 1'h1; // @[StoreQueue.scala 163:23]
        end
      end
    end else if (flush_state) begin // @[StoreQueue.scala 153:24]
      if (deq_req_empty) begin // @[StoreQueue.scala 172:28]
        flush_state <= 1'h0; // @[StoreQueue.scala 174:21]
      end
    end
    if (reset) begin // @[StoreQueue.scala 55:32]
      deq_req_counter <= 3'h0; // @[StoreQueue.scala 55:32]
    end else if (io_deq_req & ~deq_fire) begin // @[StoreQueue.scala 63:34]
      deq_req_counter <= _T_10; // @[StoreQueue.scala 64:21]
    end else if (~io_deq_req & deq_fire) begin // @[StoreQueue.scala 65:41]
      deq_req_counter <= _T_14; // @[StoreQueue.scala 66:21]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sq_0_addr = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  sq_0_wdata = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  sq_0_wmask = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  sq_0_wsize = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  sq_0_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  sq_1_addr = _RAND_5[31:0];
  _RAND_6 = {2{`RANDOM}};
  sq_1_wdata = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  sq_1_wmask = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  sq_1_wsize = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  sq_1_valid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  sq_2_addr = _RAND_10[31:0];
  _RAND_11 = {2{`RANDOM}};
  sq_2_wdata = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  sq_2_wmask = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  sq_2_wsize = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  sq_2_valid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  sq_3_addr = _RAND_15[31:0];
  _RAND_16 = {2{`RANDOM}};
  sq_3_wdata = _RAND_16[63:0];
  _RAND_17 = {1{`RANDOM}};
  sq_3_wmask = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  sq_3_wsize = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  sq_3_valid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  value = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  value_1 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  maybe_full = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  deq_state = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  enq_state = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  flush_state = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  deq_req_counter = _RAND_26[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_RRArbiter(
  input         clock,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [63:0] io_in_0_bits_wdata,
  input  [7:0]  io_in_0_bits_wmask,
  input  [1:0]  io_in_0_bits_size,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [1:0]  io_in_1_bits_size,
  input         io_out_ready,
  output        io_out_valid,
  output [3:0]  io_out_bits_id,
  output [31:0] io_out_bits_addr,
  output [63:0] io_out_bits_wdata,
  output [7:0]  io_out_bits_wmask,
  output        io_out_bits_wen,
  output [1:0]  io_out_bits_size,
  output        io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _ctrl_validMask_grantMask_lastGrant_T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg  lastGrant; // @[Reg.scala 15:16]
  wire  grantMask_1 = 1'h1 > lastGrant; // @[Arbiter.scala 67:49]
  wire  validMask_1 = io_in_1_valid & grantMask_1; // @[Arbiter.scala 68:75]
  wire  _GEN_15 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:{27,36}]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:{16,16}]
  assign io_out_bits_id = io_chosen ? 4'h2 : 4'h1; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wdata = io_chosen ? 64'h0 : io_in_0_bits_wdata; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wmask = io_chosen ? 8'h0 : io_in_0_bits_wmask; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wen = io_chosen ? 1'h0 : 1'h1; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_size = io_chosen ? io_in_1_bits_size : io_in_0_bits_size; // @[Arbiter.scala 42:{15,15}]
  assign io_chosen = validMask_1 | _GEN_15; // @[Arbiter.scala 79:{25,34}]
  always @(posedge clock) begin
    if (_ctrl_validMask_grantMask_lastGrant_T) begin // @[Reg.scala 16:19]
      lastGrant <= io_chosen; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lastGrant = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_CacheBusCrossbarNto1(
  input         clock,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [31:0] io_in_0_req_bits_addr,
  input  [63:0] io_in_0_req_bits_wdata,
  input  [7:0]  io_in_0_req_bits_wmask,
  input  [1:0]  io_in_0_req_bits_size,
  input         io_in_0_resp_ready,
  output        io_in_0_resp_valid,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [31:0] io_in_1_req_bits_addr,
  input  [1:0]  io_in_1_req_bits_size,
  input         io_in_1_resp_ready,
  output        io_in_1_resp_valid,
  output [63:0] io_in_1_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [3:0]  io_out_req_bits_id,
  output [31:0] io_out_req_bits_addr,
  output [63:0] io_out_req_bits_wdata,
  output [7:0]  io_out_req_bits_wmask,
  output        io_out_req_bits_wen,
  output [1:0]  io_out_req_bits_size,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_id,
  input  [63:0] io_out_resp_bits_rdata
);
  wire  arbiter_clock; // @[Crossbar.scala 49:23]
  wire  arbiter_io_in_0_valid; // @[Crossbar.scala 49:23]
  wire [31:0] arbiter_io_in_0_bits_addr; // @[Crossbar.scala 49:23]
  wire [63:0] arbiter_io_in_0_bits_wdata; // @[Crossbar.scala 49:23]
  wire [7:0] arbiter_io_in_0_bits_wmask; // @[Crossbar.scala 49:23]
  wire [1:0] arbiter_io_in_0_bits_size; // @[Crossbar.scala 49:23]
  wire  arbiter_io_in_1_valid; // @[Crossbar.scala 49:23]
  wire [31:0] arbiter_io_in_1_bits_addr; // @[Crossbar.scala 49:23]
  wire [1:0] arbiter_io_in_1_bits_size; // @[Crossbar.scala 49:23]
  wire  arbiter_io_out_ready; // @[Crossbar.scala 49:23]
  wire  arbiter_io_out_valid; // @[Crossbar.scala 49:23]
  wire [3:0] arbiter_io_out_bits_id; // @[Crossbar.scala 49:23]
  wire [31:0] arbiter_io_out_bits_addr; // @[Crossbar.scala 49:23]
  wire [63:0] arbiter_io_out_bits_wdata; // @[Crossbar.scala 49:23]
  wire [7:0] arbiter_io_out_bits_wmask; // @[Crossbar.scala 49:23]
  wire  arbiter_io_out_bits_wen; // @[Crossbar.scala 49:23]
  wire [1:0] arbiter_io_out_bits_size; // @[Crossbar.scala 49:23]
  wire  arbiter_io_chosen; // @[Crossbar.scala 49:23]
  wire  _GEN_0 = io_out_resp_bits_id == 4'h1 & io_in_0_resp_ready; // @[Crossbar.scala 69:23 72:46 73:25]
  ysyx_210128_RRArbiter arbiter ( // @[Crossbar.scala 49:23]
    .clock(arbiter_clock),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_0_bits_addr(arbiter_io_in_0_bits_addr),
    .io_in_0_bits_wdata(arbiter_io_in_0_bits_wdata),
    .io_in_0_bits_wmask(arbiter_io_in_0_bits_wmask),
    .io_in_0_bits_size(arbiter_io_in_0_bits_size),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_1_bits_addr(arbiter_io_in_1_bits_addr),
    .io_in_1_bits_size(arbiter_io_in_1_bits_size),
    .io_out_ready(arbiter_io_out_ready),
    .io_out_valid(arbiter_io_out_valid),
    .io_out_bits_id(arbiter_io_out_bits_id),
    .io_out_bits_addr(arbiter_io_out_bits_addr),
    .io_out_bits_wdata(arbiter_io_out_bits_wdata),
    .io_out_bits_wmask(arbiter_io_out_bits_wmask),
    .io_out_bits_wen(arbiter_io_out_bits_wen),
    .io_out_bits_size(arbiter_io_out_bits_size),
    .io_chosen(arbiter_io_chosen)
  );
  assign io_in_0_req_ready = ~arbiter_io_chosen & io_out_req_ready; // @[Crossbar.scala 57:55]
  assign io_in_0_resp_valid = io_out_resp_bits_id == 4'h1 & io_out_resp_valid; // @[Crossbar.scala 68:25 72:46 74:27]
  assign io_in_1_req_ready = arbiter_io_chosen & io_out_req_ready; // @[Crossbar.scala 57:55]
  assign io_in_1_resp_valid = io_out_resp_bits_id == 4'h2 & io_out_resp_valid; // @[Crossbar.scala 68:25 72:46 74:27]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 67:24]
  assign io_out_req_valid = arbiter_io_out_valid; // @[Crossbar.scala 61:13]
  assign io_out_req_bits_id = arbiter_io_out_bits_id; // @[Crossbar.scala 60:12]
  assign io_out_req_bits_addr = arbiter_io_out_bits_addr; // @[Crossbar.scala 60:12]
  assign io_out_req_bits_wdata = arbiter_io_out_bits_wdata; // @[Crossbar.scala 60:12]
  assign io_out_req_bits_wmask = arbiter_io_out_bits_wmask; // @[Crossbar.scala 60:12]
  assign io_out_req_bits_wen = arbiter_io_out_bits_wen; // @[Crossbar.scala 60:12]
  assign io_out_req_bits_size = arbiter_io_out_bits_size; // @[Crossbar.scala 60:12]
  assign io_out_resp_ready = io_out_resp_bits_id == 4'h2 ? io_in_1_resp_ready : _GEN_0; // @[Crossbar.scala 72:46 73:25]
  assign arbiter_clock = clock;
  assign arbiter_io_in_0_valid = io_in_0_req_valid; // @[Crossbar.scala 52:22]
  assign arbiter_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Crossbar.scala 52:22]
  assign arbiter_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Crossbar.scala 52:22]
  assign arbiter_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[Crossbar.scala 52:22]
  assign arbiter_io_in_0_bits_size = io_in_0_req_bits_size; // @[Crossbar.scala 52:22]
  assign arbiter_io_in_1_valid = io_in_1_req_valid; // @[Crossbar.scala 52:22]
  assign arbiter_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Crossbar.scala 52:22]
  assign arbiter_io_in_1_bits_size = io_in_1_req_bits_size; // @[Crossbar.scala 52:22]
  assign arbiter_io_out_ready = io_out_req_ready; // @[Crossbar.scala 62:13]
endmodule
module ysyx_210128_CacheBusCrossbar1to2_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [3:0]  io_in_req_bits_id,
  input  [31:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input  [1:0]  io_in_req_bits_size,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_id,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_0_req_ready,
  output        io_out_0_req_valid,
  output [3:0]  io_out_0_req_bits_id,
  output [31:0] io_out_0_req_bits_addr,
  output [63:0] io_out_0_req_bits_wdata,
  output [7:0]  io_out_0_req_bits_wmask,
  output        io_out_0_req_bits_wen,
  output [1:0]  io_out_0_req_bits_size,
  output        io_out_0_resp_ready,
  input         io_out_0_resp_valid,
  input  [3:0]  io_out_0_resp_bits_id,
  input  [63:0] io_out_0_resp_bits_rdata,
  input         io_out_1_req_ready,
  output        io_out_1_req_valid,
  output [3:0]  io_out_1_req_bits_id,
  output [31:0] io_out_1_req_bits_addr,
  output [63:0] io_out_1_req_bits_wdata,
  output [7:0]  io_out_1_req_bits_wmask,
  output        io_out_1_req_bits_wen,
  output [1:0]  io_out_1_req_bits_size,
  output        io_out_1_resp_ready,
  input         io_out_1_resp_valid,
  input  [3:0]  io_out_1_resp_bits_id,
  input  [63:0] io_out_1_resp_bits_rdata,
  input         io_to_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] in_flight_req_0; // @[Crossbar.scala 87:30]
  reg [7:0] in_flight_req_1; // @[Crossbar.scala 87:30]
  wire  _T = io_out_0_req_ready & io_out_0_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_1 = io_out_0_resp_ready & io_out_0_resp_valid; // @[Decoupled.scala 40:37]
  wire [7:0] _T_5 = in_flight_req_0 + 8'h1; // @[Crossbar.scala 90:44]
  wire [7:0] _T_11 = in_flight_req_0 - 8'h1; // @[Crossbar.scala 95:44]
  wire  _T_12 = io_out_1_req_ready & io_out_1_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_13 = io_out_1_resp_ready & io_out_1_resp_valid; // @[Decoupled.scala 40:37]
  wire [7:0] _T_17 = in_flight_req_1 + 8'h1; // @[Crossbar.scala 90:44]
  wire [7:0] _T_23 = in_flight_req_1 - 8'h1; // @[Crossbar.scala 95:44]
  wire  req_0_ready = in_flight_req_1 == 8'h0; // @[Crossbar.scala 102:39]
  wire  req_1_ready = in_flight_req_0 == 8'h0; // @[Crossbar.scala 103:39]
  reg  channel; // @[Crossbar.scala 105:24]
  wire  _GEN_4 = _T ? 1'h0 : channel; // @[Crossbar.scala 107:33 108:15 105:24]
  wire  _GEN_5 = _T_12 | _GEN_4; // @[Crossbar.scala 107:33 108:15]
  wire  _T_34 = ~channel; // @[Crossbar.scala 120:57]
  wire [63:0] _GEN_6 = _T_34 ? io_out_0_resp_bits_rdata : 64'h0; // @[Crossbar.scala 130:28 131:23 127:25]
  wire [3:0] _GEN_7 = _T_34 ? io_out_0_resp_bits_id : 4'h0; // @[Crossbar.scala 130:28 131:23 122:25]
  wire  _GEN_8 = _T_34 & io_out_0_resp_valid; // @[Crossbar.scala 130:28 132:24 128:25]
  assign io_in_req_ready = io_to_1 ? io_out_1_req_ready & req_1_ready : io_out_0_req_ready & req_0_ready; // @[Crossbar.scala 117:29]
  assign io_in_resp_valid = channel ? io_out_1_resp_valid : _GEN_8; // @[Crossbar.scala 130:28 132:24]
  assign io_in_resp_bits_id = channel ? io_out_1_resp_bits_id : _GEN_7; // @[Crossbar.scala 130:28 131:23]
  assign io_in_resp_bits_rdata = channel ? io_out_1_resp_bits_rdata : _GEN_6; // @[Crossbar.scala 130:28 131:23]
  assign io_out_0_req_valid = io_in_req_valid & ~io_to_1 & req_0_ready; // @[Crossbar.scala 115:54]
  assign io_out_0_req_bits_id = io_in_req_bits_id; // @[Crossbar.scala 113:23]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 113:23]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 113:23]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 113:23]
  assign io_out_0_req_bits_wen = io_in_req_bits_wen; // @[Crossbar.scala 113:23]
  assign io_out_0_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 113:23]
  assign io_out_0_resp_ready = io_in_resp_ready & ~channel; // @[Crossbar.scala 120:45]
  assign io_out_1_req_valid = io_in_req_valid & io_to_1 & req_1_ready; // @[Crossbar.scala 116:53]
  assign io_out_1_req_bits_id = io_in_req_bits_id; // @[Crossbar.scala 114:23]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 114:23]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 114:23]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 114:23]
  assign io_out_1_req_bits_wen = io_in_req_bits_wen; // @[Crossbar.scala 114:23]
  assign io_out_1_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 114:23]
  assign io_out_1_resp_ready = io_in_resp_ready & channel; // @[Crossbar.scala 121:45]
  always @(posedge clock) begin
    if (reset) begin // @[Crossbar.scala 87:30]
      in_flight_req_0 <= 8'h0; // @[Crossbar.scala 87:30]
    end else if (_T & ~_T_1) begin // @[Crossbar.scala 89:59]
      in_flight_req_0 <= _T_5; // @[Crossbar.scala 90:24]
    end else if (_T_1 & ~_T) begin // @[Crossbar.scala 94:66]
      in_flight_req_0 <= _T_11; // @[Crossbar.scala 95:24]
    end
    if (reset) begin // @[Crossbar.scala 87:30]
      in_flight_req_1 <= 8'h0; // @[Crossbar.scala 87:30]
    end else if (_T_12 & ~_T_13) begin // @[Crossbar.scala 89:59]
      in_flight_req_1 <= _T_17; // @[Crossbar.scala 90:24]
    end else if (_T_13 & ~_T_12) begin // @[Crossbar.scala 94:66]
      in_flight_req_1 <= _T_23; // @[Crossbar.scala 95:24]
    end
    if (reset) begin // @[Crossbar.scala 105:24]
      channel <= 1'h0; // @[Crossbar.scala 105:24]
    end else begin
      channel <= _GEN_5;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_flight_req_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  in_flight_req_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  channel = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_Cache_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [3:0]  io_in_req_bits_id,
  input  [31:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_id,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output        io_out_req_bits_aen,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_req_bits_wlast,
  output        io_out_req_bits_wen,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_out_resp_bits_rlast,
  input         fence_i_0,
  output        _WIRE_10_0,
  input         sq_empty_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [127:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [127:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [127:0] _RAND_222;
  reg [31:0] _RAND_223;
`endif // RANDOMIZE_REG_INIT
  wire  sram_0_clock; // @[Cache.scala 89:22]
  wire  sram_0_io_en; // @[Cache.scala 89:22]
  wire  sram_0_io_wen; // @[Cache.scala 89:22]
  wire [5:0] sram_0_io_addr; // @[Cache.scala 89:22]
  wire [127:0] sram_0_io_wdata; // @[Cache.scala 89:22]
  wire [127:0] sram_0_io_rdata; // @[Cache.scala 89:22]
  wire  sram_1_clock; // @[Cache.scala 89:22]
  wire  sram_1_io_en; // @[Cache.scala 89:22]
  wire  sram_1_io_wen; // @[Cache.scala 89:22]
  wire [5:0] sram_1_io_addr; // @[Cache.scala 89:22]
  wire [127:0] sram_1_io_wdata; // @[Cache.scala 89:22]
  wire [127:0] sram_1_io_rdata; // @[Cache.scala 89:22]
  wire  sram_2_clock; // @[Cache.scala 89:22]
  wire  sram_2_io_en; // @[Cache.scala 89:22]
  wire  sram_2_io_wen; // @[Cache.scala 89:22]
  wire [5:0] sram_2_io_addr; // @[Cache.scala 89:22]
  wire [127:0] sram_2_io_wdata; // @[Cache.scala 89:22]
  wire [127:0] sram_2_io_rdata; // @[Cache.scala 89:22]
  wire  sram_3_clock; // @[Cache.scala 89:22]
  wire  sram_3_io_en; // @[Cache.scala 89:22]
  wire  sram_3_io_wen; // @[Cache.scala 89:22]
  wire [5:0] sram_3_io_addr; // @[Cache.scala 89:22]
  wire [127:0] sram_3_io_wdata; // @[Cache.scala 89:22]
  wire [127:0] sram_3_io_rdata; // @[Cache.scala 89:22]
  wire  meta_0_clock; // @[Cache.scala 97:22]
  wire  meta_0_reset; // @[Cache.scala 97:22]
  wire [5:0] meta_0_io_idx; // @[Cache.scala 97:22]
  wire [20:0] meta_0_io_tag_r; // @[Cache.scala 97:22]
  wire [20:0] meta_0_io_tag_w; // @[Cache.scala 97:22]
  wire  meta_0_io_tag_wen; // @[Cache.scala 97:22]
  wire  meta_0_io_dirty_r_async; // @[Cache.scala 97:22]
  wire  meta_0_io_dirty_w; // @[Cache.scala 97:22]
  wire  meta_0_io_dirty_wen; // @[Cache.scala 97:22]
  wire  meta_0_io_valid_r_async; // @[Cache.scala 97:22]
  wire  meta_0_io_invalidate; // @[Cache.scala 97:22]
  wire  meta_1_clock; // @[Cache.scala 97:22]
  wire  meta_1_reset; // @[Cache.scala 97:22]
  wire [5:0] meta_1_io_idx; // @[Cache.scala 97:22]
  wire [20:0] meta_1_io_tag_r; // @[Cache.scala 97:22]
  wire [20:0] meta_1_io_tag_w; // @[Cache.scala 97:22]
  wire  meta_1_io_tag_wen; // @[Cache.scala 97:22]
  wire  meta_1_io_dirty_r_async; // @[Cache.scala 97:22]
  wire  meta_1_io_dirty_w; // @[Cache.scala 97:22]
  wire  meta_1_io_dirty_wen; // @[Cache.scala 97:22]
  wire  meta_1_io_valid_r_async; // @[Cache.scala 97:22]
  wire  meta_1_io_invalidate; // @[Cache.scala 97:22]
  wire  meta_2_clock; // @[Cache.scala 97:22]
  wire  meta_2_reset; // @[Cache.scala 97:22]
  wire [5:0] meta_2_io_idx; // @[Cache.scala 97:22]
  wire [20:0] meta_2_io_tag_r; // @[Cache.scala 97:22]
  wire [20:0] meta_2_io_tag_w; // @[Cache.scala 97:22]
  wire  meta_2_io_tag_wen; // @[Cache.scala 97:22]
  wire  meta_2_io_dirty_r_async; // @[Cache.scala 97:22]
  wire  meta_2_io_dirty_w; // @[Cache.scala 97:22]
  wire  meta_2_io_dirty_wen; // @[Cache.scala 97:22]
  wire  meta_2_io_valid_r_async; // @[Cache.scala 97:22]
  wire  meta_2_io_invalidate; // @[Cache.scala 97:22]
  wire  meta_3_clock; // @[Cache.scala 97:22]
  wire  meta_3_reset; // @[Cache.scala 97:22]
  wire [5:0] meta_3_io_idx; // @[Cache.scala 97:22]
  wire [20:0] meta_3_io_tag_r; // @[Cache.scala 97:22]
  wire [20:0] meta_3_io_tag_w; // @[Cache.scala 97:22]
  wire  meta_3_io_tag_wen; // @[Cache.scala 97:22]
  wire  meta_3_io_dirty_r_async; // @[Cache.scala 97:22]
  wire  meta_3_io_dirty_w; // @[Cache.scala 97:22]
  wire  meta_3_io_dirty_wen; // @[Cache.scala 97:22]
  wire  meta_3_io_valid_r_async; // @[Cache.scala 97:22]
  wire  meta_3_io_invalidate; // @[Cache.scala 97:22]
  reg  REG; // @[Cache.scala 123:59]
  reg  REG_1; // @[Cache.scala 123:59]
  reg  REG_2; // @[Cache.scala 123:59]
  reg  REG_3; // @[Cache.scala 123:59]
  reg  REG_4; // @[Cache.scala 124:59]
  reg  REG_5; // @[Cache.scala 124:59]
  reg  REG_6; // @[Cache.scala 124:59]
  reg  REG_7; // @[Cache.scala 124:59]
  reg  plru0_0; // @[Cache.scala 129:22]
  reg  plru0_1; // @[Cache.scala 129:22]
  reg  plru0_2; // @[Cache.scala 129:22]
  reg  plru0_3; // @[Cache.scala 129:22]
  reg  plru0_4; // @[Cache.scala 129:22]
  reg  plru0_5; // @[Cache.scala 129:22]
  reg  plru0_6; // @[Cache.scala 129:22]
  reg  plru0_7; // @[Cache.scala 129:22]
  reg  plru0_8; // @[Cache.scala 129:22]
  reg  plru0_9; // @[Cache.scala 129:22]
  reg  plru0_10; // @[Cache.scala 129:22]
  reg  plru0_11; // @[Cache.scala 129:22]
  reg  plru0_12; // @[Cache.scala 129:22]
  reg  plru0_13; // @[Cache.scala 129:22]
  reg  plru0_14; // @[Cache.scala 129:22]
  reg  plru0_15; // @[Cache.scala 129:22]
  reg  plru0_16; // @[Cache.scala 129:22]
  reg  plru0_17; // @[Cache.scala 129:22]
  reg  plru0_18; // @[Cache.scala 129:22]
  reg  plru0_19; // @[Cache.scala 129:22]
  reg  plru0_20; // @[Cache.scala 129:22]
  reg  plru0_21; // @[Cache.scala 129:22]
  reg  plru0_22; // @[Cache.scala 129:22]
  reg  plru0_23; // @[Cache.scala 129:22]
  reg  plru0_24; // @[Cache.scala 129:22]
  reg  plru0_25; // @[Cache.scala 129:22]
  reg  plru0_26; // @[Cache.scala 129:22]
  reg  plru0_27; // @[Cache.scala 129:22]
  reg  plru0_28; // @[Cache.scala 129:22]
  reg  plru0_29; // @[Cache.scala 129:22]
  reg  plru0_30; // @[Cache.scala 129:22]
  reg  plru0_31; // @[Cache.scala 129:22]
  reg  plru0_32; // @[Cache.scala 129:22]
  reg  plru0_33; // @[Cache.scala 129:22]
  reg  plru0_34; // @[Cache.scala 129:22]
  reg  plru0_35; // @[Cache.scala 129:22]
  reg  plru0_36; // @[Cache.scala 129:22]
  reg  plru0_37; // @[Cache.scala 129:22]
  reg  plru0_38; // @[Cache.scala 129:22]
  reg  plru0_39; // @[Cache.scala 129:22]
  reg  plru0_40; // @[Cache.scala 129:22]
  reg  plru0_41; // @[Cache.scala 129:22]
  reg  plru0_42; // @[Cache.scala 129:22]
  reg  plru0_43; // @[Cache.scala 129:22]
  reg  plru0_44; // @[Cache.scala 129:22]
  reg  plru0_45; // @[Cache.scala 129:22]
  reg  plru0_46; // @[Cache.scala 129:22]
  reg  plru0_47; // @[Cache.scala 129:22]
  reg  plru0_48; // @[Cache.scala 129:22]
  reg  plru0_49; // @[Cache.scala 129:22]
  reg  plru0_50; // @[Cache.scala 129:22]
  reg  plru0_51; // @[Cache.scala 129:22]
  reg  plru0_52; // @[Cache.scala 129:22]
  reg  plru0_53; // @[Cache.scala 129:22]
  reg  plru0_54; // @[Cache.scala 129:22]
  reg  plru0_55; // @[Cache.scala 129:22]
  reg  plru0_56; // @[Cache.scala 129:22]
  reg  plru0_57; // @[Cache.scala 129:22]
  reg  plru0_58; // @[Cache.scala 129:22]
  reg  plru0_59; // @[Cache.scala 129:22]
  reg  plru0_60; // @[Cache.scala 129:22]
  reg  plru0_61; // @[Cache.scala 129:22]
  reg  plru0_62; // @[Cache.scala 129:22]
  reg  plru0_63; // @[Cache.scala 129:22]
  reg  plru1_0; // @[Cache.scala 131:22]
  reg  plru1_1; // @[Cache.scala 131:22]
  reg  plru1_2; // @[Cache.scala 131:22]
  reg  plru1_3; // @[Cache.scala 131:22]
  reg  plru1_4; // @[Cache.scala 131:22]
  reg  plru1_5; // @[Cache.scala 131:22]
  reg  plru1_6; // @[Cache.scala 131:22]
  reg  plru1_7; // @[Cache.scala 131:22]
  reg  plru1_8; // @[Cache.scala 131:22]
  reg  plru1_9; // @[Cache.scala 131:22]
  reg  plru1_10; // @[Cache.scala 131:22]
  reg  plru1_11; // @[Cache.scala 131:22]
  reg  plru1_12; // @[Cache.scala 131:22]
  reg  plru1_13; // @[Cache.scala 131:22]
  reg  plru1_14; // @[Cache.scala 131:22]
  reg  plru1_15; // @[Cache.scala 131:22]
  reg  plru1_16; // @[Cache.scala 131:22]
  reg  plru1_17; // @[Cache.scala 131:22]
  reg  plru1_18; // @[Cache.scala 131:22]
  reg  plru1_19; // @[Cache.scala 131:22]
  reg  plru1_20; // @[Cache.scala 131:22]
  reg  plru1_21; // @[Cache.scala 131:22]
  reg  plru1_22; // @[Cache.scala 131:22]
  reg  plru1_23; // @[Cache.scala 131:22]
  reg  plru1_24; // @[Cache.scala 131:22]
  reg  plru1_25; // @[Cache.scala 131:22]
  reg  plru1_26; // @[Cache.scala 131:22]
  reg  plru1_27; // @[Cache.scala 131:22]
  reg  plru1_28; // @[Cache.scala 131:22]
  reg  plru1_29; // @[Cache.scala 131:22]
  reg  plru1_30; // @[Cache.scala 131:22]
  reg  plru1_31; // @[Cache.scala 131:22]
  reg  plru1_32; // @[Cache.scala 131:22]
  reg  plru1_33; // @[Cache.scala 131:22]
  reg  plru1_34; // @[Cache.scala 131:22]
  reg  plru1_35; // @[Cache.scala 131:22]
  reg  plru1_36; // @[Cache.scala 131:22]
  reg  plru1_37; // @[Cache.scala 131:22]
  reg  plru1_38; // @[Cache.scala 131:22]
  reg  plru1_39; // @[Cache.scala 131:22]
  reg  plru1_40; // @[Cache.scala 131:22]
  reg  plru1_41; // @[Cache.scala 131:22]
  reg  plru1_42; // @[Cache.scala 131:22]
  reg  plru1_43; // @[Cache.scala 131:22]
  reg  plru1_44; // @[Cache.scala 131:22]
  reg  plru1_45; // @[Cache.scala 131:22]
  reg  plru1_46; // @[Cache.scala 131:22]
  reg  plru1_47; // @[Cache.scala 131:22]
  reg  plru1_48; // @[Cache.scala 131:22]
  reg  plru1_49; // @[Cache.scala 131:22]
  reg  plru1_50; // @[Cache.scala 131:22]
  reg  plru1_51; // @[Cache.scala 131:22]
  reg  plru1_52; // @[Cache.scala 131:22]
  reg  plru1_53; // @[Cache.scala 131:22]
  reg  plru1_54; // @[Cache.scala 131:22]
  reg  plru1_55; // @[Cache.scala 131:22]
  reg  plru1_56; // @[Cache.scala 131:22]
  reg  plru1_57; // @[Cache.scala 131:22]
  reg  plru1_58; // @[Cache.scala 131:22]
  reg  plru1_59; // @[Cache.scala 131:22]
  reg  plru1_60; // @[Cache.scala 131:22]
  reg  plru1_61; // @[Cache.scala 131:22]
  reg  plru1_62; // @[Cache.scala 131:22]
  reg  plru1_63; // @[Cache.scala 131:22]
  reg  plru2_0; // @[Cache.scala 133:22]
  reg  plru2_1; // @[Cache.scala 133:22]
  reg  plru2_2; // @[Cache.scala 133:22]
  reg  plru2_3; // @[Cache.scala 133:22]
  reg  plru2_4; // @[Cache.scala 133:22]
  reg  plru2_5; // @[Cache.scala 133:22]
  reg  plru2_6; // @[Cache.scala 133:22]
  reg  plru2_7; // @[Cache.scala 133:22]
  reg  plru2_8; // @[Cache.scala 133:22]
  reg  plru2_9; // @[Cache.scala 133:22]
  reg  plru2_10; // @[Cache.scala 133:22]
  reg  plru2_11; // @[Cache.scala 133:22]
  reg  plru2_12; // @[Cache.scala 133:22]
  reg  plru2_13; // @[Cache.scala 133:22]
  reg  plru2_14; // @[Cache.scala 133:22]
  reg  plru2_15; // @[Cache.scala 133:22]
  reg  plru2_16; // @[Cache.scala 133:22]
  reg  plru2_17; // @[Cache.scala 133:22]
  reg  plru2_18; // @[Cache.scala 133:22]
  reg  plru2_19; // @[Cache.scala 133:22]
  reg  plru2_20; // @[Cache.scala 133:22]
  reg  plru2_21; // @[Cache.scala 133:22]
  reg  plru2_22; // @[Cache.scala 133:22]
  reg  plru2_23; // @[Cache.scala 133:22]
  reg  plru2_24; // @[Cache.scala 133:22]
  reg  plru2_25; // @[Cache.scala 133:22]
  reg  plru2_26; // @[Cache.scala 133:22]
  reg  plru2_27; // @[Cache.scala 133:22]
  reg  plru2_28; // @[Cache.scala 133:22]
  reg  plru2_29; // @[Cache.scala 133:22]
  reg  plru2_30; // @[Cache.scala 133:22]
  reg  plru2_31; // @[Cache.scala 133:22]
  reg  plru2_32; // @[Cache.scala 133:22]
  reg  plru2_33; // @[Cache.scala 133:22]
  reg  plru2_34; // @[Cache.scala 133:22]
  reg  plru2_35; // @[Cache.scala 133:22]
  reg  plru2_36; // @[Cache.scala 133:22]
  reg  plru2_37; // @[Cache.scala 133:22]
  reg  plru2_38; // @[Cache.scala 133:22]
  reg  plru2_39; // @[Cache.scala 133:22]
  reg  plru2_40; // @[Cache.scala 133:22]
  reg  plru2_41; // @[Cache.scala 133:22]
  reg  plru2_42; // @[Cache.scala 133:22]
  reg  plru2_43; // @[Cache.scala 133:22]
  reg  plru2_44; // @[Cache.scala 133:22]
  reg  plru2_45; // @[Cache.scala 133:22]
  reg  plru2_46; // @[Cache.scala 133:22]
  reg  plru2_47; // @[Cache.scala 133:22]
  reg  plru2_48; // @[Cache.scala 133:22]
  reg  plru2_49; // @[Cache.scala 133:22]
  reg  plru2_50; // @[Cache.scala 133:22]
  reg  plru2_51; // @[Cache.scala 133:22]
  reg  plru2_52; // @[Cache.scala 133:22]
  reg  plru2_53; // @[Cache.scala 133:22]
  reg  plru2_54; // @[Cache.scala 133:22]
  reg  plru2_55; // @[Cache.scala 133:22]
  reg  plru2_56; // @[Cache.scala 133:22]
  reg  plru2_57; // @[Cache.scala 133:22]
  reg  plru2_58; // @[Cache.scala 133:22]
  reg  plru2_59; // @[Cache.scala 133:22]
  reg  plru2_60; // @[Cache.scala 133:22]
  reg  plru2_61; // @[Cache.scala 133:22]
  reg  plru2_62; // @[Cache.scala 133:22]
  reg  plru2_63; // @[Cache.scala 133:22]
  reg  REG_9; // @[Cache.scala 275:32]
  wire [20:0] tag_out_0 = meta_0_io_tag_r;
  reg [31:0] s2_addr; // @[Cache.scala 215:25]
  wire [20:0] s2_tag = s2_addr[30:10]; // @[Cache.scala 218:25]
  wire  hit_0 = tag_out_0 == s2_tag & REG; // @[Cache.scala 230:25]
  wire [20:0] tag_out_1 = meta_1_io_tag_r;
  wire  hit_1 = tag_out_1 == s2_tag & REG_1; // @[Cache.scala 230:25]
  wire [20:0] tag_out_2 = meta_2_io_tag_r;
  wire  hit_2 = tag_out_2 == s2_tag & REG_2; // @[Cache.scala 230:25]
  wire [20:0] tag_out_3 = meta_3_io_tag_r;
  wire  hit_3 = tag_out_3 == s2_tag & REG_3; // @[Cache.scala 230:25]
  wire [3:0] _T_8 = {hit_0,hit_1,hit_2,hit_3}; // @[Cat.scala 30:58]
  wire  s2_hit = |_T_8; // @[Cache.scala 232:25]
  reg  s2_reg_hit; // @[Cache.scala 239:27]
  wire  s2_hit_real = REG_9 ? s2_hit : s2_reg_hit; // @[Cache.scala 275:24]
  reg  s2_wen; // @[Cache.scala 219:25]
  reg [3:0] state; // @[Cache.scala 213:22]
  wire  _T_18 = state == 4'h7; // @[Cache.scala 277:37]
  wire  _T_20 = s2_wen ? state == 4'h7 : state == 4'h0; // @[Cache.scala 277:22]
  wire  hit_ready = s2_hit_real & _T_20; // @[Cache.scala 276:31]
  wire  invalid_ready = state == 4'h8; // @[Cache.scala 279:30]
  wire  pipeline_ready = (hit_ready | _T_18) & io_in_resp_ready | invalid_ready; // @[Cache.scala 282:66]
  reg  fi_valid; // @[Utils.scala 34:20]
  wire  _GEN_0 = fence_i_0 | fi_valid; // @[Utils.scala 34:20 40:{20,24}]
  reg [2:0] fi_state; // @[Cache.scala 435:25]
  wire  _GEN_3564 = 3'h4 == fi_state ? 1'h0 : 3'h5 == fi_state; // @[Cache.scala 483:23]
  wire  _GEN_3567 = 3'h3 == fi_state ? 1'h0 : _GEN_3564; // @[Cache.scala 483:23]
  wire  _GEN_3570 = 3'h2 == fi_state ? 1'h0 : _GEN_3567; // @[Cache.scala 483:23]
  wire  _GEN_3577 = 3'h1 == fi_state ? 1'h0 : _GEN_3570; // @[Cache.scala 483:23]
  wire  fi_finish = 3'h0 == fi_state ? 1'h0 : _GEN_3577; // @[Cache.scala 483:23]
//   wire  _WIRE_10 = fi_finish; // @[Cache.scala 483:23]
  wire  fi_ready = pipeline_ready & sq_empty_0; // @[Cache.scala 163:33]
  wire  fi_fire = fi_valid & fi_ready; // @[Cache.scala 164:26]
  wire [5:0] s1_idx = io_in_req_bits_addr[9:4]; // @[Cache.scala 170:25]
  wire [5:0] _GEN_3 = pipeline_ready ? s1_idx : 6'h0; // @[Cache.scala 109:15 187:24 190:17]
  wire  s2_offs = s2_addr[3]; // @[Cache.scala 216:25]
  wire [5:0] s2_idx = s2_addr[9:4]; // @[Cache.scala 217:25]
  reg [63:0] s2_wdata; // @[Cache.scala 220:25]
  reg [7:0] s2_wmask; // @[Cache.scala 221:25]
  reg [3:0] s2_id; // @[Cache.scala 223:25]
  wire [3:0] _T_9 = {hit_3,hit_2,hit_1,hit_0}; // @[OneHot.scala 22:45]
  wire [1:0] hi_2 = _T_9[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] lo_2 = _T_9[1:0]; // @[OneHot.scala 31:18]
  wire  _T_10 = |hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _T_11 = hi_2 | lo_2; // @[OneHot.scala 32:28]
  wire [1:0] s2_way = {_T_10,_T_11[1]}; // @[Cat.scala 30:58]
  reg [127:0] s2_reg_rdata; // @[Cache.scala 241:29]
  reg  s2_reg_dirty; // @[Cache.scala 242:29]
  reg [20:0] s2_reg_tag_r; // @[Cache.scala 243:29]
  reg [127:0] s2_reg_dat_w; // @[Cache.scala 244:29]
  reg  REG_8; // @[Cache.scala 256:41]
  wire [127:0] sram_out_0 = sram_0_io_rdata;
  wire [127:0] sram_out_1 = sram_1_io_rdata;
  wire [127:0] _GEN_5 = 2'h1 == s2_way ? sram_out_1 : sram_out_0; // @[Cache.scala 261:{18,18}]
  wire [127:0] sram_out_2 = sram_2_io_rdata;
  wire [127:0] _GEN_6 = 2'h2 == s2_way ? sram_out_2 : _GEN_5; // @[Cache.scala 261:{18,18}]
  wire [127:0] sram_out_3 = sram_3_io_rdata;
  wire [127:0] _GEN_7 = 2'h3 == s2_way ? sram_out_3 : _GEN_6; // @[Cache.scala 261:{18,18}]
  wire  _GEN_38 = 6'h1 == s2_idx ? plru0_1 : plru0_0; // @[Cache.scala 268:{40,40}]
  wire  _GEN_39 = 6'h2 == s2_idx ? plru0_2 : _GEN_38; // @[Cache.scala 268:{40,40}]
  wire  _GEN_40 = 6'h3 == s2_idx ? plru0_3 : _GEN_39; // @[Cache.scala 268:{40,40}]
  wire  _GEN_41 = 6'h4 == s2_idx ? plru0_4 : _GEN_40; // @[Cache.scala 268:{40,40}]
  wire  _GEN_42 = 6'h5 == s2_idx ? plru0_5 : _GEN_41; // @[Cache.scala 268:{40,40}]
  wire  _GEN_43 = 6'h6 == s2_idx ? plru0_6 : _GEN_42; // @[Cache.scala 268:{40,40}]
  wire  _GEN_44 = 6'h7 == s2_idx ? plru0_7 : _GEN_43; // @[Cache.scala 268:{40,40}]
  wire  _GEN_45 = 6'h8 == s2_idx ? plru0_8 : _GEN_44; // @[Cache.scala 268:{40,40}]
  wire  _GEN_46 = 6'h9 == s2_idx ? plru0_9 : _GEN_45; // @[Cache.scala 268:{40,40}]
  wire  _GEN_47 = 6'ha == s2_idx ? plru0_10 : _GEN_46; // @[Cache.scala 268:{40,40}]
  wire  _GEN_48 = 6'hb == s2_idx ? plru0_11 : _GEN_47; // @[Cache.scala 268:{40,40}]
  wire  _GEN_49 = 6'hc == s2_idx ? plru0_12 : _GEN_48; // @[Cache.scala 268:{40,40}]
  wire  _GEN_50 = 6'hd == s2_idx ? plru0_13 : _GEN_49; // @[Cache.scala 268:{40,40}]
  wire  _GEN_51 = 6'he == s2_idx ? plru0_14 : _GEN_50; // @[Cache.scala 268:{40,40}]
  wire  _GEN_52 = 6'hf == s2_idx ? plru0_15 : _GEN_51; // @[Cache.scala 268:{40,40}]
  wire  _GEN_53 = 6'h10 == s2_idx ? plru0_16 : _GEN_52; // @[Cache.scala 268:{40,40}]
  wire  _GEN_54 = 6'h11 == s2_idx ? plru0_17 : _GEN_53; // @[Cache.scala 268:{40,40}]
  wire  _GEN_55 = 6'h12 == s2_idx ? plru0_18 : _GEN_54; // @[Cache.scala 268:{40,40}]
  wire  _GEN_56 = 6'h13 == s2_idx ? plru0_19 : _GEN_55; // @[Cache.scala 268:{40,40}]
  wire  _GEN_57 = 6'h14 == s2_idx ? plru0_20 : _GEN_56; // @[Cache.scala 268:{40,40}]
  wire  _GEN_58 = 6'h15 == s2_idx ? plru0_21 : _GEN_57; // @[Cache.scala 268:{40,40}]
  wire  _GEN_59 = 6'h16 == s2_idx ? plru0_22 : _GEN_58; // @[Cache.scala 268:{40,40}]
  wire  _GEN_60 = 6'h17 == s2_idx ? plru0_23 : _GEN_59; // @[Cache.scala 268:{40,40}]
  wire  _GEN_61 = 6'h18 == s2_idx ? plru0_24 : _GEN_60; // @[Cache.scala 268:{40,40}]
  wire  _GEN_62 = 6'h19 == s2_idx ? plru0_25 : _GEN_61; // @[Cache.scala 268:{40,40}]
  wire  _GEN_63 = 6'h1a == s2_idx ? plru0_26 : _GEN_62; // @[Cache.scala 268:{40,40}]
  wire  _GEN_64 = 6'h1b == s2_idx ? plru0_27 : _GEN_63; // @[Cache.scala 268:{40,40}]
  wire  _GEN_65 = 6'h1c == s2_idx ? plru0_28 : _GEN_64; // @[Cache.scala 268:{40,40}]
  wire  _GEN_66 = 6'h1d == s2_idx ? plru0_29 : _GEN_65; // @[Cache.scala 268:{40,40}]
  wire  _GEN_67 = 6'h1e == s2_idx ? plru0_30 : _GEN_66; // @[Cache.scala 268:{40,40}]
  wire  _GEN_68 = 6'h1f == s2_idx ? plru0_31 : _GEN_67; // @[Cache.scala 268:{40,40}]
  wire  _GEN_69 = 6'h20 == s2_idx ? plru0_32 : _GEN_68; // @[Cache.scala 268:{40,40}]
  wire  _GEN_70 = 6'h21 == s2_idx ? plru0_33 : _GEN_69; // @[Cache.scala 268:{40,40}]
  wire  _GEN_71 = 6'h22 == s2_idx ? plru0_34 : _GEN_70; // @[Cache.scala 268:{40,40}]
  wire  _GEN_72 = 6'h23 == s2_idx ? plru0_35 : _GEN_71; // @[Cache.scala 268:{40,40}]
  wire  _GEN_73 = 6'h24 == s2_idx ? plru0_36 : _GEN_72; // @[Cache.scala 268:{40,40}]
  wire  _GEN_74 = 6'h25 == s2_idx ? plru0_37 : _GEN_73; // @[Cache.scala 268:{40,40}]
  wire  _GEN_75 = 6'h26 == s2_idx ? plru0_38 : _GEN_74; // @[Cache.scala 268:{40,40}]
  wire  _GEN_76 = 6'h27 == s2_idx ? plru0_39 : _GEN_75; // @[Cache.scala 268:{40,40}]
  wire  _GEN_77 = 6'h28 == s2_idx ? plru0_40 : _GEN_76; // @[Cache.scala 268:{40,40}]
  wire  _GEN_78 = 6'h29 == s2_idx ? plru0_41 : _GEN_77; // @[Cache.scala 268:{40,40}]
  wire  _GEN_79 = 6'h2a == s2_idx ? plru0_42 : _GEN_78; // @[Cache.scala 268:{40,40}]
  wire  _GEN_80 = 6'h2b == s2_idx ? plru0_43 : _GEN_79; // @[Cache.scala 268:{40,40}]
  wire  _GEN_81 = 6'h2c == s2_idx ? plru0_44 : _GEN_80; // @[Cache.scala 268:{40,40}]
  wire  _GEN_82 = 6'h2d == s2_idx ? plru0_45 : _GEN_81; // @[Cache.scala 268:{40,40}]
  wire  _GEN_83 = 6'h2e == s2_idx ? plru0_46 : _GEN_82; // @[Cache.scala 268:{40,40}]
  wire  _GEN_84 = 6'h2f == s2_idx ? plru0_47 : _GEN_83; // @[Cache.scala 268:{40,40}]
  wire  _GEN_85 = 6'h30 == s2_idx ? plru0_48 : _GEN_84; // @[Cache.scala 268:{40,40}]
  wire  _GEN_86 = 6'h31 == s2_idx ? plru0_49 : _GEN_85; // @[Cache.scala 268:{40,40}]
  wire  _GEN_87 = 6'h32 == s2_idx ? plru0_50 : _GEN_86; // @[Cache.scala 268:{40,40}]
  wire  _GEN_88 = 6'h33 == s2_idx ? plru0_51 : _GEN_87; // @[Cache.scala 268:{40,40}]
  wire  _GEN_89 = 6'h34 == s2_idx ? plru0_52 : _GEN_88; // @[Cache.scala 268:{40,40}]
  wire  _GEN_90 = 6'h35 == s2_idx ? plru0_53 : _GEN_89; // @[Cache.scala 268:{40,40}]
  wire  _GEN_91 = 6'h36 == s2_idx ? plru0_54 : _GEN_90; // @[Cache.scala 268:{40,40}]
  wire  _GEN_92 = 6'h37 == s2_idx ? plru0_55 : _GEN_91; // @[Cache.scala 268:{40,40}]
  wire  _GEN_93 = 6'h38 == s2_idx ? plru0_56 : _GEN_92; // @[Cache.scala 268:{40,40}]
  wire  _GEN_94 = 6'h39 == s2_idx ? plru0_57 : _GEN_93; // @[Cache.scala 268:{40,40}]
  wire  _GEN_95 = 6'h3a == s2_idx ? plru0_58 : _GEN_94; // @[Cache.scala 268:{40,40}]
  wire  _GEN_96 = 6'h3b == s2_idx ? plru0_59 : _GEN_95; // @[Cache.scala 268:{40,40}]
  wire  _GEN_97 = 6'h3c == s2_idx ? plru0_60 : _GEN_96; // @[Cache.scala 268:{40,40}]
  wire  _GEN_98 = 6'h3d == s2_idx ? plru0_61 : _GEN_97; // @[Cache.scala 268:{40,40}]
  wire  _GEN_99 = 6'h3e == s2_idx ? plru0_62 : _GEN_98; // @[Cache.scala 268:{40,40}]
  wire  _GEN_100 = 6'h3f == s2_idx ? plru0_63 : _GEN_99; // @[Cache.scala 268:{40,40}]
  wire  _GEN_102 = 6'h1 == s2_idx ? plru1_1 : plru1_0; // @[Cache.scala 268:{25,25}]
  wire  _GEN_103 = 6'h2 == s2_idx ? plru1_2 : _GEN_102; // @[Cache.scala 268:{25,25}]
  wire  _GEN_104 = 6'h3 == s2_idx ? plru1_3 : _GEN_103; // @[Cache.scala 268:{25,25}]
  wire  _GEN_105 = 6'h4 == s2_idx ? plru1_4 : _GEN_104; // @[Cache.scala 268:{25,25}]
  wire  _GEN_106 = 6'h5 == s2_idx ? plru1_5 : _GEN_105; // @[Cache.scala 268:{25,25}]
  wire  _GEN_107 = 6'h6 == s2_idx ? plru1_6 : _GEN_106; // @[Cache.scala 268:{25,25}]
  wire  _GEN_108 = 6'h7 == s2_idx ? plru1_7 : _GEN_107; // @[Cache.scala 268:{25,25}]
  wire  _GEN_109 = 6'h8 == s2_idx ? plru1_8 : _GEN_108; // @[Cache.scala 268:{25,25}]
  wire  _GEN_110 = 6'h9 == s2_idx ? plru1_9 : _GEN_109; // @[Cache.scala 268:{25,25}]
  wire  _GEN_111 = 6'ha == s2_idx ? plru1_10 : _GEN_110; // @[Cache.scala 268:{25,25}]
  wire  _GEN_112 = 6'hb == s2_idx ? plru1_11 : _GEN_111; // @[Cache.scala 268:{25,25}]
  wire  _GEN_113 = 6'hc == s2_idx ? plru1_12 : _GEN_112; // @[Cache.scala 268:{25,25}]
  wire  _GEN_114 = 6'hd == s2_idx ? plru1_13 : _GEN_113; // @[Cache.scala 268:{25,25}]
  wire  _GEN_115 = 6'he == s2_idx ? plru1_14 : _GEN_114; // @[Cache.scala 268:{25,25}]
  wire  _GEN_116 = 6'hf == s2_idx ? plru1_15 : _GEN_115; // @[Cache.scala 268:{25,25}]
  wire  _GEN_117 = 6'h10 == s2_idx ? plru1_16 : _GEN_116; // @[Cache.scala 268:{25,25}]
  wire  _GEN_118 = 6'h11 == s2_idx ? plru1_17 : _GEN_117; // @[Cache.scala 268:{25,25}]
  wire  _GEN_119 = 6'h12 == s2_idx ? plru1_18 : _GEN_118; // @[Cache.scala 268:{25,25}]
  wire  _GEN_120 = 6'h13 == s2_idx ? plru1_19 : _GEN_119; // @[Cache.scala 268:{25,25}]
  wire  _GEN_121 = 6'h14 == s2_idx ? plru1_20 : _GEN_120; // @[Cache.scala 268:{25,25}]
  wire  _GEN_122 = 6'h15 == s2_idx ? plru1_21 : _GEN_121; // @[Cache.scala 268:{25,25}]
  wire  _GEN_123 = 6'h16 == s2_idx ? plru1_22 : _GEN_122; // @[Cache.scala 268:{25,25}]
  wire  _GEN_124 = 6'h17 == s2_idx ? plru1_23 : _GEN_123; // @[Cache.scala 268:{25,25}]
  wire  _GEN_125 = 6'h18 == s2_idx ? plru1_24 : _GEN_124; // @[Cache.scala 268:{25,25}]
  wire  _GEN_126 = 6'h19 == s2_idx ? plru1_25 : _GEN_125; // @[Cache.scala 268:{25,25}]
  wire  _GEN_127 = 6'h1a == s2_idx ? plru1_26 : _GEN_126; // @[Cache.scala 268:{25,25}]
  wire  _GEN_128 = 6'h1b == s2_idx ? plru1_27 : _GEN_127; // @[Cache.scala 268:{25,25}]
  wire  _GEN_129 = 6'h1c == s2_idx ? plru1_28 : _GEN_128; // @[Cache.scala 268:{25,25}]
  wire  _GEN_130 = 6'h1d == s2_idx ? plru1_29 : _GEN_129; // @[Cache.scala 268:{25,25}]
  wire  _GEN_131 = 6'h1e == s2_idx ? plru1_30 : _GEN_130; // @[Cache.scala 268:{25,25}]
  wire  _GEN_132 = 6'h1f == s2_idx ? plru1_31 : _GEN_131; // @[Cache.scala 268:{25,25}]
  wire  _GEN_133 = 6'h20 == s2_idx ? plru1_32 : _GEN_132; // @[Cache.scala 268:{25,25}]
  wire  _GEN_134 = 6'h21 == s2_idx ? plru1_33 : _GEN_133; // @[Cache.scala 268:{25,25}]
  wire  _GEN_135 = 6'h22 == s2_idx ? plru1_34 : _GEN_134; // @[Cache.scala 268:{25,25}]
  wire  _GEN_136 = 6'h23 == s2_idx ? plru1_35 : _GEN_135; // @[Cache.scala 268:{25,25}]
  wire  _GEN_137 = 6'h24 == s2_idx ? plru1_36 : _GEN_136; // @[Cache.scala 268:{25,25}]
  wire  _GEN_138 = 6'h25 == s2_idx ? plru1_37 : _GEN_137; // @[Cache.scala 268:{25,25}]
  wire  _GEN_139 = 6'h26 == s2_idx ? plru1_38 : _GEN_138; // @[Cache.scala 268:{25,25}]
  wire  _GEN_140 = 6'h27 == s2_idx ? plru1_39 : _GEN_139; // @[Cache.scala 268:{25,25}]
  wire  _GEN_141 = 6'h28 == s2_idx ? plru1_40 : _GEN_140; // @[Cache.scala 268:{25,25}]
  wire  _GEN_142 = 6'h29 == s2_idx ? plru1_41 : _GEN_141; // @[Cache.scala 268:{25,25}]
  wire  _GEN_143 = 6'h2a == s2_idx ? plru1_42 : _GEN_142; // @[Cache.scala 268:{25,25}]
  wire  _GEN_144 = 6'h2b == s2_idx ? plru1_43 : _GEN_143; // @[Cache.scala 268:{25,25}]
  wire  _GEN_145 = 6'h2c == s2_idx ? plru1_44 : _GEN_144; // @[Cache.scala 268:{25,25}]
  wire  _GEN_146 = 6'h2d == s2_idx ? plru1_45 : _GEN_145; // @[Cache.scala 268:{25,25}]
  wire  _GEN_147 = 6'h2e == s2_idx ? plru1_46 : _GEN_146; // @[Cache.scala 268:{25,25}]
  wire  _GEN_148 = 6'h2f == s2_idx ? plru1_47 : _GEN_147; // @[Cache.scala 268:{25,25}]
  wire  _GEN_149 = 6'h30 == s2_idx ? plru1_48 : _GEN_148; // @[Cache.scala 268:{25,25}]
  wire  _GEN_150 = 6'h31 == s2_idx ? plru1_49 : _GEN_149; // @[Cache.scala 268:{25,25}]
  wire  _GEN_151 = 6'h32 == s2_idx ? plru1_50 : _GEN_150; // @[Cache.scala 268:{25,25}]
  wire  _GEN_152 = 6'h33 == s2_idx ? plru1_51 : _GEN_151; // @[Cache.scala 268:{25,25}]
  wire  _GEN_153 = 6'h34 == s2_idx ? plru1_52 : _GEN_152; // @[Cache.scala 268:{25,25}]
  wire  _GEN_154 = 6'h35 == s2_idx ? plru1_53 : _GEN_153; // @[Cache.scala 268:{25,25}]
  wire  _GEN_155 = 6'h36 == s2_idx ? plru1_54 : _GEN_154; // @[Cache.scala 268:{25,25}]
  wire  _GEN_156 = 6'h37 == s2_idx ? plru1_55 : _GEN_155; // @[Cache.scala 268:{25,25}]
  wire  _GEN_157 = 6'h38 == s2_idx ? plru1_56 : _GEN_156; // @[Cache.scala 268:{25,25}]
  wire  _GEN_158 = 6'h39 == s2_idx ? plru1_57 : _GEN_157; // @[Cache.scala 268:{25,25}]
  wire  _GEN_159 = 6'h3a == s2_idx ? plru1_58 : _GEN_158; // @[Cache.scala 268:{25,25}]
  wire  _GEN_160 = 6'h3b == s2_idx ? plru1_59 : _GEN_159; // @[Cache.scala 268:{25,25}]
  wire  _GEN_161 = 6'h3c == s2_idx ? plru1_60 : _GEN_160; // @[Cache.scala 268:{25,25}]
  wire  _GEN_162 = 6'h3d == s2_idx ? plru1_61 : _GEN_161; // @[Cache.scala 268:{25,25}]
  wire  _GEN_163 = 6'h3e == s2_idx ? plru1_62 : _GEN_162; // @[Cache.scala 268:{25,25}]
  wire  _GEN_164 = 6'h3f == s2_idx ? plru1_63 : _GEN_163; // @[Cache.scala 268:{25,25}]
  wire  _GEN_166 = 6'h1 == s2_idx ? plru2_1 : plru2_0; // @[Cache.scala 268:{25,25}]
  wire  _GEN_167 = 6'h2 == s2_idx ? plru2_2 : _GEN_166; // @[Cache.scala 268:{25,25}]
  wire  _GEN_168 = 6'h3 == s2_idx ? plru2_3 : _GEN_167; // @[Cache.scala 268:{25,25}]
  wire  _GEN_169 = 6'h4 == s2_idx ? plru2_4 : _GEN_168; // @[Cache.scala 268:{25,25}]
  wire  _GEN_170 = 6'h5 == s2_idx ? plru2_5 : _GEN_169; // @[Cache.scala 268:{25,25}]
  wire  _GEN_171 = 6'h6 == s2_idx ? plru2_6 : _GEN_170; // @[Cache.scala 268:{25,25}]
  wire  _GEN_172 = 6'h7 == s2_idx ? plru2_7 : _GEN_171; // @[Cache.scala 268:{25,25}]
  wire  _GEN_173 = 6'h8 == s2_idx ? plru2_8 : _GEN_172; // @[Cache.scala 268:{25,25}]
  wire  _GEN_174 = 6'h9 == s2_idx ? plru2_9 : _GEN_173; // @[Cache.scala 268:{25,25}]
  wire  _GEN_175 = 6'ha == s2_idx ? plru2_10 : _GEN_174; // @[Cache.scala 268:{25,25}]
  wire  _GEN_176 = 6'hb == s2_idx ? plru2_11 : _GEN_175; // @[Cache.scala 268:{25,25}]
  wire  _GEN_177 = 6'hc == s2_idx ? plru2_12 : _GEN_176; // @[Cache.scala 268:{25,25}]
  wire  _GEN_178 = 6'hd == s2_idx ? plru2_13 : _GEN_177; // @[Cache.scala 268:{25,25}]
  wire  _GEN_179 = 6'he == s2_idx ? plru2_14 : _GEN_178; // @[Cache.scala 268:{25,25}]
  wire  _GEN_180 = 6'hf == s2_idx ? plru2_15 : _GEN_179; // @[Cache.scala 268:{25,25}]
  wire  _GEN_181 = 6'h10 == s2_idx ? plru2_16 : _GEN_180; // @[Cache.scala 268:{25,25}]
  wire  _GEN_182 = 6'h11 == s2_idx ? plru2_17 : _GEN_181; // @[Cache.scala 268:{25,25}]
  wire  _GEN_183 = 6'h12 == s2_idx ? plru2_18 : _GEN_182; // @[Cache.scala 268:{25,25}]
  wire  _GEN_184 = 6'h13 == s2_idx ? plru2_19 : _GEN_183; // @[Cache.scala 268:{25,25}]
  wire  _GEN_185 = 6'h14 == s2_idx ? plru2_20 : _GEN_184; // @[Cache.scala 268:{25,25}]
  wire  _GEN_186 = 6'h15 == s2_idx ? plru2_21 : _GEN_185; // @[Cache.scala 268:{25,25}]
  wire  _GEN_187 = 6'h16 == s2_idx ? plru2_22 : _GEN_186; // @[Cache.scala 268:{25,25}]
  wire  _GEN_188 = 6'h17 == s2_idx ? plru2_23 : _GEN_187; // @[Cache.scala 268:{25,25}]
  wire  _GEN_189 = 6'h18 == s2_idx ? plru2_24 : _GEN_188; // @[Cache.scala 268:{25,25}]
  wire  _GEN_190 = 6'h19 == s2_idx ? plru2_25 : _GEN_189; // @[Cache.scala 268:{25,25}]
  wire  _GEN_191 = 6'h1a == s2_idx ? plru2_26 : _GEN_190; // @[Cache.scala 268:{25,25}]
  wire  _GEN_192 = 6'h1b == s2_idx ? plru2_27 : _GEN_191; // @[Cache.scala 268:{25,25}]
  wire  _GEN_193 = 6'h1c == s2_idx ? plru2_28 : _GEN_192; // @[Cache.scala 268:{25,25}]
  wire  _GEN_194 = 6'h1d == s2_idx ? plru2_29 : _GEN_193; // @[Cache.scala 268:{25,25}]
  wire  _GEN_195 = 6'h1e == s2_idx ? plru2_30 : _GEN_194; // @[Cache.scala 268:{25,25}]
  wire  _GEN_196 = 6'h1f == s2_idx ? plru2_31 : _GEN_195; // @[Cache.scala 268:{25,25}]
  wire  _GEN_197 = 6'h20 == s2_idx ? plru2_32 : _GEN_196; // @[Cache.scala 268:{25,25}]
  wire  _GEN_198 = 6'h21 == s2_idx ? plru2_33 : _GEN_197; // @[Cache.scala 268:{25,25}]
  wire  _GEN_199 = 6'h22 == s2_idx ? plru2_34 : _GEN_198; // @[Cache.scala 268:{25,25}]
  wire  _GEN_200 = 6'h23 == s2_idx ? plru2_35 : _GEN_199; // @[Cache.scala 268:{25,25}]
  wire  _GEN_201 = 6'h24 == s2_idx ? plru2_36 : _GEN_200; // @[Cache.scala 268:{25,25}]
  wire  _GEN_202 = 6'h25 == s2_idx ? plru2_37 : _GEN_201; // @[Cache.scala 268:{25,25}]
  wire  _GEN_203 = 6'h26 == s2_idx ? plru2_38 : _GEN_202; // @[Cache.scala 268:{25,25}]
  wire  _GEN_204 = 6'h27 == s2_idx ? plru2_39 : _GEN_203; // @[Cache.scala 268:{25,25}]
  wire  _GEN_205 = 6'h28 == s2_idx ? plru2_40 : _GEN_204; // @[Cache.scala 268:{25,25}]
  wire  _GEN_206 = 6'h29 == s2_idx ? plru2_41 : _GEN_205; // @[Cache.scala 268:{25,25}]
  wire  _GEN_207 = 6'h2a == s2_idx ? plru2_42 : _GEN_206; // @[Cache.scala 268:{25,25}]
  wire  _GEN_208 = 6'h2b == s2_idx ? plru2_43 : _GEN_207; // @[Cache.scala 268:{25,25}]
  wire  _GEN_209 = 6'h2c == s2_idx ? plru2_44 : _GEN_208; // @[Cache.scala 268:{25,25}]
  wire  _GEN_210 = 6'h2d == s2_idx ? plru2_45 : _GEN_209; // @[Cache.scala 268:{25,25}]
  wire  _GEN_211 = 6'h2e == s2_idx ? plru2_46 : _GEN_210; // @[Cache.scala 268:{25,25}]
  wire  _GEN_212 = 6'h2f == s2_idx ? plru2_47 : _GEN_211; // @[Cache.scala 268:{25,25}]
  wire  _GEN_213 = 6'h30 == s2_idx ? plru2_48 : _GEN_212; // @[Cache.scala 268:{25,25}]
  wire  _GEN_214 = 6'h31 == s2_idx ? plru2_49 : _GEN_213; // @[Cache.scala 268:{25,25}]
  wire  _GEN_215 = 6'h32 == s2_idx ? plru2_50 : _GEN_214; // @[Cache.scala 268:{25,25}]
  wire  _GEN_216 = 6'h33 == s2_idx ? plru2_51 : _GEN_215; // @[Cache.scala 268:{25,25}]
  wire  _GEN_217 = 6'h34 == s2_idx ? plru2_52 : _GEN_216; // @[Cache.scala 268:{25,25}]
  wire  _GEN_218 = 6'h35 == s2_idx ? plru2_53 : _GEN_217; // @[Cache.scala 268:{25,25}]
  wire  _GEN_219 = 6'h36 == s2_idx ? plru2_54 : _GEN_218; // @[Cache.scala 268:{25,25}]
  wire  _GEN_220 = 6'h37 == s2_idx ? plru2_55 : _GEN_219; // @[Cache.scala 268:{25,25}]
  wire  _GEN_221 = 6'h38 == s2_idx ? plru2_56 : _GEN_220; // @[Cache.scala 268:{25,25}]
  wire  _GEN_222 = 6'h39 == s2_idx ? plru2_57 : _GEN_221; // @[Cache.scala 268:{25,25}]
  wire  _GEN_223 = 6'h3a == s2_idx ? plru2_58 : _GEN_222; // @[Cache.scala 268:{25,25}]
  wire  _GEN_224 = 6'h3b == s2_idx ? plru2_59 : _GEN_223; // @[Cache.scala 268:{25,25}]
  wire  _GEN_225 = 6'h3c == s2_idx ? plru2_60 : _GEN_224; // @[Cache.scala 268:{25,25}]
  wire  _GEN_226 = 6'h3d == s2_idx ? plru2_61 : _GEN_225; // @[Cache.scala 268:{25,25}]
  wire  _GEN_227 = 6'h3e == s2_idx ? plru2_62 : _GEN_226; // @[Cache.scala 268:{25,25}]
  wire  _GEN_228 = 6'h3f == s2_idx ? plru2_63 : _GEN_227; // @[Cache.scala 268:{25,25}]
  wire  _T_16 = ~_GEN_100 ? _GEN_164 : _GEN_228; // @[Cache.scala 268:25]
  wire [1:0] replace_way = {_GEN_100,_T_16}; // @[Cat.scala 30:58]
  wire  _GEN_9 = 2'h1 == replace_way ? REG_5 : REG_4; // @[Cache.scala 262:{18,18}]
  wire  _GEN_10 = 2'h2 == replace_way ? REG_6 : _GEN_9; // @[Cache.scala 262:{18,18}]
  wire [20:0] _GEN_13 = 2'h1 == replace_way ? tag_out_1 : tag_out_0; // @[Cache.scala 263:{18,18}]
  wire [20:0] _GEN_14 = 2'h2 == replace_way ? tag_out_2 : _GEN_13; // @[Cache.scala 263:{18,18}]
  wire [127:0] _GEN_17 = 2'h1 == replace_way ? sram_out_1 : sram_out_0; // @[Cache.scala 264:{18,18}]
  wire [127:0] _GEN_18 = 2'h2 == replace_way ? sram_out_2 : _GEN_17; // @[Cache.scala 264:{18,18}]
  wire  _GEN_27 = pipeline_ready ? io_in_req_bits_wen : s2_wen; // @[Cache.scala 246:24 249:14 219:25]
  reg [63:0] wdata1; // @[Cache.scala 270:23]
  reg [63:0] wdata2; // @[Cache.scala 271:23]
  reg  REG_10; // @[Cache.scala 320:20]
  wire [63:0] _T_36 = s2_offs ? _GEN_7[127:64] : _GEN_7[63:0]; // @[Cache.scala 321:34]
  wire [63:0] _T_40 = s2_offs ? s2_reg_rdata[127:64] : s2_reg_rdata[63:0]; // @[Cache.scala 323:34]
  wire [63:0] _GEN_229 = REG_10 ? _T_36 : _T_40; // @[Cache.scala 320:37 321:28 323:28]
  reg  REG_11; // @[Cache.scala 325:20]
  wire  _T_42 = ~s2_way[1]; // @[Cache.scala 136:19]
  wire  _GEN_230 = 6'h0 == s2_idx ? ~s2_way[1] : plru0_0; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_231 = 6'h1 == s2_idx ? ~s2_way[1] : plru0_1; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_232 = 6'h2 == s2_idx ? ~s2_way[1] : plru0_2; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_233 = 6'h3 == s2_idx ? ~s2_way[1] : plru0_3; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_234 = 6'h4 == s2_idx ? ~s2_way[1] : plru0_4; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_235 = 6'h5 == s2_idx ? ~s2_way[1] : plru0_5; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_236 = 6'h6 == s2_idx ? ~s2_way[1] : plru0_6; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_237 = 6'h7 == s2_idx ? ~s2_way[1] : plru0_7; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_238 = 6'h8 == s2_idx ? ~s2_way[1] : plru0_8; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_239 = 6'h9 == s2_idx ? ~s2_way[1] : plru0_9; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_240 = 6'ha == s2_idx ? ~s2_way[1] : plru0_10; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_241 = 6'hb == s2_idx ? ~s2_way[1] : plru0_11; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_242 = 6'hc == s2_idx ? ~s2_way[1] : plru0_12; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_243 = 6'hd == s2_idx ? ~s2_way[1] : plru0_13; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_244 = 6'he == s2_idx ? ~s2_way[1] : plru0_14; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_245 = 6'hf == s2_idx ? ~s2_way[1] : plru0_15; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_246 = 6'h10 == s2_idx ? ~s2_way[1] : plru0_16; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_247 = 6'h11 == s2_idx ? ~s2_way[1] : plru0_17; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_248 = 6'h12 == s2_idx ? ~s2_way[1] : plru0_18; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_249 = 6'h13 == s2_idx ? ~s2_way[1] : plru0_19; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_250 = 6'h14 == s2_idx ? ~s2_way[1] : plru0_20; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_251 = 6'h15 == s2_idx ? ~s2_way[1] : plru0_21; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_252 = 6'h16 == s2_idx ? ~s2_way[1] : plru0_22; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_253 = 6'h17 == s2_idx ? ~s2_way[1] : plru0_23; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_254 = 6'h18 == s2_idx ? ~s2_way[1] : plru0_24; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_255 = 6'h19 == s2_idx ? ~s2_way[1] : plru0_25; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_256 = 6'h1a == s2_idx ? ~s2_way[1] : plru0_26; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_257 = 6'h1b == s2_idx ? ~s2_way[1] : plru0_27; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_258 = 6'h1c == s2_idx ? ~s2_way[1] : plru0_28; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_259 = 6'h1d == s2_idx ? ~s2_way[1] : plru0_29; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_260 = 6'h1e == s2_idx ? ~s2_way[1] : plru0_30; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_261 = 6'h1f == s2_idx ? ~s2_way[1] : plru0_31; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_262 = 6'h20 == s2_idx ? ~s2_way[1] : plru0_32; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_263 = 6'h21 == s2_idx ? ~s2_way[1] : plru0_33; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_264 = 6'h22 == s2_idx ? ~s2_way[1] : plru0_34; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_265 = 6'h23 == s2_idx ? ~s2_way[1] : plru0_35; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_266 = 6'h24 == s2_idx ? ~s2_way[1] : plru0_36; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_267 = 6'h25 == s2_idx ? ~s2_way[1] : plru0_37; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_268 = 6'h26 == s2_idx ? ~s2_way[1] : plru0_38; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_269 = 6'h27 == s2_idx ? ~s2_way[1] : plru0_39; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_270 = 6'h28 == s2_idx ? ~s2_way[1] : plru0_40; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_271 = 6'h29 == s2_idx ? ~s2_way[1] : plru0_41; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_272 = 6'h2a == s2_idx ? ~s2_way[1] : plru0_42; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_273 = 6'h2b == s2_idx ? ~s2_way[1] : plru0_43; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_274 = 6'h2c == s2_idx ? ~s2_way[1] : plru0_44; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_275 = 6'h2d == s2_idx ? ~s2_way[1] : plru0_45; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_276 = 6'h2e == s2_idx ? ~s2_way[1] : plru0_46; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_277 = 6'h2f == s2_idx ? ~s2_way[1] : plru0_47; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_278 = 6'h30 == s2_idx ? ~s2_way[1] : plru0_48; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_279 = 6'h31 == s2_idx ? ~s2_way[1] : plru0_49; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_280 = 6'h32 == s2_idx ? ~s2_way[1] : plru0_50; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_281 = 6'h33 == s2_idx ? ~s2_way[1] : plru0_51; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_282 = 6'h34 == s2_idx ? ~s2_way[1] : plru0_52; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_283 = 6'h35 == s2_idx ? ~s2_way[1] : plru0_53; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_284 = 6'h36 == s2_idx ? ~s2_way[1] : plru0_54; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_285 = 6'h37 == s2_idx ? ~s2_way[1] : plru0_55; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_286 = 6'h38 == s2_idx ? ~s2_way[1] : plru0_56; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_287 = 6'h39 == s2_idx ? ~s2_way[1] : plru0_57; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_288 = 6'h3a == s2_idx ? ~s2_way[1] : plru0_58; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_289 = 6'h3b == s2_idx ? ~s2_way[1] : plru0_59; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_290 = 6'h3c == s2_idx ? ~s2_way[1] : plru0_60; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_291 = 6'h3d == s2_idx ? ~s2_way[1] : plru0_61; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_292 = 6'h3e == s2_idx ? ~s2_way[1] : plru0_62; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_293 = 6'h3f == s2_idx ? ~s2_way[1] : plru0_63; // @[Cache.scala 136:{16,16} 129:22]
  wire  _T_46 = ~s2_way[0]; // @[Cache.scala 138:21]
  wire  _GEN_294 = 6'h0 == s2_idx ? ~s2_way[0] : plru1_0; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_295 = 6'h1 == s2_idx ? ~s2_way[0] : plru1_1; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_296 = 6'h2 == s2_idx ? ~s2_way[0] : plru1_2; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_297 = 6'h3 == s2_idx ? ~s2_way[0] : plru1_3; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_298 = 6'h4 == s2_idx ? ~s2_way[0] : plru1_4; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_299 = 6'h5 == s2_idx ? ~s2_way[0] : plru1_5; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_300 = 6'h6 == s2_idx ? ~s2_way[0] : plru1_6; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_301 = 6'h7 == s2_idx ? ~s2_way[0] : plru1_7; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_302 = 6'h8 == s2_idx ? ~s2_way[0] : plru1_8; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_303 = 6'h9 == s2_idx ? ~s2_way[0] : plru1_9; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_304 = 6'ha == s2_idx ? ~s2_way[0] : plru1_10; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_305 = 6'hb == s2_idx ? ~s2_way[0] : plru1_11; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_306 = 6'hc == s2_idx ? ~s2_way[0] : plru1_12; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_307 = 6'hd == s2_idx ? ~s2_way[0] : plru1_13; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_308 = 6'he == s2_idx ? ~s2_way[0] : plru1_14; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_309 = 6'hf == s2_idx ? ~s2_way[0] : plru1_15; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_310 = 6'h10 == s2_idx ? ~s2_way[0] : plru1_16; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_311 = 6'h11 == s2_idx ? ~s2_way[0] : plru1_17; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_312 = 6'h12 == s2_idx ? ~s2_way[0] : plru1_18; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_313 = 6'h13 == s2_idx ? ~s2_way[0] : plru1_19; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_314 = 6'h14 == s2_idx ? ~s2_way[0] : plru1_20; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_315 = 6'h15 == s2_idx ? ~s2_way[0] : plru1_21; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_316 = 6'h16 == s2_idx ? ~s2_way[0] : plru1_22; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_317 = 6'h17 == s2_idx ? ~s2_way[0] : plru1_23; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_318 = 6'h18 == s2_idx ? ~s2_way[0] : plru1_24; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_319 = 6'h19 == s2_idx ? ~s2_way[0] : plru1_25; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_320 = 6'h1a == s2_idx ? ~s2_way[0] : plru1_26; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_321 = 6'h1b == s2_idx ? ~s2_way[0] : plru1_27; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_322 = 6'h1c == s2_idx ? ~s2_way[0] : plru1_28; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_323 = 6'h1d == s2_idx ? ~s2_way[0] : plru1_29; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_324 = 6'h1e == s2_idx ? ~s2_way[0] : plru1_30; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_325 = 6'h1f == s2_idx ? ~s2_way[0] : plru1_31; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_326 = 6'h20 == s2_idx ? ~s2_way[0] : plru1_32; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_327 = 6'h21 == s2_idx ? ~s2_way[0] : plru1_33; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_328 = 6'h22 == s2_idx ? ~s2_way[0] : plru1_34; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_329 = 6'h23 == s2_idx ? ~s2_way[0] : plru1_35; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_330 = 6'h24 == s2_idx ? ~s2_way[0] : plru1_36; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_331 = 6'h25 == s2_idx ? ~s2_way[0] : plru1_37; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_332 = 6'h26 == s2_idx ? ~s2_way[0] : plru1_38; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_333 = 6'h27 == s2_idx ? ~s2_way[0] : plru1_39; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_334 = 6'h28 == s2_idx ? ~s2_way[0] : plru1_40; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_335 = 6'h29 == s2_idx ? ~s2_way[0] : plru1_41; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_336 = 6'h2a == s2_idx ? ~s2_way[0] : plru1_42; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_337 = 6'h2b == s2_idx ? ~s2_way[0] : plru1_43; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_338 = 6'h2c == s2_idx ? ~s2_way[0] : plru1_44; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_339 = 6'h2d == s2_idx ? ~s2_way[0] : plru1_45; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_340 = 6'h2e == s2_idx ? ~s2_way[0] : plru1_46; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_341 = 6'h2f == s2_idx ? ~s2_way[0] : plru1_47; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_342 = 6'h30 == s2_idx ? ~s2_way[0] : plru1_48; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_343 = 6'h31 == s2_idx ? ~s2_way[0] : plru1_49; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_344 = 6'h32 == s2_idx ? ~s2_way[0] : plru1_50; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_345 = 6'h33 == s2_idx ? ~s2_way[0] : plru1_51; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_346 = 6'h34 == s2_idx ? ~s2_way[0] : plru1_52; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_347 = 6'h35 == s2_idx ? ~s2_way[0] : plru1_53; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_348 = 6'h36 == s2_idx ? ~s2_way[0] : plru1_54; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_349 = 6'h37 == s2_idx ? ~s2_way[0] : plru1_55; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_350 = 6'h38 == s2_idx ? ~s2_way[0] : plru1_56; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_351 = 6'h39 == s2_idx ? ~s2_way[0] : plru1_57; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_352 = 6'h3a == s2_idx ? ~s2_way[0] : plru1_58; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_353 = 6'h3b == s2_idx ? ~s2_way[0] : plru1_59; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_354 = 6'h3c == s2_idx ? ~s2_way[0] : plru1_60; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_355 = 6'h3d == s2_idx ? ~s2_way[0] : plru1_61; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_356 = 6'h3e == s2_idx ? ~s2_way[0] : plru1_62; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_357 = 6'h3f == s2_idx ? ~s2_way[0] : plru1_63; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_358 = 6'h0 == s2_idx ? _T_46 : plru2_0; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_359 = 6'h1 == s2_idx ? _T_46 : plru2_1; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_360 = 6'h2 == s2_idx ? _T_46 : plru2_2; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_361 = 6'h3 == s2_idx ? _T_46 : plru2_3; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_362 = 6'h4 == s2_idx ? _T_46 : plru2_4; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_363 = 6'h5 == s2_idx ? _T_46 : plru2_5; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_364 = 6'h6 == s2_idx ? _T_46 : plru2_6; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_365 = 6'h7 == s2_idx ? _T_46 : plru2_7; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_366 = 6'h8 == s2_idx ? _T_46 : plru2_8; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_367 = 6'h9 == s2_idx ? _T_46 : plru2_9; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_368 = 6'ha == s2_idx ? _T_46 : plru2_10; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_369 = 6'hb == s2_idx ? _T_46 : plru2_11; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_370 = 6'hc == s2_idx ? _T_46 : plru2_12; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_371 = 6'hd == s2_idx ? _T_46 : plru2_13; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_372 = 6'he == s2_idx ? _T_46 : plru2_14; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_373 = 6'hf == s2_idx ? _T_46 : plru2_15; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_374 = 6'h10 == s2_idx ? _T_46 : plru2_16; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_375 = 6'h11 == s2_idx ? _T_46 : plru2_17; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_376 = 6'h12 == s2_idx ? _T_46 : plru2_18; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_377 = 6'h13 == s2_idx ? _T_46 : plru2_19; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_378 = 6'h14 == s2_idx ? _T_46 : plru2_20; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_379 = 6'h15 == s2_idx ? _T_46 : plru2_21; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_380 = 6'h16 == s2_idx ? _T_46 : plru2_22; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_381 = 6'h17 == s2_idx ? _T_46 : plru2_23; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_382 = 6'h18 == s2_idx ? _T_46 : plru2_24; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_383 = 6'h19 == s2_idx ? _T_46 : plru2_25; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_384 = 6'h1a == s2_idx ? _T_46 : plru2_26; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_385 = 6'h1b == s2_idx ? _T_46 : plru2_27; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_386 = 6'h1c == s2_idx ? _T_46 : plru2_28; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_387 = 6'h1d == s2_idx ? _T_46 : plru2_29; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_388 = 6'h1e == s2_idx ? _T_46 : plru2_30; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_389 = 6'h1f == s2_idx ? _T_46 : plru2_31; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_390 = 6'h20 == s2_idx ? _T_46 : plru2_32; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_391 = 6'h21 == s2_idx ? _T_46 : plru2_33; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_392 = 6'h22 == s2_idx ? _T_46 : plru2_34; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_393 = 6'h23 == s2_idx ? _T_46 : plru2_35; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_394 = 6'h24 == s2_idx ? _T_46 : plru2_36; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_395 = 6'h25 == s2_idx ? _T_46 : plru2_37; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_396 = 6'h26 == s2_idx ? _T_46 : plru2_38; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_397 = 6'h27 == s2_idx ? _T_46 : plru2_39; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_398 = 6'h28 == s2_idx ? _T_46 : plru2_40; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_399 = 6'h29 == s2_idx ? _T_46 : plru2_41; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_400 = 6'h2a == s2_idx ? _T_46 : plru2_42; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_401 = 6'h2b == s2_idx ? _T_46 : plru2_43; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_402 = 6'h2c == s2_idx ? _T_46 : plru2_44; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_403 = 6'h2d == s2_idx ? _T_46 : plru2_45; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_404 = 6'h2e == s2_idx ? _T_46 : plru2_46; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_405 = 6'h2f == s2_idx ? _T_46 : plru2_47; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_406 = 6'h30 == s2_idx ? _T_46 : plru2_48; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_407 = 6'h31 == s2_idx ? _T_46 : plru2_49; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_408 = 6'h32 == s2_idx ? _T_46 : plru2_50; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_409 = 6'h33 == s2_idx ? _T_46 : plru2_51; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_410 = 6'h34 == s2_idx ? _T_46 : plru2_52; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_411 = 6'h35 == s2_idx ? _T_46 : plru2_53; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_412 = 6'h36 == s2_idx ? _T_46 : plru2_54; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_413 = 6'h37 == s2_idx ? _T_46 : plru2_55; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_414 = 6'h38 == s2_idx ? _T_46 : plru2_56; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_415 = 6'h39 == s2_idx ? _T_46 : plru2_57; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_416 = 6'h3a == s2_idx ? _T_46 : plru2_58; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_417 = 6'h3b == s2_idx ? _T_46 : plru2_59; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_418 = 6'h3c == s2_idx ? _T_46 : plru2_60; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_419 = 6'h3d == s2_idx ? _T_46 : plru2_61; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_420 = 6'h3e == s2_idx ? _T_46 : plru2_62; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_421 = 6'h3f == s2_idx ? _T_46 : plru2_63; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_422 = _T_42 ? _GEN_294 : plru1_0; // @[Cache.scala 131:22 137:27]
  wire  _GEN_423 = _T_42 ? _GEN_295 : plru1_1; // @[Cache.scala 131:22 137:27]
  wire  _GEN_424 = _T_42 ? _GEN_296 : plru1_2; // @[Cache.scala 131:22 137:27]
  wire  _GEN_425 = _T_42 ? _GEN_297 : plru1_3; // @[Cache.scala 131:22 137:27]
  wire  _GEN_426 = _T_42 ? _GEN_298 : plru1_4; // @[Cache.scala 131:22 137:27]
  wire  _GEN_427 = _T_42 ? _GEN_299 : plru1_5; // @[Cache.scala 131:22 137:27]
  wire  _GEN_428 = _T_42 ? _GEN_300 : plru1_6; // @[Cache.scala 131:22 137:27]
  wire  _GEN_429 = _T_42 ? _GEN_301 : plru1_7; // @[Cache.scala 131:22 137:27]
  wire  _GEN_430 = _T_42 ? _GEN_302 : plru1_8; // @[Cache.scala 131:22 137:27]
  wire  _GEN_431 = _T_42 ? _GEN_303 : plru1_9; // @[Cache.scala 131:22 137:27]
  wire  _GEN_432 = _T_42 ? _GEN_304 : plru1_10; // @[Cache.scala 131:22 137:27]
  wire  _GEN_433 = _T_42 ? _GEN_305 : plru1_11; // @[Cache.scala 131:22 137:27]
  wire  _GEN_434 = _T_42 ? _GEN_306 : plru1_12; // @[Cache.scala 131:22 137:27]
  wire  _GEN_435 = _T_42 ? _GEN_307 : plru1_13; // @[Cache.scala 131:22 137:27]
  wire  _GEN_436 = _T_42 ? _GEN_308 : plru1_14; // @[Cache.scala 131:22 137:27]
  wire  _GEN_437 = _T_42 ? _GEN_309 : plru1_15; // @[Cache.scala 131:22 137:27]
  wire  _GEN_438 = _T_42 ? _GEN_310 : plru1_16; // @[Cache.scala 131:22 137:27]
  wire  _GEN_439 = _T_42 ? _GEN_311 : plru1_17; // @[Cache.scala 131:22 137:27]
  wire  _GEN_440 = _T_42 ? _GEN_312 : plru1_18; // @[Cache.scala 131:22 137:27]
  wire  _GEN_441 = _T_42 ? _GEN_313 : plru1_19; // @[Cache.scala 131:22 137:27]
  wire  _GEN_442 = _T_42 ? _GEN_314 : plru1_20; // @[Cache.scala 131:22 137:27]
  wire  _GEN_443 = _T_42 ? _GEN_315 : plru1_21; // @[Cache.scala 131:22 137:27]
  wire  _GEN_444 = _T_42 ? _GEN_316 : plru1_22; // @[Cache.scala 131:22 137:27]
  wire  _GEN_445 = _T_42 ? _GEN_317 : plru1_23; // @[Cache.scala 131:22 137:27]
  wire  _GEN_446 = _T_42 ? _GEN_318 : plru1_24; // @[Cache.scala 131:22 137:27]
  wire  _GEN_447 = _T_42 ? _GEN_319 : plru1_25; // @[Cache.scala 131:22 137:27]
  wire  _GEN_448 = _T_42 ? _GEN_320 : plru1_26; // @[Cache.scala 131:22 137:27]
  wire  _GEN_449 = _T_42 ? _GEN_321 : plru1_27; // @[Cache.scala 131:22 137:27]
  wire  _GEN_450 = _T_42 ? _GEN_322 : plru1_28; // @[Cache.scala 131:22 137:27]
  wire  _GEN_451 = _T_42 ? _GEN_323 : plru1_29; // @[Cache.scala 131:22 137:27]
  wire  _GEN_452 = _T_42 ? _GEN_324 : plru1_30; // @[Cache.scala 131:22 137:27]
  wire  _GEN_453 = _T_42 ? _GEN_325 : plru1_31; // @[Cache.scala 131:22 137:27]
  wire  _GEN_454 = _T_42 ? _GEN_326 : plru1_32; // @[Cache.scala 131:22 137:27]
  wire  _GEN_455 = _T_42 ? _GEN_327 : plru1_33; // @[Cache.scala 131:22 137:27]
  wire  _GEN_456 = _T_42 ? _GEN_328 : plru1_34; // @[Cache.scala 131:22 137:27]
  wire  _GEN_457 = _T_42 ? _GEN_329 : plru1_35; // @[Cache.scala 131:22 137:27]
  wire  _GEN_458 = _T_42 ? _GEN_330 : plru1_36; // @[Cache.scala 131:22 137:27]
  wire  _GEN_459 = _T_42 ? _GEN_331 : plru1_37; // @[Cache.scala 131:22 137:27]
  wire  _GEN_460 = _T_42 ? _GEN_332 : plru1_38; // @[Cache.scala 131:22 137:27]
  wire  _GEN_461 = _T_42 ? _GEN_333 : plru1_39; // @[Cache.scala 131:22 137:27]
  wire  _GEN_462 = _T_42 ? _GEN_334 : plru1_40; // @[Cache.scala 131:22 137:27]
  wire  _GEN_463 = _T_42 ? _GEN_335 : plru1_41; // @[Cache.scala 131:22 137:27]
  wire  _GEN_464 = _T_42 ? _GEN_336 : plru1_42; // @[Cache.scala 131:22 137:27]
  wire  _GEN_465 = _T_42 ? _GEN_337 : plru1_43; // @[Cache.scala 131:22 137:27]
  wire  _GEN_466 = _T_42 ? _GEN_338 : plru1_44; // @[Cache.scala 131:22 137:27]
  wire  _GEN_467 = _T_42 ? _GEN_339 : plru1_45; // @[Cache.scala 131:22 137:27]
  wire  _GEN_468 = _T_42 ? _GEN_340 : plru1_46; // @[Cache.scala 131:22 137:27]
  wire  _GEN_469 = _T_42 ? _GEN_341 : plru1_47; // @[Cache.scala 131:22 137:27]
  wire  _GEN_470 = _T_42 ? _GEN_342 : plru1_48; // @[Cache.scala 131:22 137:27]
  wire  _GEN_471 = _T_42 ? _GEN_343 : plru1_49; // @[Cache.scala 131:22 137:27]
  wire  _GEN_472 = _T_42 ? _GEN_344 : plru1_50; // @[Cache.scala 131:22 137:27]
  wire  _GEN_473 = _T_42 ? _GEN_345 : plru1_51; // @[Cache.scala 131:22 137:27]
  wire  _GEN_474 = _T_42 ? _GEN_346 : plru1_52; // @[Cache.scala 131:22 137:27]
  wire  _GEN_475 = _T_42 ? _GEN_347 : plru1_53; // @[Cache.scala 131:22 137:27]
  wire  _GEN_476 = _T_42 ? _GEN_348 : plru1_54; // @[Cache.scala 131:22 137:27]
  wire  _GEN_477 = _T_42 ? _GEN_349 : plru1_55; // @[Cache.scala 131:22 137:27]
  wire  _GEN_478 = _T_42 ? _GEN_350 : plru1_56; // @[Cache.scala 131:22 137:27]
  wire  _GEN_479 = _T_42 ? _GEN_351 : plru1_57; // @[Cache.scala 131:22 137:27]
  wire  _GEN_480 = _T_42 ? _GEN_352 : plru1_58; // @[Cache.scala 131:22 137:27]
  wire  _GEN_481 = _T_42 ? _GEN_353 : plru1_59; // @[Cache.scala 131:22 137:27]
  wire  _GEN_482 = _T_42 ? _GEN_354 : plru1_60; // @[Cache.scala 131:22 137:27]
  wire  _GEN_483 = _T_42 ? _GEN_355 : plru1_61; // @[Cache.scala 131:22 137:27]
  wire  _GEN_484 = _T_42 ? _GEN_356 : plru1_62; // @[Cache.scala 131:22 137:27]
  wire  _GEN_485 = _T_42 ? _GEN_357 : plru1_63; // @[Cache.scala 131:22 137:27]
  wire  _GEN_486 = _T_42 ? plru2_0 : _GEN_358; // @[Cache.scala 133:22 137:27]
  wire  _GEN_487 = _T_42 ? plru2_1 : _GEN_359; // @[Cache.scala 133:22 137:27]
  wire  _GEN_488 = _T_42 ? plru2_2 : _GEN_360; // @[Cache.scala 133:22 137:27]
  wire  _GEN_489 = _T_42 ? plru2_3 : _GEN_361; // @[Cache.scala 133:22 137:27]
  wire  _GEN_490 = _T_42 ? plru2_4 : _GEN_362; // @[Cache.scala 133:22 137:27]
  wire  _GEN_491 = _T_42 ? plru2_5 : _GEN_363; // @[Cache.scala 133:22 137:27]
  wire  _GEN_492 = _T_42 ? plru2_6 : _GEN_364; // @[Cache.scala 133:22 137:27]
  wire  _GEN_493 = _T_42 ? plru2_7 : _GEN_365; // @[Cache.scala 133:22 137:27]
  wire  _GEN_494 = _T_42 ? plru2_8 : _GEN_366; // @[Cache.scala 133:22 137:27]
  wire  _GEN_495 = _T_42 ? plru2_9 : _GEN_367; // @[Cache.scala 133:22 137:27]
  wire  _GEN_496 = _T_42 ? plru2_10 : _GEN_368; // @[Cache.scala 133:22 137:27]
  wire  _GEN_497 = _T_42 ? plru2_11 : _GEN_369; // @[Cache.scala 133:22 137:27]
  wire  _GEN_498 = _T_42 ? plru2_12 : _GEN_370; // @[Cache.scala 133:22 137:27]
  wire  _GEN_499 = _T_42 ? plru2_13 : _GEN_371; // @[Cache.scala 133:22 137:27]
  wire  _GEN_500 = _T_42 ? plru2_14 : _GEN_372; // @[Cache.scala 133:22 137:27]
  wire  _GEN_501 = _T_42 ? plru2_15 : _GEN_373; // @[Cache.scala 133:22 137:27]
  wire  _GEN_502 = _T_42 ? plru2_16 : _GEN_374; // @[Cache.scala 133:22 137:27]
  wire  _GEN_503 = _T_42 ? plru2_17 : _GEN_375; // @[Cache.scala 133:22 137:27]
  wire  _GEN_504 = _T_42 ? plru2_18 : _GEN_376; // @[Cache.scala 133:22 137:27]
  wire  _GEN_505 = _T_42 ? plru2_19 : _GEN_377; // @[Cache.scala 133:22 137:27]
  wire  _GEN_506 = _T_42 ? plru2_20 : _GEN_378; // @[Cache.scala 133:22 137:27]
  wire  _GEN_507 = _T_42 ? plru2_21 : _GEN_379; // @[Cache.scala 133:22 137:27]
  wire  _GEN_508 = _T_42 ? plru2_22 : _GEN_380; // @[Cache.scala 133:22 137:27]
  wire  _GEN_509 = _T_42 ? plru2_23 : _GEN_381; // @[Cache.scala 133:22 137:27]
  wire  _GEN_510 = _T_42 ? plru2_24 : _GEN_382; // @[Cache.scala 133:22 137:27]
  wire  _GEN_511 = _T_42 ? plru2_25 : _GEN_383; // @[Cache.scala 133:22 137:27]
  wire  _GEN_512 = _T_42 ? plru2_26 : _GEN_384; // @[Cache.scala 133:22 137:27]
  wire  _GEN_513 = _T_42 ? plru2_27 : _GEN_385; // @[Cache.scala 133:22 137:27]
  wire  _GEN_514 = _T_42 ? plru2_28 : _GEN_386; // @[Cache.scala 133:22 137:27]
  wire  _GEN_515 = _T_42 ? plru2_29 : _GEN_387; // @[Cache.scala 133:22 137:27]
  wire  _GEN_516 = _T_42 ? plru2_30 : _GEN_388; // @[Cache.scala 133:22 137:27]
  wire  _GEN_517 = _T_42 ? plru2_31 : _GEN_389; // @[Cache.scala 133:22 137:27]
  wire  _GEN_518 = _T_42 ? plru2_32 : _GEN_390; // @[Cache.scala 133:22 137:27]
  wire  _GEN_519 = _T_42 ? plru2_33 : _GEN_391; // @[Cache.scala 133:22 137:27]
  wire  _GEN_520 = _T_42 ? plru2_34 : _GEN_392; // @[Cache.scala 133:22 137:27]
  wire  _GEN_521 = _T_42 ? plru2_35 : _GEN_393; // @[Cache.scala 133:22 137:27]
  wire  _GEN_522 = _T_42 ? plru2_36 : _GEN_394; // @[Cache.scala 133:22 137:27]
  wire  _GEN_523 = _T_42 ? plru2_37 : _GEN_395; // @[Cache.scala 133:22 137:27]
  wire  _GEN_524 = _T_42 ? plru2_38 : _GEN_396; // @[Cache.scala 133:22 137:27]
  wire  _GEN_525 = _T_42 ? plru2_39 : _GEN_397; // @[Cache.scala 133:22 137:27]
  wire  _GEN_526 = _T_42 ? plru2_40 : _GEN_398; // @[Cache.scala 133:22 137:27]
  wire  _GEN_527 = _T_42 ? plru2_41 : _GEN_399; // @[Cache.scala 133:22 137:27]
  wire  _GEN_528 = _T_42 ? plru2_42 : _GEN_400; // @[Cache.scala 133:22 137:27]
  wire  _GEN_529 = _T_42 ? plru2_43 : _GEN_401; // @[Cache.scala 133:22 137:27]
  wire  _GEN_530 = _T_42 ? plru2_44 : _GEN_402; // @[Cache.scala 133:22 137:27]
  wire  _GEN_531 = _T_42 ? plru2_45 : _GEN_403; // @[Cache.scala 133:22 137:27]
  wire  _GEN_532 = _T_42 ? plru2_46 : _GEN_404; // @[Cache.scala 133:22 137:27]
  wire  _GEN_533 = _T_42 ? plru2_47 : _GEN_405; // @[Cache.scala 133:22 137:27]
  wire  _GEN_534 = _T_42 ? plru2_48 : _GEN_406; // @[Cache.scala 133:22 137:27]
  wire  _GEN_535 = _T_42 ? plru2_49 : _GEN_407; // @[Cache.scala 133:22 137:27]
  wire  _GEN_536 = _T_42 ? plru2_50 : _GEN_408; // @[Cache.scala 133:22 137:27]
  wire  _GEN_537 = _T_42 ? plru2_51 : _GEN_409; // @[Cache.scala 133:22 137:27]
  wire  _GEN_538 = _T_42 ? plru2_52 : _GEN_410; // @[Cache.scala 133:22 137:27]
  wire  _GEN_539 = _T_42 ? plru2_53 : _GEN_411; // @[Cache.scala 133:22 137:27]
  wire  _GEN_540 = _T_42 ? plru2_54 : _GEN_412; // @[Cache.scala 133:22 137:27]
  wire  _GEN_541 = _T_42 ? plru2_55 : _GEN_413; // @[Cache.scala 133:22 137:27]
  wire  _GEN_542 = _T_42 ? plru2_56 : _GEN_414; // @[Cache.scala 133:22 137:27]
  wire  _GEN_543 = _T_42 ? plru2_57 : _GEN_415; // @[Cache.scala 133:22 137:27]
  wire  _GEN_544 = _T_42 ? plru2_58 : _GEN_416; // @[Cache.scala 133:22 137:27]
  wire  _GEN_545 = _T_42 ? plru2_59 : _GEN_417; // @[Cache.scala 133:22 137:27]
  wire  _GEN_546 = _T_42 ? plru2_60 : _GEN_418; // @[Cache.scala 133:22 137:27]
  wire  _GEN_547 = _T_42 ? plru2_61 : _GEN_419; // @[Cache.scala 133:22 137:27]
  wire  _GEN_548 = _T_42 ? plru2_62 : _GEN_420; // @[Cache.scala 133:22 137:27]
  wire  _GEN_549 = _T_42 ? plru2_63 : _GEN_421; // @[Cache.scala 133:22 137:27]
  wire  _T_50 = s2_way == 2'h0; // @[Cache.scala 331:26]
  wire [7:0] _T_62 = s2_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_64 = s2_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_66 = s2_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_68 = s2_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_70 = s2_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_72 = s2_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74 = s2_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76 = s2_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_77 = {_T_76,_T_74,_T_72,_T_70,_T_68,_T_66,_T_64,_T_62}; // @[Cat.scala 30:58]
  wire [63:0] _T_78 = s2_wdata & _T_77; // @[Utils.scala 20:15]
  wire [63:0] _T_79 = ~_T_77; // @[Utils.scala 20:37]
  wire [63:0] _T_80 = _GEN_7[127:64] & _T_79; // @[Utils.scala 20:35]
  wire [63:0] _T_81 = _T_78 | _T_80; // @[Utils.scala 20:23]
  wire [127:0] _T_83 = {_T_81,_GEN_7[63:0]}; // @[Cat.scala 30:58]
  wire [63:0] _T_113 = _GEN_7[63:0] & _T_79; // @[Utils.scala 20:35]
  wire [63:0] _T_114 = _T_78 | _T_113; // @[Utils.scala 20:23]
  wire [127:0] _T_115 = {_GEN_7[127:64],_T_114}; // @[Cat.scala 30:58]
  wire [127:0] _T_116 = s2_offs ? _T_83 : _T_115; // @[Cache.scala 335:38]
  wire  _GEN_742 = s2_way == 2'h0 | pipeline_ready; // @[Cache.scala 331:35 332:29]
  wire [5:0] _GEN_744 = s2_way == 2'h0 ? s2_idx : _GEN_3; // @[Cache.scala 331:35 334:31]
  wire [127:0] _GEN_745 = s2_way == 2'h0 ? _T_116 : 128'h0; // @[Cache.scala 110:16 331:35 335:32]
  wire  _T_117 = s2_way == 2'h1; // @[Cache.scala 331:26]
  wire  _GEN_746 = s2_way == 2'h1 | pipeline_ready; // @[Cache.scala 331:35 332:29]
  wire [5:0] _GEN_748 = s2_way == 2'h1 ? s2_idx : _GEN_3; // @[Cache.scala 331:35 334:31]
  wire [127:0] _GEN_749 = s2_way == 2'h1 ? _T_116 : 128'h0; // @[Cache.scala 110:16 331:35 335:32]
  wire  _T_184 = s2_way == 2'h2; // @[Cache.scala 331:26]
  wire  _GEN_750 = s2_way == 2'h2 | pipeline_ready; // @[Cache.scala 331:35 332:29]
  wire [5:0] _GEN_752 = s2_way == 2'h2 ? s2_idx : _GEN_3; // @[Cache.scala 331:35 334:31]
  wire [127:0] _GEN_753 = s2_way == 2'h2 ? _T_116 : 128'h0; // @[Cache.scala 110:16 331:35 335:32]
  wire  _T_251 = s2_way == 2'h3; // @[Cache.scala 331:26]
  wire  _GEN_754 = s2_way == 2'h3 | pipeline_ready; // @[Cache.scala 331:35 332:29]
  wire [5:0] _GEN_756 = s2_way == 2'h3 ? s2_idx : _GEN_3; // @[Cache.scala 331:35 334:31]
  wire [127:0] _GEN_757 = s2_way == 2'h3 ? _T_116 : 128'h0; // @[Cache.scala 110:16 331:35 335:32]
  wire [3:0] _GEN_758 = ~s2_hit ? 4'h1 : state; // @[Cache.scala 344:31 345:17 213:22]
  wire  _GEN_759 = s2_hit & s2_wen ? _GEN_742 : pipeline_ready; // @[Cache.scala 329:33]
  wire  _GEN_760 = s2_hit & s2_wen & _T_50; // @[Cache.scala 108:14 329:33]
  wire [5:0] _GEN_761 = s2_hit & s2_wen ? _GEN_744 : _GEN_3; // @[Cache.scala 329:33]
  wire [127:0] _GEN_762 = s2_hit & s2_wen ? _GEN_745 : 128'h0; // @[Cache.scala 110:16 329:33]
  wire  _GEN_763 = s2_hit & s2_wen ? _GEN_746 : pipeline_ready; // @[Cache.scala 329:33]
  wire  _GEN_764 = s2_hit & s2_wen & _T_117; // @[Cache.scala 108:14 329:33]
  wire [5:0] _GEN_765 = s2_hit & s2_wen ? _GEN_748 : _GEN_3; // @[Cache.scala 329:33]
  wire [127:0] _GEN_766 = s2_hit & s2_wen ? _GEN_749 : 128'h0; // @[Cache.scala 110:16 329:33]
  wire  _GEN_767 = s2_hit & s2_wen ? _GEN_750 : pipeline_ready; // @[Cache.scala 329:33]
  wire  _GEN_768 = s2_hit & s2_wen & _T_184; // @[Cache.scala 108:14 329:33]
  wire [5:0] _GEN_769 = s2_hit & s2_wen ? _GEN_752 : _GEN_3; // @[Cache.scala 329:33]
  wire [127:0] _GEN_770 = s2_hit & s2_wen ? _GEN_753 : 128'h0; // @[Cache.scala 110:16 329:33]
  wire  _GEN_771 = s2_hit & s2_wen ? _GEN_754 : pipeline_ready; // @[Cache.scala 329:33]
  wire  _GEN_772 = s2_hit & s2_wen & _T_251; // @[Cache.scala 108:14 329:33]
  wire [5:0] _GEN_773 = s2_hit & s2_wen ? _GEN_756 : _GEN_3; // @[Cache.scala 329:33]
  wire [127:0] _GEN_774 = s2_hit & s2_wen ? _GEN_757 : 128'h0; // @[Cache.scala 110:16 329:33]
  wire [3:0] _GEN_775 = s2_hit & s2_wen ? 4'h7 : _GEN_758; // @[Cache.scala 329:33 343:17]
  wire  _GEN_968 = REG_11 ? _GEN_759 : pipeline_ready; // @[Cache.scala 325:37]
  wire  _GEN_969 = REG_11 & _GEN_760; // @[Cache.scala 108:14 325:37]
  wire [5:0] _GEN_970 = REG_11 ? _GEN_761 : _GEN_3; // @[Cache.scala 325:37]
  wire [127:0] _GEN_971 = REG_11 ? _GEN_762 : 128'h0; // @[Cache.scala 110:16 325:37]
  wire  _GEN_972 = REG_11 ? _GEN_763 : pipeline_ready; // @[Cache.scala 325:37]
  wire  _GEN_973 = REG_11 & _GEN_764; // @[Cache.scala 108:14 325:37]
  wire [5:0] _GEN_974 = REG_11 ? _GEN_765 : _GEN_3; // @[Cache.scala 325:37]
  wire [127:0] _GEN_975 = REG_11 ? _GEN_766 : 128'h0; // @[Cache.scala 110:16 325:37]
  wire  _GEN_976 = REG_11 ? _GEN_767 : pipeline_ready; // @[Cache.scala 325:37]
  wire  _GEN_977 = REG_11 & _GEN_768; // @[Cache.scala 108:14 325:37]
  wire [5:0] _GEN_978 = REG_11 ? _GEN_769 : _GEN_3; // @[Cache.scala 325:37]
  wire [127:0] _GEN_979 = REG_11 ? _GEN_770 : 128'h0; // @[Cache.scala 110:16 325:37]
  wire  _GEN_980 = REG_11 ? _GEN_771 : pipeline_ready; // @[Cache.scala 325:37]
  wire  _GEN_981 = REG_11 & _GEN_772; // @[Cache.scala 108:14 325:37]
  wire [5:0] _GEN_982 = REG_11 ? _GEN_773 : _GEN_3; // @[Cache.scala 325:37]
  wire [127:0] _GEN_983 = REG_11 ? _GEN_774 : 128'h0; // @[Cache.scala 110:16 325:37]
  wire [3:0] _GEN_984 = REG_11 ? _GEN_775 : state; // @[Cache.scala 213:22 325:37]
  wire  _T_320 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_985 = _T_320 ? 4'h2 : state; // @[Cache.scala 350:29 351:15 213:22]
  wire  _T_322 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_986 = ~io_out_resp_bits_rlast ? io_out_resp_bits_rdata : wdata1; // @[Cache.scala 356:37 357:18 270:23]
  wire [63:0] _GEN_987 = ~io_out_resp_bits_rlast ? wdata2 : io_out_resp_bits_rdata; // @[Cache.scala 271:23 356:37 359:18]
  wire [3:0] _GEN_988 = ~io_out_resp_bits_rlast ? state : 4'h3; // @[Cache.scala 213:22 356:37 360:17]
  wire [63:0] _GEN_989 = _T_322 ? _GEN_986 : wdata1; // @[Cache.scala 270:23 355:30]
  wire [63:0] _GEN_990 = _T_322 ? _GEN_987 : wdata2; // @[Cache.scala 271:23 355:30]
  wire [3:0] _GEN_991 = _T_322 ? _GEN_988 : state; // @[Cache.scala 213:22 355:30]
  wire  _T_325 = replace_way == 2'h0; // @[Cache.scala 366:27]
  wire [63:0] _T_354 = wdata2 & _T_79; // @[Utils.scala 20:35]
  wire [63:0] _T_355 = _T_78 | _T_354; // @[Utils.scala 20:23]
  wire [127:0] _T_356 = {_T_355,wdata1}; // @[Cat.scala 30:58]
  wire [63:0] _T_384 = wdata1 & _T_79; // @[Utils.scala 20:35]
  wire [63:0] _T_385 = _T_78 | _T_384; // @[Utils.scala 20:23]
  wire [127:0] _T_386 = {wdata2,_T_385}; // @[Cat.scala 30:58]
  wire [127:0] _T_387 = s2_offs ? _T_356 : _T_386; // @[Cache.scala 371:36]
  wire [127:0] _T_388 = {wdata2,wdata1}; // @[Cat.scala 30:58]
  wire [127:0] _GEN_992 = s2_wen ? _T_387 : _T_388; // @[Cache.scala 370:25 371:30 375:30]
  wire  _GEN_993 = replace_way == 2'h0 | pipeline_ready; // @[Cache.scala 366:36 367:25]
  wire [5:0] _GEN_995 = replace_way == 2'h0 ? s2_idx : _GEN_3; // @[Cache.scala 366:36 369:27]
  wire [127:0] _GEN_996 = replace_way == 2'h0 ? _GEN_992 : 128'h0; // @[Cache.scala 110:16 366:36]
  wire [20:0] _GEN_997 = replace_way == 2'h0 ? s2_tag : 21'h0; // @[Cache.scala 114:16 366:36 380:28]
  wire  _GEN_998 = replace_way == 2'h0 & s2_wen; // @[Cache.scala 116:18 366:36 382:30]
  wire  _T_389 = replace_way == 2'h1; // @[Cache.scala 366:27]
  wire  _GEN_1000 = replace_way == 2'h1 | pipeline_ready; // @[Cache.scala 366:36 367:25]
  wire [5:0] _GEN_1002 = replace_way == 2'h1 ? s2_idx : _GEN_3; // @[Cache.scala 366:36 369:27]
  wire [127:0] _GEN_1003 = replace_way == 2'h1 ? _GEN_992 : 128'h0; // @[Cache.scala 110:16 366:36]
  wire [20:0] _GEN_1004 = replace_way == 2'h1 ? s2_tag : 21'h0; // @[Cache.scala 114:16 366:36 380:28]
  wire  _GEN_1005 = replace_way == 2'h1 & s2_wen; // @[Cache.scala 116:18 366:36 382:30]
  wire  _T_453 = replace_way == 2'h2; // @[Cache.scala 366:27]
  wire  _GEN_1007 = replace_way == 2'h2 | pipeline_ready; // @[Cache.scala 366:36 367:25]
  wire [5:0] _GEN_1009 = replace_way == 2'h2 ? s2_idx : _GEN_3; // @[Cache.scala 366:36 369:27]
  wire [127:0] _GEN_1010 = replace_way == 2'h2 ? _GEN_992 : 128'h0; // @[Cache.scala 110:16 366:36]
  wire [20:0] _GEN_1011 = replace_way == 2'h2 ? s2_tag : 21'h0; // @[Cache.scala 114:16 366:36 380:28]
  wire  _GEN_1012 = replace_way == 2'h2 & s2_wen; // @[Cache.scala 116:18 366:36 382:30]
  wire  _T_517 = replace_way == 2'h3; // @[Cache.scala 366:27]
  wire  _GEN_1014 = replace_way == 2'h3 | pipeline_ready; // @[Cache.scala 366:36 367:25]
  wire [5:0] _GEN_1016 = replace_way == 2'h3 ? s2_idx : _GEN_3; // @[Cache.scala 366:36 369:27]
  wire [127:0] _GEN_1017 = replace_way == 2'h3 ? _GEN_992 : 128'h0; // @[Cache.scala 110:16 366:36]
  wire [20:0] _GEN_1018 = replace_way == 2'h3 ? s2_tag : 21'h0; // @[Cache.scala 114:16 366:36 380:28]
  wire  _GEN_1019 = replace_way == 2'h3 & s2_wen; // @[Cache.scala 116:18 366:36 382:30]
  wire  _T_582 = ~replace_way[1]; // @[Cache.scala 136:19]
  wire  _GEN_1020 = 6'h0 == s2_idx ? ~replace_way[1] : plru0_0; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1021 = 6'h1 == s2_idx ? ~replace_way[1] : plru0_1; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1022 = 6'h2 == s2_idx ? ~replace_way[1] : plru0_2; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1023 = 6'h3 == s2_idx ? ~replace_way[1] : plru0_3; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1024 = 6'h4 == s2_idx ? ~replace_way[1] : plru0_4; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1025 = 6'h5 == s2_idx ? ~replace_way[1] : plru0_5; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1026 = 6'h6 == s2_idx ? ~replace_way[1] : plru0_6; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1027 = 6'h7 == s2_idx ? ~replace_way[1] : plru0_7; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1028 = 6'h8 == s2_idx ? ~replace_way[1] : plru0_8; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1029 = 6'h9 == s2_idx ? ~replace_way[1] : plru0_9; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1030 = 6'ha == s2_idx ? ~replace_way[1] : plru0_10; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1031 = 6'hb == s2_idx ? ~replace_way[1] : plru0_11; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1032 = 6'hc == s2_idx ? ~replace_way[1] : plru0_12; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1033 = 6'hd == s2_idx ? ~replace_way[1] : plru0_13; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1034 = 6'he == s2_idx ? ~replace_way[1] : plru0_14; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1035 = 6'hf == s2_idx ? ~replace_way[1] : plru0_15; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1036 = 6'h10 == s2_idx ? ~replace_way[1] : plru0_16; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1037 = 6'h11 == s2_idx ? ~replace_way[1] : plru0_17; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1038 = 6'h12 == s2_idx ? ~replace_way[1] : plru0_18; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1039 = 6'h13 == s2_idx ? ~replace_way[1] : plru0_19; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1040 = 6'h14 == s2_idx ? ~replace_way[1] : plru0_20; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1041 = 6'h15 == s2_idx ? ~replace_way[1] : plru0_21; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1042 = 6'h16 == s2_idx ? ~replace_way[1] : plru0_22; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1043 = 6'h17 == s2_idx ? ~replace_way[1] : plru0_23; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1044 = 6'h18 == s2_idx ? ~replace_way[1] : plru0_24; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1045 = 6'h19 == s2_idx ? ~replace_way[1] : plru0_25; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1046 = 6'h1a == s2_idx ? ~replace_way[1] : plru0_26; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1047 = 6'h1b == s2_idx ? ~replace_way[1] : plru0_27; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1048 = 6'h1c == s2_idx ? ~replace_way[1] : plru0_28; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1049 = 6'h1d == s2_idx ? ~replace_way[1] : plru0_29; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1050 = 6'h1e == s2_idx ? ~replace_way[1] : plru0_30; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1051 = 6'h1f == s2_idx ? ~replace_way[1] : plru0_31; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1052 = 6'h20 == s2_idx ? ~replace_way[1] : plru0_32; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1053 = 6'h21 == s2_idx ? ~replace_way[1] : plru0_33; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1054 = 6'h22 == s2_idx ? ~replace_way[1] : plru0_34; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1055 = 6'h23 == s2_idx ? ~replace_way[1] : plru0_35; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1056 = 6'h24 == s2_idx ? ~replace_way[1] : plru0_36; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1057 = 6'h25 == s2_idx ? ~replace_way[1] : plru0_37; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1058 = 6'h26 == s2_idx ? ~replace_way[1] : plru0_38; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1059 = 6'h27 == s2_idx ? ~replace_way[1] : plru0_39; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1060 = 6'h28 == s2_idx ? ~replace_way[1] : plru0_40; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1061 = 6'h29 == s2_idx ? ~replace_way[1] : plru0_41; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1062 = 6'h2a == s2_idx ? ~replace_way[1] : plru0_42; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1063 = 6'h2b == s2_idx ? ~replace_way[1] : plru0_43; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1064 = 6'h2c == s2_idx ? ~replace_way[1] : plru0_44; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1065 = 6'h2d == s2_idx ? ~replace_way[1] : plru0_45; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1066 = 6'h2e == s2_idx ? ~replace_way[1] : plru0_46; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1067 = 6'h2f == s2_idx ? ~replace_way[1] : plru0_47; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1068 = 6'h30 == s2_idx ? ~replace_way[1] : plru0_48; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1069 = 6'h31 == s2_idx ? ~replace_way[1] : plru0_49; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1070 = 6'h32 == s2_idx ? ~replace_way[1] : plru0_50; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1071 = 6'h33 == s2_idx ? ~replace_way[1] : plru0_51; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1072 = 6'h34 == s2_idx ? ~replace_way[1] : plru0_52; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1073 = 6'h35 == s2_idx ? ~replace_way[1] : plru0_53; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1074 = 6'h36 == s2_idx ? ~replace_way[1] : plru0_54; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1075 = 6'h37 == s2_idx ? ~replace_way[1] : plru0_55; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1076 = 6'h38 == s2_idx ? ~replace_way[1] : plru0_56; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1077 = 6'h39 == s2_idx ? ~replace_way[1] : plru0_57; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1078 = 6'h3a == s2_idx ? ~replace_way[1] : plru0_58; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1079 = 6'h3b == s2_idx ? ~replace_way[1] : plru0_59; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1080 = 6'h3c == s2_idx ? ~replace_way[1] : plru0_60; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1081 = 6'h3d == s2_idx ? ~replace_way[1] : plru0_61; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1082 = 6'h3e == s2_idx ? ~replace_way[1] : plru0_62; // @[Cache.scala 136:{16,16} 129:22]
  wire  _GEN_1083 = 6'h3f == s2_idx ? ~replace_way[1] : plru0_63; // @[Cache.scala 136:{16,16} 129:22]
  wire  _T_586 = ~replace_way[0]; // @[Cache.scala 138:21]
  wire  _GEN_1084 = 6'h0 == s2_idx ? ~replace_way[0] : plru1_0; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1085 = 6'h1 == s2_idx ? ~replace_way[0] : plru1_1; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1086 = 6'h2 == s2_idx ? ~replace_way[0] : plru1_2; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1087 = 6'h3 == s2_idx ? ~replace_way[0] : plru1_3; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1088 = 6'h4 == s2_idx ? ~replace_way[0] : plru1_4; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1089 = 6'h5 == s2_idx ? ~replace_way[0] : plru1_5; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1090 = 6'h6 == s2_idx ? ~replace_way[0] : plru1_6; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1091 = 6'h7 == s2_idx ? ~replace_way[0] : plru1_7; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1092 = 6'h8 == s2_idx ? ~replace_way[0] : plru1_8; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1093 = 6'h9 == s2_idx ? ~replace_way[0] : plru1_9; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1094 = 6'ha == s2_idx ? ~replace_way[0] : plru1_10; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1095 = 6'hb == s2_idx ? ~replace_way[0] : plru1_11; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1096 = 6'hc == s2_idx ? ~replace_way[0] : plru1_12; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1097 = 6'hd == s2_idx ? ~replace_way[0] : plru1_13; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1098 = 6'he == s2_idx ? ~replace_way[0] : plru1_14; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1099 = 6'hf == s2_idx ? ~replace_way[0] : plru1_15; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1100 = 6'h10 == s2_idx ? ~replace_way[0] : plru1_16; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1101 = 6'h11 == s2_idx ? ~replace_way[0] : plru1_17; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1102 = 6'h12 == s2_idx ? ~replace_way[0] : plru1_18; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1103 = 6'h13 == s2_idx ? ~replace_way[0] : plru1_19; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1104 = 6'h14 == s2_idx ? ~replace_way[0] : plru1_20; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1105 = 6'h15 == s2_idx ? ~replace_way[0] : plru1_21; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1106 = 6'h16 == s2_idx ? ~replace_way[0] : plru1_22; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1107 = 6'h17 == s2_idx ? ~replace_way[0] : plru1_23; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1108 = 6'h18 == s2_idx ? ~replace_way[0] : plru1_24; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1109 = 6'h19 == s2_idx ? ~replace_way[0] : plru1_25; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1110 = 6'h1a == s2_idx ? ~replace_way[0] : plru1_26; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1111 = 6'h1b == s2_idx ? ~replace_way[0] : plru1_27; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1112 = 6'h1c == s2_idx ? ~replace_way[0] : plru1_28; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1113 = 6'h1d == s2_idx ? ~replace_way[0] : plru1_29; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1114 = 6'h1e == s2_idx ? ~replace_way[0] : plru1_30; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1115 = 6'h1f == s2_idx ? ~replace_way[0] : plru1_31; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1116 = 6'h20 == s2_idx ? ~replace_way[0] : plru1_32; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1117 = 6'h21 == s2_idx ? ~replace_way[0] : plru1_33; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1118 = 6'h22 == s2_idx ? ~replace_way[0] : plru1_34; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1119 = 6'h23 == s2_idx ? ~replace_way[0] : plru1_35; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1120 = 6'h24 == s2_idx ? ~replace_way[0] : plru1_36; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1121 = 6'h25 == s2_idx ? ~replace_way[0] : plru1_37; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1122 = 6'h26 == s2_idx ? ~replace_way[0] : plru1_38; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1123 = 6'h27 == s2_idx ? ~replace_way[0] : plru1_39; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1124 = 6'h28 == s2_idx ? ~replace_way[0] : plru1_40; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1125 = 6'h29 == s2_idx ? ~replace_way[0] : plru1_41; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1126 = 6'h2a == s2_idx ? ~replace_way[0] : plru1_42; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1127 = 6'h2b == s2_idx ? ~replace_way[0] : plru1_43; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1128 = 6'h2c == s2_idx ? ~replace_way[0] : plru1_44; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1129 = 6'h2d == s2_idx ? ~replace_way[0] : plru1_45; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1130 = 6'h2e == s2_idx ? ~replace_way[0] : plru1_46; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1131 = 6'h2f == s2_idx ? ~replace_way[0] : plru1_47; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1132 = 6'h30 == s2_idx ? ~replace_way[0] : plru1_48; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1133 = 6'h31 == s2_idx ? ~replace_way[0] : plru1_49; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1134 = 6'h32 == s2_idx ? ~replace_way[0] : plru1_50; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1135 = 6'h33 == s2_idx ? ~replace_way[0] : plru1_51; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1136 = 6'h34 == s2_idx ? ~replace_way[0] : plru1_52; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1137 = 6'h35 == s2_idx ? ~replace_way[0] : plru1_53; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1138 = 6'h36 == s2_idx ? ~replace_way[0] : plru1_54; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1139 = 6'h37 == s2_idx ? ~replace_way[0] : plru1_55; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1140 = 6'h38 == s2_idx ? ~replace_way[0] : plru1_56; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1141 = 6'h39 == s2_idx ? ~replace_way[0] : plru1_57; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1142 = 6'h3a == s2_idx ? ~replace_way[0] : plru1_58; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1143 = 6'h3b == s2_idx ? ~replace_way[0] : plru1_59; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1144 = 6'h3c == s2_idx ? ~replace_way[0] : plru1_60; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1145 = 6'h3d == s2_idx ? ~replace_way[0] : plru1_61; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1146 = 6'h3e == s2_idx ? ~replace_way[0] : plru1_62; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1147 = 6'h3f == s2_idx ? ~replace_way[0] : plru1_63; // @[Cache.scala 138:{18,18} 131:22]
  wire  _GEN_1148 = 6'h0 == s2_idx ? _T_586 : plru2_0; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1149 = 6'h1 == s2_idx ? _T_586 : plru2_1; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1150 = 6'h2 == s2_idx ? _T_586 : plru2_2; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1151 = 6'h3 == s2_idx ? _T_586 : plru2_3; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1152 = 6'h4 == s2_idx ? _T_586 : plru2_4; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1153 = 6'h5 == s2_idx ? _T_586 : plru2_5; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1154 = 6'h6 == s2_idx ? _T_586 : plru2_6; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1155 = 6'h7 == s2_idx ? _T_586 : plru2_7; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1156 = 6'h8 == s2_idx ? _T_586 : plru2_8; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1157 = 6'h9 == s2_idx ? _T_586 : plru2_9; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1158 = 6'ha == s2_idx ? _T_586 : plru2_10; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1159 = 6'hb == s2_idx ? _T_586 : plru2_11; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1160 = 6'hc == s2_idx ? _T_586 : plru2_12; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1161 = 6'hd == s2_idx ? _T_586 : plru2_13; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1162 = 6'he == s2_idx ? _T_586 : plru2_14; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1163 = 6'hf == s2_idx ? _T_586 : plru2_15; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1164 = 6'h10 == s2_idx ? _T_586 : plru2_16; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1165 = 6'h11 == s2_idx ? _T_586 : plru2_17; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1166 = 6'h12 == s2_idx ? _T_586 : plru2_18; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1167 = 6'h13 == s2_idx ? _T_586 : plru2_19; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1168 = 6'h14 == s2_idx ? _T_586 : plru2_20; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1169 = 6'h15 == s2_idx ? _T_586 : plru2_21; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1170 = 6'h16 == s2_idx ? _T_586 : plru2_22; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1171 = 6'h17 == s2_idx ? _T_586 : plru2_23; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1172 = 6'h18 == s2_idx ? _T_586 : plru2_24; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1173 = 6'h19 == s2_idx ? _T_586 : plru2_25; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1174 = 6'h1a == s2_idx ? _T_586 : plru2_26; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1175 = 6'h1b == s2_idx ? _T_586 : plru2_27; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1176 = 6'h1c == s2_idx ? _T_586 : plru2_28; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1177 = 6'h1d == s2_idx ? _T_586 : plru2_29; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1178 = 6'h1e == s2_idx ? _T_586 : plru2_30; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1179 = 6'h1f == s2_idx ? _T_586 : plru2_31; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1180 = 6'h20 == s2_idx ? _T_586 : plru2_32; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1181 = 6'h21 == s2_idx ? _T_586 : plru2_33; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1182 = 6'h22 == s2_idx ? _T_586 : plru2_34; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1183 = 6'h23 == s2_idx ? _T_586 : plru2_35; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1184 = 6'h24 == s2_idx ? _T_586 : plru2_36; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1185 = 6'h25 == s2_idx ? _T_586 : plru2_37; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1186 = 6'h26 == s2_idx ? _T_586 : plru2_38; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1187 = 6'h27 == s2_idx ? _T_586 : plru2_39; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1188 = 6'h28 == s2_idx ? _T_586 : plru2_40; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1189 = 6'h29 == s2_idx ? _T_586 : plru2_41; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1190 = 6'h2a == s2_idx ? _T_586 : plru2_42; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1191 = 6'h2b == s2_idx ? _T_586 : plru2_43; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1192 = 6'h2c == s2_idx ? _T_586 : plru2_44; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1193 = 6'h2d == s2_idx ? _T_586 : plru2_45; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1194 = 6'h2e == s2_idx ? _T_586 : plru2_46; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1195 = 6'h2f == s2_idx ? _T_586 : plru2_47; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1196 = 6'h30 == s2_idx ? _T_586 : plru2_48; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1197 = 6'h31 == s2_idx ? _T_586 : plru2_49; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1198 = 6'h32 == s2_idx ? _T_586 : plru2_50; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1199 = 6'h33 == s2_idx ? _T_586 : plru2_51; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1200 = 6'h34 == s2_idx ? _T_586 : plru2_52; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1201 = 6'h35 == s2_idx ? _T_586 : plru2_53; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1202 = 6'h36 == s2_idx ? _T_586 : plru2_54; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1203 = 6'h37 == s2_idx ? _T_586 : plru2_55; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1204 = 6'h38 == s2_idx ? _T_586 : plru2_56; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1205 = 6'h39 == s2_idx ? _T_586 : plru2_57; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1206 = 6'h3a == s2_idx ? _T_586 : plru2_58; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1207 = 6'h3b == s2_idx ? _T_586 : plru2_59; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1208 = 6'h3c == s2_idx ? _T_586 : plru2_60; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1209 = 6'h3d == s2_idx ? _T_586 : plru2_61; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1210 = 6'h3e == s2_idx ? _T_586 : plru2_62; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1211 = 6'h3f == s2_idx ? _T_586 : plru2_63; // @[Cache.scala 140:{18,18} 133:22]
  wire  _GEN_1212 = _T_582 ? _GEN_1084 : plru1_0; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1213 = _T_582 ? _GEN_1085 : plru1_1; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1214 = _T_582 ? _GEN_1086 : plru1_2; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1215 = _T_582 ? _GEN_1087 : plru1_3; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1216 = _T_582 ? _GEN_1088 : plru1_4; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1217 = _T_582 ? _GEN_1089 : plru1_5; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1218 = _T_582 ? _GEN_1090 : plru1_6; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1219 = _T_582 ? _GEN_1091 : plru1_7; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1220 = _T_582 ? _GEN_1092 : plru1_8; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1221 = _T_582 ? _GEN_1093 : plru1_9; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1222 = _T_582 ? _GEN_1094 : plru1_10; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1223 = _T_582 ? _GEN_1095 : plru1_11; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1224 = _T_582 ? _GEN_1096 : plru1_12; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1225 = _T_582 ? _GEN_1097 : plru1_13; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1226 = _T_582 ? _GEN_1098 : plru1_14; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1227 = _T_582 ? _GEN_1099 : plru1_15; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1228 = _T_582 ? _GEN_1100 : plru1_16; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1229 = _T_582 ? _GEN_1101 : plru1_17; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1230 = _T_582 ? _GEN_1102 : plru1_18; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1231 = _T_582 ? _GEN_1103 : plru1_19; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1232 = _T_582 ? _GEN_1104 : plru1_20; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1233 = _T_582 ? _GEN_1105 : plru1_21; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1234 = _T_582 ? _GEN_1106 : plru1_22; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1235 = _T_582 ? _GEN_1107 : plru1_23; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1236 = _T_582 ? _GEN_1108 : plru1_24; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1237 = _T_582 ? _GEN_1109 : plru1_25; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1238 = _T_582 ? _GEN_1110 : plru1_26; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1239 = _T_582 ? _GEN_1111 : plru1_27; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1240 = _T_582 ? _GEN_1112 : plru1_28; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1241 = _T_582 ? _GEN_1113 : plru1_29; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1242 = _T_582 ? _GEN_1114 : plru1_30; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1243 = _T_582 ? _GEN_1115 : plru1_31; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1244 = _T_582 ? _GEN_1116 : plru1_32; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1245 = _T_582 ? _GEN_1117 : plru1_33; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1246 = _T_582 ? _GEN_1118 : plru1_34; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1247 = _T_582 ? _GEN_1119 : plru1_35; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1248 = _T_582 ? _GEN_1120 : plru1_36; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1249 = _T_582 ? _GEN_1121 : plru1_37; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1250 = _T_582 ? _GEN_1122 : plru1_38; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1251 = _T_582 ? _GEN_1123 : plru1_39; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1252 = _T_582 ? _GEN_1124 : plru1_40; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1253 = _T_582 ? _GEN_1125 : plru1_41; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1254 = _T_582 ? _GEN_1126 : plru1_42; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1255 = _T_582 ? _GEN_1127 : plru1_43; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1256 = _T_582 ? _GEN_1128 : plru1_44; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1257 = _T_582 ? _GEN_1129 : plru1_45; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1258 = _T_582 ? _GEN_1130 : plru1_46; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1259 = _T_582 ? _GEN_1131 : plru1_47; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1260 = _T_582 ? _GEN_1132 : plru1_48; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1261 = _T_582 ? _GEN_1133 : plru1_49; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1262 = _T_582 ? _GEN_1134 : plru1_50; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1263 = _T_582 ? _GEN_1135 : plru1_51; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1264 = _T_582 ? _GEN_1136 : plru1_52; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1265 = _T_582 ? _GEN_1137 : plru1_53; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1266 = _T_582 ? _GEN_1138 : plru1_54; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1267 = _T_582 ? _GEN_1139 : plru1_55; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1268 = _T_582 ? _GEN_1140 : plru1_56; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1269 = _T_582 ? _GEN_1141 : plru1_57; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1270 = _T_582 ? _GEN_1142 : plru1_58; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1271 = _T_582 ? _GEN_1143 : plru1_59; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1272 = _T_582 ? _GEN_1144 : plru1_60; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1273 = _T_582 ? _GEN_1145 : plru1_61; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1274 = _T_582 ? _GEN_1146 : plru1_62; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1275 = _T_582 ? _GEN_1147 : plru1_63; // @[Cache.scala 131:22 137:27]
  wire  _GEN_1276 = _T_582 ? plru2_0 : _GEN_1148; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1277 = _T_582 ? plru2_1 : _GEN_1149; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1278 = _T_582 ? plru2_2 : _GEN_1150; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1279 = _T_582 ? plru2_3 : _GEN_1151; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1280 = _T_582 ? plru2_4 : _GEN_1152; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1281 = _T_582 ? plru2_5 : _GEN_1153; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1282 = _T_582 ? plru2_6 : _GEN_1154; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1283 = _T_582 ? plru2_7 : _GEN_1155; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1284 = _T_582 ? plru2_8 : _GEN_1156; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1285 = _T_582 ? plru2_9 : _GEN_1157; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1286 = _T_582 ? plru2_10 : _GEN_1158; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1287 = _T_582 ? plru2_11 : _GEN_1159; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1288 = _T_582 ? plru2_12 : _GEN_1160; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1289 = _T_582 ? plru2_13 : _GEN_1161; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1290 = _T_582 ? plru2_14 : _GEN_1162; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1291 = _T_582 ? plru2_15 : _GEN_1163; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1292 = _T_582 ? plru2_16 : _GEN_1164; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1293 = _T_582 ? plru2_17 : _GEN_1165; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1294 = _T_582 ? plru2_18 : _GEN_1166; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1295 = _T_582 ? plru2_19 : _GEN_1167; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1296 = _T_582 ? plru2_20 : _GEN_1168; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1297 = _T_582 ? plru2_21 : _GEN_1169; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1298 = _T_582 ? plru2_22 : _GEN_1170; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1299 = _T_582 ? plru2_23 : _GEN_1171; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1300 = _T_582 ? plru2_24 : _GEN_1172; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1301 = _T_582 ? plru2_25 : _GEN_1173; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1302 = _T_582 ? plru2_26 : _GEN_1174; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1303 = _T_582 ? plru2_27 : _GEN_1175; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1304 = _T_582 ? plru2_28 : _GEN_1176; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1305 = _T_582 ? plru2_29 : _GEN_1177; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1306 = _T_582 ? plru2_30 : _GEN_1178; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1307 = _T_582 ? plru2_31 : _GEN_1179; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1308 = _T_582 ? plru2_32 : _GEN_1180; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1309 = _T_582 ? plru2_33 : _GEN_1181; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1310 = _T_582 ? plru2_34 : _GEN_1182; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1311 = _T_582 ? plru2_35 : _GEN_1183; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1312 = _T_582 ? plru2_36 : _GEN_1184; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1313 = _T_582 ? plru2_37 : _GEN_1185; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1314 = _T_582 ? plru2_38 : _GEN_1186; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1315 = _T_582 ? plru2_39 : _GEN_1187; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1316 = _T_582 ? plru2_40 : _GEN_1188; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1317 = _T_582 ? plru2_41 : _GEN_1189; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1318 = _T_582 ? plru2_42 : _GEN_1190; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1319 = _T_582 ? plru2_43 : _GEN_1191; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1320 = _T_582 ? plru2_44 : _GEN_1192; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1321 = _T_582 ? plru2_45 : _GEN_1193; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1322 = _T_582 ? plru2_46 : _GEN_1194; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1323 = _T_582 ? plru2_47 : _GEN_1195; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1324 = _T_582 ? plru2_48 : _GEN_1196; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1325 = _T_582 ? plru2_49 : _GEN_1197; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1326 = _T_582 ? plru2_50 : _GEN_1198; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1327 = _T_582 ? plru2_51 : _GEN_1199; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1328 = _T_582 ? plru2_52 : _GEN_1200; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1329 = _T_582 ? plru2_53 : _GEN_1201; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1330 = _T_582 ? plru2_54 : _GEN_1202; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1331 = _T_582 ? plru2_55 : _GEN_1203; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1332 = _T_582 ? plru2_56 : _GEN_1204; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1333 = _T_582 ? plru2_57 : _GEN_1205; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1334 = _T_582 ? plru2_58 : _GEN_1206; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1335 = _T_582 ? plru2_59 : _GEN_1207; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1336 = _T_582 ? plru2_60 : _GEN_1208; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1337 = _T_582 ? plru2_61 : _GEN_1209; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1338 = _T_582 ? plru2_62 : _GEN_1210; // @[Cache.scala 133:22 137:27]
  wire  _GEN_1339 = _T_582 ? plru2_63 : _GEN_1211; // @[Cache.scala 133:22 137:27]
  wire [3:0] _GEN_1340 = s2_reg_dirty ? 4'h4 : 4'h7; // @[Cache.scala 385:27 386:15 389:15]
  wire  _GEN_1341 = s2_reg_dirty ? plru0_0 : _GEN_1020; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1342 = s2_reg_dirty ? plru0_1 : _GEN_1021; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1343 = s2_reg_dirty ? plru0_2 : _GEN_1022; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1344 = s2_reg_dirty ? plru0_3 : _GEN_1023; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1345 = s2_reg_dirty ? plru0_4 : _GEN_1024; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1346 = s2_reg_dirty ? plru0_5 : _GEN_1025; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1347 = s2_reg_dirty ? plru0_6 : _GEN_1026; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1348 = s2_reg_dirty ? plru0_7 : _GEN_1027; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1349 = s2_reg_dirty ? plru0_8 : _GEN_1028; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1350 = s2_reg_dirty ? plru0_9 : _GEN_1029; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1351 = s2_reg_dirty ? plru0_10 : _GEN_1030; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1352 = s2_reg_dirty ? plru0_11 : _GEN_1031; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1353 = s2_reg_dirty ? plru0_12 : _GEN_1032; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1354 = s2_reg_dirty ? plru0_13 : _GEN_1033; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1355 = s2_reg_dirty ? plru0_14 : _GEN_1034; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1356 = s2_reg_dirty ? plru0_15 : _GEN_1035; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1357 = s2_reg_dirty ? plru0_16 : _GEN_1036; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1358 = s2_reg_dirty ? plru0_17 : _GEN_1037; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1359 = s2_reg_dirty ? plru0_18 : _GEN_1038; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1360 = s2_reg_dirty ? plru0_19 : _GEN_1039; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1361 = s2_reg_dirty ? plru0_20 : _GEN_1040; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1362 = s2_reg_dirty ? plru0_21 : _GEN_1041; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1363 = s2_reg_dirty ? plru0_22 : _GEN_1042; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1364 = s2_reg_dirty ? plru0_23 : _GEN_1043; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1365 = s2_reg_dirty ? plru0_24 : _GEN_1044; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1366 = s2_reg_dirty ? plru0_25 : _GEN_1045; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1367 = s2_reg_dirty ? plru0_26 : _GEN_1046; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1368 = s2_reg_dirty ? plru0_27 : _GEN_1047; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1369 = s2_reg_dirty ? plru0_28 : _GEN_1048; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1370 = s2_reg_dirty ? plru0_29 : _GEN_1049; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1371 = s2_reg_dirty ? plru0_30 : _GEN_1050; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1372 = s2_reg_dirty ? plru0_31 : _GEN_1051; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1373 = s2_reg_dirty ? plru0_32 : _GEN_1052; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1374 = s2_reg_dirty ? plru0_33 : _GEN_1053; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1375 = s2_reg_dirty ? plru0_34 : _GEN_1054; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1376 = s2_reg_dirty ? plru0_35 : _GEN_1055; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1377 = s2_reg_dirty ? plru0_36 : _GEN_1056; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1378 = s2_reg_dirty ? plru0_37 : _GEN_1057; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1379 = s2_reg_dirty ? plru0_38 : _GEN_1058; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1380 = s2_reg_dirty ? plru0_39 : _GEN_1059; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1381 = s2_reg_dirty ? plru0_40 : _GEN_1060; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1382 = s2_reg_dirty ? plru0_41 : _GEN_1061; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1383 = s2_reg_dirty ? plru0_42 : _GEN_1062; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1384 = s2_reg_dirty ? plru0_43 : _GEN_1063; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1385 = s2_reg_dirty ? plru0_44 : _GEN_1064; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1386 = s2_reg_dirty ? plru0_45 : _GEN_1065; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1387 = s2_reg_dirty ? plru0_46 : _GEN_1066; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1388 = s2_reg_dirty ? plru0_47 : _GEN_1067; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1389 = s2_reg_dirty ? plru0_48 : _GEN_1068; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1390 = s2_reg_dirty ? plru0_49 : _GEN_1069; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1391 = s2_reg_dirty ? plru0_50 : _GEN_1070; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1392 = s2_reg_dirty ? plru0_51 : _GEN_1071; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1393 = s2_reg_dirty ? plru0_52 : _GEN_1072; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1394 = s2_reg_dirty ? plru0_53 : _GEN_1073; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1395 = s2_reg_dirty ? plru0_54 : _GEN_1074; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1396 = s2_reg_dirty ? plru0_55 : _GEN_1075; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1397 = s2_reg_dirty ? plru0_56 : _GEN_1076; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1398 = s2_reg_dirty ? plru0_57 : _GEN_1077; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1399 = s2_reg_dirty ? plru0_58 : _GEN_1078; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1400 = s2_reg_dirty ? plru0_59 : _GEN_1079; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1401 = s2_reg_dirty ? plru0_60 : _GEN_1080; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1402 = s2_reg_dirty ? plru0_61 : _GEN_1081; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1403 = s2_reg_dirty ? plru0_62 : _GEN_1082; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1404 = s2_reg_dirty ? plru0_63 : _GEN_1083; // @[Cache.scala 129:22 385:27]
  wire  _GEN_1405 = s2_reg_dirty ? plru1_0 : _GEN_1212; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1406 = s2_reg_dirty ? plru1_1 : _GEN_1213; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1407 = s2_reg_dirty ? plru1_2 : _GEN_1214; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1408 = s2_reg_dirty ? plru1_3 : _GEN_1215; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1409 = s2_reg_dirty ? plru1_4 : _GEN_1216; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1410 = s2_reg_dirty ? plru1_5 : _GEN_1217; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1411 = s2_reg_dirty ? plru1_6 : _GEN_1218; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1412 = s2_reg_dirty ? plru1_7 : _GEN_1219; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1413 = s2_reg_dirty ? plru1_8 : _GEN_1220; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1414 = s2_reg_dirty ? plru1_9 : _GEN_1221; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1415 = s2_reg_dirty ? plru1_10 : _GEN_1222; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1416 = s2_reg_dirty ? plru1_11 : _GEN_1223; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1417 = s2_reg_dirty ? plru1_12 : _GEN_1224; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1418 = s2_reg_dirty ? plru1_13 : _GEN_1225; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1419 = s2_reg_dirty ? plru1_14 : _GEN_1226; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1420 = s2_reg_dirty ? plru1_15 : _GEN_1227; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1421 = s2_reg_dirty ? plru1_16 : _GEN_1228; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1422 = s2_reg_dirty ? plru1_17 : _GEN_1229; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1423 = s2_reg_dirty ? plru1_18 : _GEN_1230; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1424 = s2_reg_dirty ? plru1_19 : _GEN_1231; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1425 = s2_reg_dirty ? plru1_20 : _GEN_1232; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1426 = s2_reg_dirty ? plru1_21 : _GEN_1233; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1427 = s2_reg_dirty ? plru1_22 : _GEN_1234; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1428 = s2_reg_dirty ? plru1_23 : _GEN_1235; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1429 = s2_reg_dirty ? plru1_24 : _GEN_1236; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1430 = s2_reg_dirty ? plru1_25 : _GEN_1237; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1431 = s2_reg_dirty ? plru1_26 : _GEN_1238; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1432 = s2_reg_dirty ? plru1_27 : _GEN_1239; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1433 = s2_reg_dirty ? plru1_28 : _GEN_1240; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1434 = s2_reg_dirty ? plru1_29 : _GEN_1241; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1435 = s2_reg_dirty ? plru1_30 : _GEN_1242; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1436 = s2_reg_dirty ? plru1_31 : _GEN_1243; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1437 = s2_reg_dirty ? plru1_32 : _GEN_1244; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1438 = s2_reg_dirty ? plru1_33 : _GEN_1245; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1439 = s2_reg_dirty ? plru1_34 : _GEN_1246; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1440 = s2_reg_dirty ? plru1_35 : _GEN_1247; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1441 = s2_reg_dirty ? plru1_36 : _GEN_1248; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1442 = s2_reg_dirty ? plru1_37 : _GEN_1249; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1443 = s2_reg_dirty ? plru1_38 : _GEN_1250; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1444 = s2_reg_dirty ? plru1_39 : _GEN_1251; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1445 = s2_reg_dirty ? plru1_40 : _GEN_1252; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1446 = s2_reg_dirty ? plru1_41 : _GEN_1253; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1447 = s2_reg_dirty ? plru1_42 : _GEN_1254; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1448 = s2_reg_dirty ? plru1_43 : _GEN_1255; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1449 = s2_reg_dirty ? plru1_44 : _GEN_1256; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1450 = s2_reg_dirty ? plru1_45 : _GEN_1257; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1451 = s2_reg_dirty ? plru1_46 : _GEN_1258; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1452 = s2_reg_dirty ? plru1_47 : _GEN_1259; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1453 = s2_reg_dirty ? plru1_48 : _GEN_1260; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1454 = s2_reg_dirty ? plru1_49 : _GEN_1261; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1455 = s2_reg_dirty ? plru1_50 : _GEN_1262; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1456 = s2_reg_dirty ? plru1_51 : _GEN_1263; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1457 = s2_reg_dirty ? plru1_52 : _GEN_1264; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1458 = s2_reg_dirty ? plru1_53 : _GEN_1265; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1459 = s2_reg_dirty ? plru1_54 : _GEN_1266; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1460 = s2_reg_dirty ? plru1_55 : _GEN_1267; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1461 = s2_reg_dirty ? plru1_56 : _GEN_1268; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1462 = s2_reg_dirty ? plru1_57 : _GEN_1269; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1463 = s2_reg_dirty ? plru1_58 : _GEN_1270; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1464 = s2_reg_dirty ? plru1_59 : _GEN_1271; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1465 = s2_reg_dirty ? plru1_60 : _GEN_1272; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1466 = s2_reg_dirty ? plru1_61 : _GEN_1273; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1467 = s2_reg_dirty ? plru1_62 : _GEN_1274; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1468 = s2_reg_dirty ? plru1_63 : _GEN_1275; // @[Cache.scala 131:22 385:27]
  wire  _GEN_1469 = s2_reg_dirty ? plru2_0 : _GEN_1276; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1470 = s2_reg_dirty ? plru2_1 : _GEN_1277; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1471 = s2_reg_dirty ? plru2_2 : _GEN_1278; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1472 = s2_reg_dirty ? plru2_3 : _GEN_1279; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1473 = s2_reg_dirty ? plru2_4 : _GEN_1280; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1474 = s2_reg_dirty ? plru2_5 : _GEN_1281; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1475 = s2_reg_dirty ? plru2_6 : _GEN_1282; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1476 = s2_reg_dirty ? plru2_7 : _GEN_1283; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1477 = s2_reg_dirty ? plru2_8 : _GEN_1284; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1478 = s2_reg_dirty ? plru2_9 : _GEN_1285; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1479 = s2_reg_dirty ? plru2_10 : _GEN_1286; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1480 = s2_reg_dirty ? plru2_11 : _GEN_1287; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1481 = s2_reg_dirty ? plru2_12 : _GEN_1288; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1482 = s2_reg_dirty ? plru2_13 : _GEN_1289; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1483 = s2_reg_dirty ? plru2_14 : _GEN_1290; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1484 = s2_reg_dirty ? plru2_15 : _GEN_1291; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1485 = s2_reg_dirty ? plru2_16 : _GEN_1292; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1486 = s2_reg_dirty ? plru2_17 : _GEN_1293; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1487 = s2_reg_dirty ? plru2_18 : _GEN_1294; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1488 = s2_reg_dirty ? plru2_19 : _GEN_1295; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1489 = s2_reg_dirty ? plru2_20 : _GEN_1296; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1490 = s2_reg_dirty ? plru2_21 : _GEN_1297; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1491 = s2_reg_dirty ? plru2_22 : _GEN_1298; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1492 = s2_reg_dirty ? plru2_23 : _GEN_1299; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1493 = s2_reg_dirty ? plru2_24 : _GEN_1300; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1494 = s2_reg_dirty ? plru2_25 : _GEN_1301; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1495 = s2_reg_dirty ? plru2_26 : _GEN_1302; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1496 = s2_reg_dirty ? plru2_27 : _GEN_1303; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1497 = s2_reg_dirty ? plru2_28 : _GEN_1304; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1498 = s2_reg_dirty ? plru2_29 : _GEN_1305; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1499 = s2_reg_dirty ? plru2_30 : _GEN_1306; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1500 = s2_reg_dirty ? plru2_31 : _GEN_1307; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1501 = s2_reg_dirty ? plru2_32 : _GEN_1308; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1502 = s2_reg_dirty ? plru2_33 : _GEN_1309; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1503 = s2_reg_dirty ? plru2_34 : _GEN_1310; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1504 = s2_reg_dirty ? plru2_35 : _GEN_1311; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1505 = s2_reg_dirty ? plru2_36 : _GEN_1312; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1506 = s2_reg_dirty ? plru2_37 : _GEN_1313; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1507 = s2_reg_dirty ? plru2_38 : _GEN_1314; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1508 = s2_reg_dirty ? plru2_39 : _GEN_1315; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1509 = s2_reg_dirty ? plru2_40 : _GEN_1316; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1510 = s2_reg_dirty ? plru2_41 : _GEN_1317; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1511 = s2_reg_dirty ? plru2_42 : _GEN_1318; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1512 = s2_reg_dirty ? plru2_43 : _GEN_1319; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1513 = s2_reg_dirty ? plru2_44 : _GEN_1320; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1514 = s2_reg_dirty ? plru2_45 : _GEN_1321; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1515 = s2_reg_dirty ? plru2_46 : _GEN_1322; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1516 = s2_reg_dirty ? plru2_47 : _GEN_1323; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1517 = s2_reg_dirty ? plru2_48 : _GEN_1324; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1518 = s2_reg_dirty ? plru2_49 : _GEN_1325; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1519 = s2_reg_dirty ? plru2_50 : _GEN_1326; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1520 = s2_reg_dirty ? plru2_51 : _GEN_1327; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1521 = s2_reg_dirty ? plru2_52 : _GEN_1328; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1522 = s2_reg_dirty ? plru2_53 : _GEN_1329; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1523 = s2_reg_dirty ? plru2_54 : _GEN_1330; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1524 = s2_reg_dirty ? plru2_55 : _GEN_1331; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1525 = s2_reg_dirty ? plru2_56 : _GEN_1332; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1526 = s2_reg_dirty ? plru2_57 : _GEN_1333; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1527 = s2_reg_dirty ? plru2_58 : _GEN_1334; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1528 = s2_reg_dirty ? plru2_59 : _GEN_1335; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1529 = s2_reg_dirty ? plru2_60 : _GEN_1336; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1530 = s2_reg_dirty ? plru2_61 : _GEN_1337; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1531 = s2_reg_dirty ? plru2_62 : _GEN_1338; // @[Cache.scala 133:22 385:27]
  wire  _GEN_1532 = s2_reg_dirty ? plru2_63 : _GEN_1339; // @[Cache.scala 133:22 385:27]
  wire [3:0] _GEN_1533 = _T_320 ? 4'h5 : state; // @[Cache.scala 393:29 394:15 213:22]
  wire [3:0] _GEN_1534 = _T_320 ? 4'h6 : state; // @[Cache.scala 398:29 399:15 213:22]
  wire  _GEN_1855 = _T_322 ? _GEN_1020 : plru0_0; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1856 = _T_322 ? _GEN_1021 : plru0_1; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1857 = _T_322 ? _GEN_1022 : plru0_2; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1858 = _T_322 ? _GEN_1023 : plru0_3; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1859 = _T_322 ? _GEN_1024 : plru0_4; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1860 = _T_322 ? _GEN_1025 : plru0_5; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1861 = _T_322 ? _GEN_1026 : plru0_6; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1862 = _T_322 ? _GEN_1027 : plru0_7; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1863 = _T_322 ? _GEN_1028 : plru0_8; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1864 = _T_322 ? _GEN_1029 : plru0_9; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1865 = _T_322 ? _GEN_1030 : plru0_10; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1866 = _T_322 ? _GEN_1031 : plru0_11; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1867 = _T_322 ? _GEN_1032 : plru0_12; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1868 = _T_322 ? _GEN_1033 : plru0_13; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1869 = _T_322 ? _GEN_1034 : plru0_14; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1870 = _T_322 ? _GEN_1035 : plru0_15; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1871 = _T_322 ? _GEN_1036 : plru0_16; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1872 = _T_322 ? _GEN_1037 : plru0_17; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1873 = _T_322 ? _GEN_1038 : plru0_18; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1874 = _T_322 ? _GEN_1039 : plru0_19; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1875 = _T_322 ? _GEN_1040 : plru0_20; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1876 = _T_322 ? _GEN_1041 : plru0_21; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1877 = _T_322 ? _GEN_1042 : plru0_22; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1878 = _T_322 ? _GEN_1043 : plru0_23; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1879 = _T_322 ? _GEN_1044 : plru0_24; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1880 = _T_322 ? _GEN_1045 : plru0_25; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1881 = _T_322 ? _GEN_1046 : plru0_26; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1882 = _T_322 ? _GEN_1047 : plru0_27; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1883 = _T_322 ? _GEN_1048 : plru0_28; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1884 = _T_322 ? _GEN_1049 : plru0_29; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1885 = _T_322 ? _GEN_1050 : plru0_30; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1886 = _T_322 ? _GEN_1051 : plru0_31; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1887 = _T_322 ? _GEN_1052 : plru0_32; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1888 = _T_322 ? _GEN_1053 : plru0_33; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1889 = _T_322 ? _GEN_1054 : plru0_34; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1890 = _T_322 ? _GEN_1055 : plru0_35; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1891 = _T_322 ? _GEN_1056 : plru0_36; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1892 = _T_322 ? _GEN_1057 : plru0_37; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1893 = _T_322 ? _GEN_1058 : plru0_38; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1894 = _T_322 ? _GEN_1059 : plru0_39; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1895 = _T_322 ? _GEN_1060 : plru0_40; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1896 = _T_322 ? _GEN_1061 : plru0_41; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1897 = _T_322 ? _GEN_1062 : plru0_42; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1898 = _T_322 ? _GEN_1063 : plru0_43; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1899 = _T_322 ? _GEN_1064 : plru0_44; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1900 = _T_322 ? _GEN_1065 : plru0_45; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1901 = _T_322 ? _GEN_1066 : plru0_46; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1902 = _T_322 ? _GEN_1067 : plru0_47; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1903 = _T_322 ? _GEN_1068 : plru0_48; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1904 = _T_322 ? _GEN_1069 : plru0_49; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1905 = _T_322 ? _GEN_1070 : plru0_50; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1906 = _T_322 ? _GEN_1071 : plru0_51; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1907 = _T_322 ? _GEN_1072 : plru0_52; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1908 = _T_322 ? _GEN_1073 : plru0_53; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1909 = _T_322 ? _GEN_1074 : plru0_54; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1910 = _T_322 ? _GEN_1075 : plru0_55; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1911 = _T_322 ? _GEN_1076 : plru0_56; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1912 = _T_322 ? _GEN_1077 : plru0_57; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1913 = _T_322 ? _GEN_1078 : plru0_58; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1914 = _T_322 ? _GEN_1079 : plru0_59; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1915 = _T_322 ? _GEN_1080 : plru0_60; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1916 = _T_322 ? _GEN_1081 : plru0_61; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1917 = _T_322 ? _GEN_1082 : plru0_62; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1918 = _T_322 ? _GEN_1083 : plru0_63; // @[Cache.scala 129:22 404:30]
  wire  _GEN_1919 = _T_322 ? _GEN_1212 : plru1_0; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1920 = _T_322 ? _GEN_1213 : plru1_1; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1921 = _T_322 ? _GEN_1214 : plru1_2; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1922 = _T_322 ? _GEN_1215 : plru1_3; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1923 = _T_322 ? _GEN_1216 : plru1_4; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1924 = _T_322 ? _GEN_1217 : plru1_5; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1925 = _T_322 ? _GEN_1218 : plru1_6; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1926 = _T_322 ? _GEN_1219 : plru1_7; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1927 = _T_322 ? _GEN_1220 : plru1_8; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1928 = _T_322 ? _GEN_1221 : plru1_9; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1929 = _T_322 ? _GEN_1222 : plru1_10; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1930 = _T_322 ? _GEN_1223 : plru1_11; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1931 = _T_322 ? _GEN_1224 : plru1_12; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1932 = _T_322 ? _GEN_1225 : plru1_13; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1933 = _T_322 ? _GEN_1226 : plru1_14; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1934 = _T_322 ? _GEN_1227 : plru1_15; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1935 = _T_322 ? _GEN_1228 : plru1_16; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1936 = _T_322 ? _GEN_1229 : plru1_17; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1937 = _T_322 ? _GEN_1230 : plru1_18; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1938 = _T_322 ? _GEN_1231 : plru1_19; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1939 = _T_322 ? _GEN_1232 : plru1_20; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1940 = _T_322 ? _GEN_1233 : plru1_21; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1941 = _T_322 ? _GEN_1234 : plru1_22; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1942 = _T_322 ? _GEN_1235 : plru1_23; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1943 = _T_322 ? _GEN_1236 : plru1_24; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1944 = _T_322 ? _GEN_1237 : plru1_25; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1945 = _T_322 ? _GEN_1238 : plru1_26; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1946 = _T_322 ? _GEN_1239 : plru1_27; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1947 = _T_322 ? _GEN_1240 : plru1_28; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1948 = _T_322 ? _GEN_1241 : plru1_29; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1949 = _T_322 ? _GEN_1242 : plru1_30; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1950 = _T_322 ? _GEN_1243 : plru1_31; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1951 = _T_322 ? _GEN_1244 : plru1_32; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1952 = _T_322 ? _GEN_1245 : plru1_33; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1953 = _T_322 ? _GEN_1246 : plru1_34; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1954 = _T_322 ? _GEN_1247 : plru1_35; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1955 = _T_322 ? _GEN_1248 : plru1_36; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1956 = _T_322 ? _GEN_1249 : plru1_37; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1957 = _T_322 ? _GEN_1250 : plru1_38; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1958 = _T_322 ? _GEN_1251 : plru1_39; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1959 = _T_322 ? _GEN_1252 : plru1_40; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1960 = _T_322 ? _GEN_1253 : plru1_41; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1961 = _T_322 ? _GEN_1254 : plru1_42; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1962 = _T_322 ? _GEN_1255 : plru1_43; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1963 = _T_322 ? _GEN_1256 : plru1_44; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1964 = _T_322 ? _GEN_1257 : plru1_45; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1965 = _T_322 ? _GEN_1258 : plru1_46; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1966 = _T_322 ? _GEN_1259 : plru1_47; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1967 = _T_322 ? _GEN_1260 : plru1_48; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1968 = _T_322 ? _GEN_1261 : plru1_49; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1969 = _T_322 ? _GEN_1262 : plru1_50; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1970 = _T_322 ? _GEN_1263 : plru1_51; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1971 = _T_322 ? _GEN_1264 : plru1_52; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1972 = _T_322 ? _GEN_1265 : plru1_53; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1973 = _T_322 ? _GEN_1266 : plru1_54; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1974 = _T_322 ? _GEN_1267 : plru1_55; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1975 = _T_322 ? _GEN_1268 : plru1_56; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1976 = _T_322 ? _GEN_1269 : plru1_57; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1977 = _T_322 ? _GEN_1270 : plru1_58; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1978 = _T_322 ? _GEN_1271 : plru1_59; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1979 = _T_322 ? _GEN_1272 : plru1_60; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1980 = _T_322 ? _GEN_1273 : plru1_61; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1981 = _T_322 ? _GEN_1274 : plru1_62; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1982 = _T_322 ? _GEN_1275 : plru1_63; // @[Cache.scala 131:22 404:30]
  wire  _GEN_1983 = _T_322 ? _GEN_1276 : plru2_0; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1984 = _T_322 ? _GEN_1277 : plru2_1; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1985 = _T_322 ? _GEN_1278 : plru2_2; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1986 = _T_322 ? _GEN_1279 : plru2_3; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1987 = _T_322 ? _GEN_1280 : plru2_4; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1988 = _T_322 ? _GEN_1281 : plru2_5; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1989 = _T_322 ? _GEN_1282 : plru2_6; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1990 = _T_322 ? _GEN_1283 : plru2_7; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1991 = _T_322 ? _GEN_1284 : plru2_8; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1992 = _T_322 ? _GEN_1285 : plru2_9; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1993 = _T_322 ? _GEN_1286 : plru2_10; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1994 = _T_322 ? _GEN_1287 : plru2_11; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1995 = _T_322 ? _GEN_1288 : plru2_12; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1996 = _T_322 ? _GEN_1289 : plru2_13; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1997 = _T_322 ? _GEN_1290 : plru2_14; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1998 = _T_322 ? _GEN_1291 : plru2_15; // @[Cache.scala 133:22 404:30]
  wire  _GEN_1999 = _T_322 ? _GEN_1292 : plru2_16; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2000 = _T_322 ? _GEN_1293 : plru2_17; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2001 = _T_322 ? _GEN_1294 : plru2_18; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2002 = _T_322 ? _GEN_1295 : plru2_19; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2003 = _T_322 ? _GEN_1296 : plru2_20; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2004 = _T_322 ? _GEN_1297 : plru2_21; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2005 = _T_322 ? _GEN_1298 : plru2_22; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2006 = _T_322 ? _GEN_1299 : plru2_23; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2007 = _T_322 ? _GEN_1300 : plru2_24; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2008 = _T_322 ? _GEN_1301 : plru2_25; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2009 = _T_322 ? _GEN_1302 : plru2_26; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2010 = _T_322 ? _GEN_1303 : plru2_27; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2011 = _T_322 ? _GEN_1304 : plru2_28; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2012 = _T_322 ? _GEN_1305 : plru2_29; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2013 = _T_322 ? _GEN_1306 : plru2_30; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2014 = _T_322 ? _GEN_1307 : plru2_31; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2015 = _T_322 ? _GEN_1308 : plru2_32; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2016 = _T_322 ? _GEN_1309 : plru2_33; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2017 = _T_322 ? _GEN_1310 : plru2_34; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2018 = _T_322 ? _GEN_1311 : plru2_35; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2019 = _T_322 ? _GEN_1312 : plru2_36; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2020 = _T_322 ? _GEN_1313 : plru2_37; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2021 = _T_322 ? _GEN_1314 : plru2_38; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2022 = _T_322 ? _GEN_1315 : plru2_39; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2023 = _T_322 ? _GEN_1316 : plru2_40; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2024 = _T_322 ? _GEN_1317 : plru2_41; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2025 = _T_322 ? _GEN_1318 : plru2_42; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2026 = _T_322 ? _GEN_1319 : plru2_43; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2027 = _T_322 ? _GEN_1320 : plru2_44; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2028 = _T_322 ? _GEN_1321 : plru2_45; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2029 = _T_322 ? _GEN_1322 : plru2_46; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2030 = _T_322 ? _GEN_1323 : plru2_47; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2031 = _T_322 ? _GEN_1324 : plru2_48; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2032 = _T_322 ? _GEN_1325 : plru2_49; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2033 = _T_322 ? _GEN_1326 : plru2_50; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2034 = _T_322 ? _GEN_1327 : plru2_51; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2035 = _T_322 ? _GEN_1328 : plru2_52; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2036 = _T_322 ? _GEN_1329 : plru2_53; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2037 = _T_322 ? _GEN_1330 : plru2_54; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2038 = _T_322 ? _GEN_1331 : plru2_55; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2039 = _T_322 ? _GEN_1332 : plru2_56; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2040 = _T_322 ? _GEN_1333 : plru2_57; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2041 = _T_322 ? _GEN_1334 : plru2_58; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2042 = _T_322 ? _GEN_1335 : plru2_59; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2043 = _T_322 ? _GEN_1336 : plru2_60; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2044 = _T_322 ? _GEN_1337 : plru2_61; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2045 = _T_322 ? _GEN_1338 : plru2_62; // @[Cache.scala 133:22 404:30]
  wire  _GEN_2046 = _T_322 ? _GEN_1339 : plru2_63; // @[Cache.scala 133:22 404:30]
  wire [3:0] _GEN_2047 = _T_322 ? 4'h7 : state; // @[Cache.scala 404:30 406:15 213:22]
  reg [63:0] REG_12; // @[Cache.scala 410:36]
  wire  _T_606 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_2048 = _T_606 ? 4'h8 : state; // @[Cache.scala 411:29 412:15 213:22]
  wire [63:0] _GEN_2049 = 4'h7 == state ? REG_12 : 64'h0; // @[Cache.scala 318:18 289:22 410:26]
  wire [3:0] _GEN_2050 = 4'h7 == state ? _GEN_2048 : state; // @[Cache.scala 318:18 213:22]
  wire  _GEN_2051 = 4'h6 == state ? 1'h0 : _GEN_27; // @[Cache.scala 318:18 403:14]
  wire  _GEN_2052 = 4'h6 == state ? _GEN_1855 : plru0_0; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2053 = 4'h6 == state ? _GEN_1856 : plru0_1; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2054 = 4'h6 == state ? _GEN_1857 : plru0_2; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2055 = 4'h6 == state ? _GEN_1858 : plru0_3; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2056 = 4'h6 == state ? _GEN_1859 : plru0_4; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2057 = 4'h6 == state ? _GEN_1860 : plru0_5; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2058 = 4'h6 == state ? _GEN_1861 : plru0_6; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2059 = 4'h6 == state ? _GEN_1862 : plru0_7; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2060 = 4'h6 == state ? _GEN_1863 : plru0_8; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2061 = 4'h6 == state ? _GEN_1864 : plru0_9; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2062 = 4'h6 == state ? _GEN_1865 : plru0_10; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2063 = 4'h6 == state ? _GEN_1866 : plru0_11; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2064 = 4'h6 == state ? _GEN_1867 : plru0_12; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2065 = 4'h6 == state ? _GEN_1868 : plru0_13; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2066 = 4'h6 == state ? _GEN_1869 : plru0_14; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2067 = 4'h6 == state ? _GEN_1870 : plru0_15; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2068 = 4'h6 == state ? _GEN_1871 : plru0_16; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2069 = 4'h6 == state ? _GEN_1872 : plru0_17; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2070 = 4'h6 == state ? _GEN_1873 : plru0_18; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2071 = 4'h6 == state ? _GEN_1874 : plru0_19; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2072 = 4'h6 == state ? _GEN_1875 : plru0_20; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2073 = 4'h6 == state ? _GEN_1876 : plru0_21; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2074 = 4'h6 == state ? _GEN_1877 : plru0_22; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2075 = 4'h6 == state ? _GEN_1878 : plru0_23; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2076 = 4'h6 == state ? _GEN_1879 : plru0_24; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2077 = 4'h6 == state ? _GEN_1880 : plru0_25; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2078 = 4'h6 == state ? _GEN_1881 : plru0_26; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2079 = 4'h6 == state ? _GEN_1882 : plru0_27; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2080 = 4'h6 == state ? _GEN_1883 : plru0_28; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2081 = 4'h6 == state ? _GEN_1884 : plru0_29; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2082 = 4'h6 == state ? _GEN_1885 : plru0_30; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2083 = 4'h6 == state ? _GEN_1886 : plru0_31; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2084 = 4'h6 == state ? _GEN_1887 : plru0_32; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2085 = 4'h6 == state ? _GEN_1888 : plru0_33; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2086 = 4'h6 == state ? _GEN_1889 : plru0_34; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2087 = 4'h6 == state ? _GEN_1890 : plru0_35; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2088 = 4'h6 == state ? _GEN_1891 : plru0_36; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2089 = 4'h6 == state ? _GEN_1892 : plru0_37; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2090 = 4'h6 == state ? _GEN_1893 : plru0_38; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2091 = 4'h6 == state ? _GEN_1894 : plru0_39; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2092 = 4'h6 == state ? _GEN_1895 : plru0_40; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2093 = 4'h6 == state ? _GEN_1896 : plru0_41; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2094 = 4'h6 == state ? _GEN_1897 : plru0_42; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2095 = 4'h6 == state ? _GEN_1898 : plru0_43; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2096 = 4'h6 == state ? _GEN_1899 : plru0_44; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2097 = 4'h6 == state ? _GEN_1900 : plru0_45; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2098 = 4'h6 == state ? _GEN_1901 : plru0_46; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2099 = 4'h6 == state ? _GEN_1902 : plru0_47; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2100 = 4'h6 == state ? _GEN_1903 : plru0_48; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2101 = 4'h6 == state ? _GEN_1904 : plru0_49; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2102 = 4'h6 == state ? _GEN_1905 : plru0_50; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2103 = 4'h6 == state ? _GEN_1906 : plru0_51; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2104 = 4'h6 == state ? _GEN_1907 : plru0_52; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2105 = 4'h6 == state ? _GEN_1908 : plru0_53; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2106 = 4'h6 == state ? _GEN_1909 : plru0_54; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2107 = 4'h6 == state ? _GEN_1910 : plru0_55; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2108 = 4'h6 == state ? _GEN_1911 : plru0_56; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2109 = 4'h6 == state ? _GEN_1912 : plru0_57; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2110 = 4'h6 == state ? _GEN_1913 : plru0_58; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2111 = 4'h6 == state ? _GEN_1914 : plru0_59; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2112 = 4'h6 == state ? _GEN_1915 : plru0_60; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2113 = 4'h6 == state ? _GEN_1916 : plru0_61; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2114 = 4'h6 == state ? _GEN_1917 : plru0_62; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2115 = 4'h6 == state ? _GEN_1918 : plru0_63; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2116 = 4'h6 == state ? _GEN_1919 : plru1_0; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2117 = 4'h6 == state ? _GEN_1920 : plru1_1; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2118 = 4'h6 == state ? _GEN_1921 : plru1_2; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2119 = 4'h6 == state ? _GEN_1922 : plru1_3; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2120 = 4'h6 == state ? _GEN_1923 : plru1_4; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2121 = 4'h6 == state ? _GEN_1924 : plru1_5; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2122 = 4'h6 == state ? _GEN_1925 : plru1_6; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2123 = 4'h6 == state ? _GEN_1926 : plru1_7; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2124 = 4'h6 == state ? _GEN_1927 : plru1_8; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2125 = 4'h6 == state ? _GEN_1928 : plru1_9; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2126 = 4'h6 == state ? _GEN_1929 : plru1_10; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2127 = 4'h6 == state ? _GEN_1930 : plru1_11; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2128 = 4'h6 == state ? _GEN_1931 : plru1_12; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2129 = 4'h6 == state ? _GEN_1932 : plru1_13; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2130 = 4'h6 == state ? _GEN_1933 : plru1_14; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2131 = 4'h6 == state ? _GEN_1934 : plru1_15; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2132 = 4'h6 == state ? _GEN_1935 : plru1_16; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2133 = 4'h6 == state ? _GEN_1936 : plru1_17; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2134 = 4'h6 == state ? _GEN_1937 : plru1_18; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2135 = 4'h6 == state ? _GEN_1938 : plru1_19; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2136 = 4'h6 == state ? _GEN_1939 : plru1_20; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2137 = 4'h6 == state ? _GEN_1940 : plru1_21; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2138 = 4'h6 == state ? _GEN_1941 : plru1_22; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2139 = 4'h6 == state ? _GEN_1942 : plru1_23; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2140 = 4'h6 == state ? _GEN_1943 : plru1_24; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2141 = 4'h6 == state ? _GEN_1944 : plru1_25; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2142 = 4'h6 == state ? _GEN_1945 : plru1_26; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2143 = 4'h6 == state ? _GEN_1946 : plru1_27; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2144 = 4'h6 == state ? _GEN_1947 : plru1_28; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2145 = 4'h6 == state ? _GEN_1948 : plru1_29; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2146 = 4'h6 == state ? _GEN_1949 : plru1_30; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2147 = 4'h6 == state ? _GEN_1950 : plru1_31; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2148 = 4'h6 == state ? _GEN_1951 : plru1_32; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2149 = 4'h6 == state ? _GEN_1952 : plru1_33; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2150 = 4'h6 == state ? _GEN_1953 : plru1_34; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2151 = 4'h6 == state ? _GEN_1954 : plru1_35; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2152 = 4'h6 == state ? _GEN_1955 : plru1_36; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2153 = 4'h6 == state ? _GEN_1956 : plru1_37; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2154 = 4'h6 == state ? _GEN_1957 : plru1_38; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2155 = 4'h6 == state ? _GEN_1958 : plru1_39; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2156 = 4'h6 == state ? _GEN_1959 : plru1_40; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2157 = 4'h6 == state ? _GEN_1960 : plru1_41; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2158 = 4'h6 == state ? _GEN_1961 : plru1_42; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2159 = 4'h6 == state ? _GEN_1962 : plru1_43; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2160 = 4'h6 == state ? _GEN_1963 : plru1_44; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2161 = 4'h6 == state ? _GEN_1964 : plru1_45; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2162 = 4'h6 == state ? _GEN_1965 : plru1_46; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2163 = 4'h6 == state ? _GEN_1966 : plru1_47; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2164 = 4'h6 == state ? _GEN_1967 : plru1_48; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2165 = 4'h6 == state ? _GEN_1968 : plru1_49; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2166 = 4'h6 == state ? _GEN_1969 : plru1_50; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2167 = 4'h6 == state ? _GEN_1970 : plru1_51; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2168 = 4'h6 == state ? _GEN_1971 : plru1_52; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2169 = 4'h6 == state ? _GEN_1972 : plru1_53; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2170 = 4'h6 == state ? _GEN_1973 : plru1_54; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2171 = 4'h6 == state ? _GEN_1974 : plru1_55; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2172 = 4'h6 == state ? _GEN_1975 : plru1_56; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2173 = 4'h6 == state ? _GEN_1976 : plru1_57; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2174 = 4'h6 == state ? _GEN_1977 : plru1_58; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2175 = 4'h6 == state ? _GEN_1978 : plru1_59; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2176 = 4'h6 == state ? _GEN_1979 : plru1_60; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2177 = 4'h6 == state ? _GEN_1980 : plru1_61; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2178 = 4'h6 == state ? _GEN_1981 : plru1_62; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2179 = 4'h6 == state ? _GEN_1982 : plru1_63; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2180 = 4'h6 == state ? _GEN_1983 : plru2_0; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2181 = 4'h6 == state ? _GEN_1984 : plru2_1; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2182 = 4'h6 == state ? _GEN_1985 : plru2_2; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2183 = 4'h6 == state ? _GEN_1986 : plru2_3; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2184 = 4'h6 == state ? _GEN_1987 : plru2_4; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2185 = 4'h6 == state ? _GEN_1988 : plru2_5; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2186 = 4'h6 == state ? _GEN_1989 : plru2_6; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2187 = 4'h6 == state ? _GEN_1990 : plru2_7; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2188 = 4'h6 == state ? _GEN_1991 : plru2_8; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2189 = 4'h6 == state ? _GEN_1992 : plru2_9; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2190 = 4'h6 == state ? _GEN_1993 : plru2_10; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2191 = 4'h6 == state ? _GEN_1994 : plru2_11; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2192 = 4'h6 == state ? _GEN_1995 : plru2_12; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2193 = 4'h6 == state ? _GEN_1996 : plru2_13; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2194 = 4'h6 == state ? _GEN_1997 : plru2_14; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2195 = 4'h6 == state ? _GEN_1998 : plru2_15; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2196 = 4'h6 == state ? _GEN_1999 : plru2_16; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2197 = 4'h6 == state ? _GEN_2000 : plru2_17; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2198 = 4'h6 == state ? _GEN_2001 : plru2_18; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2199 = 4'h6 == state ? _GEN_2002 : plru2_19; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2200 = 4'h6 == state ? _GEN_2003 : plru2_20; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2201 = 4'h6 == state ? _GEN_2004 : plru2_21; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2202 = 4'h6 == state ? _GEN_2005 : plru2_22; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2203 = 4'h6 == state ? _GEN_2006 : plru2_23; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2204 = 4'h6 == state ? _GEN_2007 : plru2_24; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2205 = 4'h6 == state ? _GEN_2008 : plru2_25; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2206 = 4'h6 == state ? _GEN_2009 : plru2_26; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2207 = 4'h6 == state ? _GEN_2010 : plru2_27; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2208 = 4'h6 == state ? _GEN_2011 : plru2_28; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2209 = 4'h6 == state ? _GEN_2012 : plru2_29; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2210 = 4'h6 == state ? _GEN_2013 : plru2_30; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2211 = 4'h6 == state ? _GEN_2014 : plru2_31; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2212 = 4'h6 == state ? _GEN_2015 : plru2_32; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2213 = 4'h6 == state ? _GEN_2016 : plru2_33; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2214 = 4'h6 == state ? _GEN_2017 : plru2_34; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2215 = 4'h6 == state ? _GEN_2018 : plru2_35; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2216 = 4'h6 == state ? _GEN_2019 : plru2_36; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2217 = 4'h6 == state ? _GEN_2020 : plru2_37; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2218 = 4'h6 == state ? _GEN_2021 : plru2_38; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2219 = 4'h6 == state ? _GEN_2022 : plru2_39; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2220 = 4'h6 == state ? _GEN_2023 : plru2_40; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2221 = 4'h6 == state ? _GEN_2024 : plru2_41; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2222 = 4'h6 == state ? _GEN_2025 : plru2_42; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2223 = 4'h6 == state ? _GEN_2026 : plru2_43; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2224 = 4'h6 == state ? _GEN_2027 : plru2_44; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2225 = 4'h6 == state ? _GEN_2028 : plru2_45; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2226 = 4'h6 == state ? _GEN_2029 : plru2_46; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2227 = 4'h6 == state ? _GEN_2030 : plru2_47; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2228 = 4'h6 == state ? _GEN_2031 : plru2_48; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2229 = 4'h6 == state ? _GEN_2032 : plru2_49; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2230 = 4'h6 == state ? _GEN_2033 : plru2_50; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2231 = 4'h6 == state ? _GEN_2034 : plru2_51; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2232 = 4'h6 == state ? _GEN_2035 : plru2_52; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2233 = 4'h6 == state ? _GEN_2036 : plru2_53; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2234 = 4'h6 == state ? _GEN_2037 : plru2_54; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2235 = 4'h6 == state ? _GEN_2038 : plru2_55; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2236 = 4'h6 == state ? _GEN_2039 : plru2_56; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2237 = 4'h6 == state ? _GEN_2040 : plru2_57; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2238 = 4'h6 == state ? _GEN_2041 : plru2_58; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2239 = 4'h6 == state ? _GEN_2042 : plru2_59; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2240 = 4'h6 == state ? _GEN_2043 : plru2_60; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2241 = 4'h6 == state ? _GEN_2044 : plru2_61; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2242 = 4'h6 == state ? _GEN_2045 : plru2_62; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2243 = 4'h6 == state ? _GEN_2046 : plru2_63; // @[Cache.scala 318:18 133:22]
  wire [3:0] _GEN_2244 = 4'h6 == state ? _GEN_2047 : _GEN_2050; // @[Cache.scala 318:18]
  wire [63:0] _GEN_2245 = 4'h6 == state ? 64'h0 : _GEN_2049; // @[Cache.scala 318:18 289:22]
  wire [3:0] _GEN_2246 = 4'h5 == state ? _GEN_1534 : _GEN_2244; // @[Cache.scala 318:18]
  wire  _GEN_2247 = 4'h5 == state ? _GEN_27 : _GEN_2051; // @[Cache.scala 318:18]
  wire  _GEN_2248 = 4'h5 == state ? plru0_0 : _GEN_2052; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2249 = 4'h5 == state ? plru0_1 : _GEN_2053; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2250 = 4'h5 == state ? plru0_2 : _GEN_2054; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2251 = 4'h5 == state ? plru0_3 : _GEN_2055; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2252 = 4'h5 == state ? plru0_4 : _GEN_2056; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2253 = 4'h5 == state ? plru0_5 : _GEN_2057; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2254 = 4'h5 == state ? plru0_6 : _GEN_2058; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2255 = 4'h5 == state ? plru0_7 : _GEN_2059; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2256 = 4'h5 == state ? plru0_8 : _GEN_2060; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2257 = 4'h5 == state ? plru0_9 : _GEN_2061; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2258 = 4'h5 == state ? plru0_10 : _GEN_2062; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2259 = 4'h5 == state ? plru0_11 : _GEN_2063; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2260 = 4'h5 == state ? plru0_12 : _GEN_2064; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2261 = 4'h5 == state ? plru0_13 : _GEN_2065; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2262 = 4'h5 == state ? plru0_14 : _GEN_2066; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2263 = 4'h5 == state ? plru0_15 : _GEN_2067; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2264 = 4'h5 == state ? plru0_16 : _GEN_2068; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2265 = 4'h5 == state ? plru0_17 : _GEN_2069; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2266 = 4'h5 == state ? plru0_18 : _GEN_2070; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2267 = 4'h5 == state ? plru0_19 : _GEN_2071; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2268 = 4'h5 == state ? plru0_20 : _GEN_2072; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2269 = 4'h5 == state ? plru0_21 : _GEN_2073; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2270 = 4'h5 == state ? plru0_22 : _GEN_2074; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2271 = 4'h5 == state ? plru0_23 : _GEN_2075; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2272 = 4'h5 == state ? plru0_24 : _GEN_2076; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2273 = 4'h5 == state ? plru0_25 : _GEN_2077; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2274 = 4'h5 == state ? plru0_26 : _GEN_2078; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2275 = 4'h5 == state ? plru0_27 : _GEN_2079; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2276 = 4'h5 == state ? plru0_28 : _GEN_2080; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2277 = 4'h5 == state ? plru0_29 : _GEN_2081; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2278 = 4'h5 == state ? plru0_30 : _GEN_2082; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2279 = 4'h5 == state ? plru0_31 : _GEN_2083; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2280 = 4'h5 == state ? plru0_32 : _GEN_2084; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2281 = 4'h5 == state ? plru0_33 : _GEN_2085; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2282 = 4'h5 == state ? plru0_34 : _GEN_2086; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2283 = 4'h5 == state ? plru0_35 : _GEN_2087; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2284 = 4'h5 == state ? plru0_36 : _GEN_2088; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2285 = 4'h5 == state ? plru0_37 : _GEN_2089; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2286 = 4'h5 == state ? plru0_38 : _GEN_2090; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2287 = 4'h5 == state ? plru0_39 : _GEN_2091; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2288 = 4'h5 == state ? plru0_40 : _GEN_2092; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2289 = 4'h5 == state ? plru0_41 : _GEN_2093; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2290 = 4'h5 == state ? plru0_42 : _GEN_2094; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2291 = 4'h5 == state ? plru0_43 : _GEN_2095; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2292 = 4'h5 == state ? plru0_44 : _GEN_2096; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2293 = 4'h5 == state ? plru0_45 : _GEN_2097; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2294 = 4'h5 == state ? plru0_46 : _GEN_2098; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2295 = 4'h5 == state ? plru0_47 : _GEN_2099; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2296 = 4'h5 == state ? plru0_48 : _GEN_2100; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2297 = 4'h5 == state ? plru0_49 : _GEN_2101; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2298 = 4'h5 == state ? plru0_50 : _GEN_2102; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2299 = 4'h5 == state ? plru0_51 : _GEN_2103; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2300 = 4'h5 == state ? plru0_52 : _GEN_2104; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2301 = 4'h5 == state ? plru0_53 : _GEN_2105; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2302 = 4'h5 == state ? plru0_54 : _GEN_2106; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2303 = 4'h5 == state ? plru0_55 : _GEN_2107; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2304 = 4'h5 == state ? plru0_56 : _GEN_2108; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2305 = 4'h5 == state ? plru0_57 : _GEN_2109; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2306 = 4'h5 == state ? plru0_58 : _GEN_2110; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2307 = 4'h5 == state ? plru0_59 : _GEN_2111; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2308 = 4'h5 == state ? plru0_60 : _GEN_2112; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2309 = 4'h5 == state ? plru0_61 : _GEN_2113; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2310 = 4'h5 == state ? plru0_62 : _GEN_2114; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2311 = 4'h5 == state ? plru0_63 : _GEN_2115; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2312 = 4'h5 == state ? plru1_0 : _GEN_2116; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2313 = 4'h5 == state ? plru1_1 : _GEN_2117; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2314 = 4'h5 == state ? plru1_2 : _GEN_2118; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2315 = 4'h5 == state ? plru1_3 : _GEN_2119; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2316 = 4'h5 == state ? plru1_4 : _GEN_2120; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2317 = 4'h5 == state ? plru1_5 : _GEN_2121; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2318 = 4'h5 == state ? plru1_6 : _GEN_2122; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2319 = 4'h5 == state ? plru1_7 : _GEN_2123; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2320 = 4'h5 == state ? plru1_8 : _GEN_2124; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2321 = 4'h5 == state ? plru1_9 : _GEN_2125; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2322 = 4'h5 == state ? plru1_10 : _GEN_2126; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2323 = 4'h5 == state ? plru1_11 : _GEN_2127; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2324 = 4'h5 == state ? plru1_12 : _GEN_2128; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2325 = 4'h5 == state ? plru1_13 : _GEN_2129; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2326 = 4'h5 == state ? plru1_14 : _GEN_2130; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2327 = 4'h5 == state ? plru1_15 : _GEN_2131; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2328 = 4'h5 == state ? plru1_16 : _GEN_2132; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2329 = 4'h5 == state ? plru1_17 : _GEN_2133; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2330 = 4'h5 == state ? plru1_18 : _GEN_2134; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2331 = 4'h5 == state ? plru1_19 : _GEN_2135; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2332 = 4'h5 == state ? plru1_20 : _GEN_2136; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2333 = 4'h5 == state ? plru1_21 : _GEN_2137; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2334 = 4'h5 == state ? plru1_22 : _GEN_2138; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2335 = 4'h5 == state ? plru1_23 : _GEN_2139; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2336 = 4'h5 == state ? plru1_24 : _GEN_2140; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2337 = 4'h5 == state ? plru1_25 : _GEN_2141; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2338 = 4'h5 == state ? plru1_26 : _GEN_2142; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2339 = 4'h5 == state ? plru1_27 : _GEN_2143; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2340 = 4'h5 == state ? plru1_28 : _GEN_2144; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2341 = 4'h5 == state ? plru1_29 : _GEN_2145; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2342 = 4'h5 == state ? plru1_30 : _GEN_2146; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2343 = 4'h5 == state ? plru1_31 : _GEN_2147; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2344 = 4'h5 == state ? plru1_32 : _GEN_2148; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2345 = 4'h5 == state ? plru1_33 : _GEN_2149; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2346 = 4'h5 == state ? plru1_34 : _GEN_2150; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2347 = 4'h5 == state ? plru1_35 : _GEN_2151; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2348 = 4'h5 == state ? plru1_36 : _GEN_2152; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2349 = 4'h5 == state ? plru1_37 : _GEN_2153; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2350 = 4'h5 == state ? plru1_38 : _GEN_2154; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2351 = 4'h5 == state ? plru1_39 : _GEN_2155; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2352 = 4'h5 == state ? plru1_40 : _GEN_2156; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2353 = 4'h5 == state ? plru1_41 : _GEN_2157; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2354 = 4'h5 == state ? plru1_42 : _GEN_2158; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2355 = 4'h5 == state ? plru1_43 : _GEN_2159; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2356 = 4'h5 == state ? plru1_44 : _GEN_2160; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2357 = 4'h5 == state ? plru1_45 : _GEN_2161; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2358 = 4'h5 == state ? plru1_46 : _GEN_2162; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2359 = 4'h5 == state ? plru1_47 : _GEN_2163; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2360 = 4'h5 == state ? plru1_48 : _GEN_2164; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2361 = 4'h5 == state ? plru1_49 : _GEN_2165; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2362 = 4'h5 == state ? plru1_50 : _GEN_2166; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2363 = 4'h5 == state ? plru1_51 : _GEN_2167; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2364 = 4'h5 == state ? plru1_52 : _GEN_2168; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2365 = 4'h5 == state ? plru1_53 : _GEN_2169; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2366 = 4'h5 == state ? plru1_54 : _GEN_2170; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2367 = 4'h5 == state ? plru1_55 : _GEN_2171; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2368 = 4'h5 == state ? plru1_56 : _GEN_2172; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2369 = 4'h5 == state ? plru1_57 : _GEN_2173; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2370 = 4'h5 == state ? plru1_58 : _GEN_2174; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2371 = 4'h5 == state ? plru1_59 : _GEN_2175; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2372 = 4'h5 == state ? plru1_60 : _GEN_2176; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2373 = 4'h5 == state ? plru1_61 : _GEN_2177; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2374 = 4'h5 == state ? plru1_62 : _GEN_2178; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2375 = 4'h5 == state ? plru1_63 : _GEN_2179; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2376 = 4'h5 == state ? plru2_0 : _GEN_2180; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2377 = 4'h5 == state ? plru2_1 : _GEN_2181; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2378 = 4'h5 == state ? plru2_2 : _GEN_2182; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2379 = 4'h5 == state ? plru2_3 : _GEN_2183; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2380 = 4'h5 == state ? plru2_4 : _GEN_2184; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2381 = 4'h5 == state ? plru2_5 : _GEN_2185; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2382 = 4'h5 == state ? plru2_6 : _GEN_2186; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2383 = 4'h5 == state ? plru2_7 : _GEN_2187; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2384 = 4'h5 == state ? plru2_8 : _GEN_2188; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2385 = 4'h5 == state ? plru2_9 : _GEN_2189; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2386 = 4'h5 == state ? plru2_10 : _GEN_2190; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2387 = 4'h5 == state ? plru2_11 : _GEN_2191; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2388 = 4'h5 == state ? plru2_12 : _GEN_2192; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2389 = 4'h5 == state ? plru2_13 : _GEN_2193; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2390 = 4'h5 == state ? plru2_14 : _GEN_2194; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2391 = 4'h5 == state ? plru2_15 : _GEN_2195; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2392 = 4'h5 == state ? plru2_16 : _GEN_2196; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2393 = 4'h5 == state ? plru2_17 : _GEN_2197; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2394 = 4'h5 == state ? plru2_18 : _GEN_2198; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2395 = 4'h5 == state ? plru2_19 : _GEN_2199; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2396 = 4'h5 == state ? plru2_20 : _GEN_2200; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2397 = 4'h5 == state ? plru2_21 : _GEN_2201; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2398 = 4'h5 == state ? plru2_22 : _GEN_2202; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2399 = 4'h5 == state ? plru2_23 : _GEN_2203; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2400 = 4'h5 == state ? plru2_24 : _GEN_2204; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2401 = 4'h5 == state ? plru2_25 : _GEN_2205; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2402 = 4'h5 == state ? plru2_26 : _GEN_2206; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2403 = 4'h5 == state ? plru2_27 : _GEN_2207; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2404 = 4'h5 == state ? plru2_28 : _GEN_2208; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2405 = 4'h5 == state ? plru2_29 : _GEN_2209; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2406 = 4'h5 == state ? plru2_30 : _GEN_2210; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2407 = 4'h5 == state ? plru2_31 : _GEN_2211; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2408 = 4'h5 == state ? plru2_32 : _GEN_2212; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2409 = 4'h5 == state ? plru2_33 : _GEN_2213; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2410 = 4'h5 == state ? plru2_34 : _GEN_2214; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2411 = 4'h5 == state ? plru2_35 : _GEN_2215; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2412 = 4'h5 == state ? plru2_36 : _GEN_2216; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2413 = 4'h5 == state ? plru2_37 : _GEN_2217; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2414 = 4'h5 == state ? plru2_38 : _GEN_2218; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2415 = 4'h5 == state ? plru2_39 : _GEN_2219; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2416 = 4'h5 == state ? plru2_40 : _GEN_2220; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2417 = 4'h5 == state ? plru2_41 : _GEN_2221; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2418 = 4'h5 == state ? plru2_42 : _GEN_2222; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2419 = 4'h5 == state ? plru2_43 : _GEN_2223; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2420 = 4'h5 == state ? plru2_44 : _GEN_2224; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2421 = 4'h5 == state ? plru2_45 : _GEN_2225; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2422 = 4'h5 == state ? plru2_46 : _GEN_2226; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2423 = 4'h5 == state ? plru2_47 : _GEN_2227; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2424 = 4'h5 == state ? plru2_48 : _GEN_2228; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2425 = 4'h5 == state ? plru2_49 : _GEN_2229; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2426 = 4'h5 == state ? plru2_50 : _GEN_2230; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2427 = 4'h5 == state ? plru2_51 : _GEN_2231; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2428 = 4'h5 == state ? plru2_52 : _GEN_2232; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2429 = 4'h5 == state ? plru2_53 : _GEN_2233; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2430 = 4'h5 == state ? plru2_54 : _GEN_2234; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2431 = 4'h5 == state ? plru2_55 : _GEN_2235; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2432 = 4'h5 == state ? plru2_56 : _GEN_2236; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2433 = 4'h5 == state ? plru2_57 : _GEN_2237; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2434 = 4'h5 == state ? plru2_58 : _GEN_2238; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2435 = 4'h5 == state ? plru2_59 : _GEN_2239; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2436 = 4'h5 == state ? plru2_60 : _GEN_2240; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2437 = 4'h5 == state ? plru2_61 : _GEN_2241; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2438 = 4'h5 == state ? plru2_62 : _GEN_2242; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2439 = 4'h5 == state ? plru2_63 : _GEN_2243; // @[Cache.scala 318:18 133:22]
  wire [63:0] _GEN_2440 = 4'h5 == state ? 64'h0 : _GEN_2245; // @[Cache.scala 318:18 289:22]
  wire [3:0] _GEN_2441 = 4'h4 == state ? _GEN_1533 : _GEN_2246; // @[Cache.scala 318:18]
  wire  _GEN_2442 = 4'h4 == state ? _GEN_27 : _GEN_2247; // @[Cache.scala 318:18]
  wire  _GEN_2443 = 4'h4 == state ? plru0_0 : _GEN_2248; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2444 = 4'h4 == state ? plru0_1 : _GEN_2249; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2445 = 4'h4 == state ? plru0_2 : _GEN_2250; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2446 = 4'h4 == state ? plru0_3 : _GEN_2251; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2447 = 4'h4 == state ? plru0_4 : _GEN_2252; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2448 = 4'h4 == state ? plru0_5 : _GEN_2253; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2449 = 4'h4 == state ? plru0_6 : _GEN_2254; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2450 = 4'h4 == state ? plru0_7 : _GEN_2255; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2451 = 4'h4 == state ? plru0_8 : _GEN_2256; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2452 = 4'h4 == state ? plru0_9 : _GEN_2257; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2453 = 4'h4 == state ? plru0_10 : _GEN_2258; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2454 = 4'h4 == state ? plru0_11 : _GEN_2259; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2455 = 4'h4 == state ? plru0_12 : _GEN_2260; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2456 = 4'h4 == state ? plru0_13 : _GEN_2261; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2457 = 4'h4 == state ? plru0_14 : _GEN_2262; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2458 = 4'h4 == state ? plru0_15 : _GEN_2263; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2459 = 4'h4 == state ? plru0_16 : _GEN_2264; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2460 = 4'h4 == state ? plru0_17 : _GEN_2265; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2461 = 4'h4 == state ? plru0_18 : _GEN_2266; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2462 = 4'h4 == state ? plru0_19 : _GEN_2267; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2463 = 4'h4 == state ? plru0_20 : _GEN_2268; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2464 = 4'h4 == state ? plru0_21 : _GEN_2269; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2465 = 4'h4 == state ? plru0_22 : _GEN_2270; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2466 = 4'h4 == state ? plru0_23 : _GEN_2271; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2467 = 4'h4 == state ? plru0_24 : _GEN_2272; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2468 = 4'h4 == state ? plru0_25 : _GEN_2273; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2469 = 4'h4 == state ? plru0_26 : _GEN_2274; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2470 = 4'h4 == state ? plru0_27 : _GEN_2275; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2471 = 4'h4 == state ? plru0_28 : _GEN_2276; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2472 = 4'h4 == state ? plru0_29 : _GEN_2277; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2473 = 4'h4 == state ? plru0_30 : _GEN_2278; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2474 = 4'h4 == state ? plru0_31 : _GEN_2279; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2475 = 4'h4 == state ? plru0_32 : _GEN_2280; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2476 = 4'h4 == state ? plru0_33 : _GEN_2281; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2477 = 4'h4 == state ? plru0_34 : _GEN_2282; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2478 = 4'h4 == state ? plru0_35 : _GEN_2283; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2479 = 4'h4 == state ? plru0_36 : _GEN_2284; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2480 = 4'h4 == state ? plru0_37 : _GEN_2285; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2481 = 4'h4 == state ? plru0_38 : _GEN_2286; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2482 = 4'h4 == state ? plru0_39 : _GEN_2287; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2483 = 4'h4 == state ? plru0_40 : _GEN_2288; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2484 = 4'h4 == state ? plru0_41 : _GEN_2289; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2485 = 4'h4 == state ? plru0_42 : _GEN_2290; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2486 = 4'h4 == state ? plru0_43 : _GEN_2291; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2487 = 4'h4 == state ? plru0_44 : _GEN_2292; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2488 = 4'h4 == state ? plru0_45 : _GEN_2293; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2489 = 4'h4 == state ? plru0_46 : _GEN_2294; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2490 = 4'h4 == state ? plru0_47 : _GEN_2295; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2491 = 4'h4 == state ? plru0_48 : _GEN_2296; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2492 = 4'h4 == state ? plru0_49 : _GEN_2297; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2493 = 4'h4 == state ? plru0_50 : _GEN_2298; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2494 = 4'h4 == state ? plru0_51 : _GEN_2299; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2495 = 4'h4 == state ? plru0_52 : _GEN_2300; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2496 = 4'h4 == state ? plru0_53 : _GEN_2301; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2497 = 4'h4 == state ? plru0_54 : _GEN_2302; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2498 = 4'h4 == state ? plru0_55 : _GEN_2303; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2499 = 4'h4 == state ? plru0_56 : _GEN_2304; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2500 = 4'h4 == state ? plru0_57 : _GEN_2305; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2501 = 4'h4 == state ? plru0_58 : _GEN_2306; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2502 = 4'h4 == state ? plru0_59 : _GEN_2307; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2503 = 4'h4 == state ? plru0_60 : _GEN_2308; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2504 = 4'h4 == state ? plru0_61 : _GEN_2309; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2505 = 4'h4 == state ? plru0_62 : _GEN_2310; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2506 = 4'h4 == state ? plru0_63 : _GEN_2311; // @[Cache.scala 318:18 129:22]
  wire  _GEN_2507 = 4'h4 == state ? plru1_0 : _GEN_2312; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2508 = 4'h4 == state ? plru1_1 : _GEN_2313; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2509 = 4'h4 == state ? plru1_2 : _GEN_2314; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2510 = 4'h4 == state ? plru1_3 : _GEN_2315; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2511 = 4'h4 == state ? plru1_4 : _GEN_2316; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2512 = 4'h4 == state ? plru1_5 : _GEN_2317; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2513 = 4'h4 == state ? plru1_6 : _GEN_2318; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2514 = 4'h4 == state ? plru1_7 : _GEN_2319; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2515 = 4'h4 == state ? plru1_8 : _GEN_2320; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2516 = 4'h4 == state ? plru1_9 : _GEN_2321; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2517 = 4'h4 == state ? plru1_10 : _GEN_2322; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2518 = 4'h4 == state ? plru1_11 : _GEN_2323; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2519 = 4'h4 == state ? plru1_12 : _GEN_2324; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2520 = 4'h4 == state ? plru1_13 : _GEN_2325; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2521 = 4'h4 == state ? plru1_14 : _GEN_2326; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2522 = 4'h4 == state ? plru1_15 : _GEN_2327; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2523 = 4'h4 == state ? plru1_16 : _GEN_2328; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2524 = 4'h4 == state ? plru1_17 : _GEN_2329; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2525 = 4'h4 == state ? plru1_18 : _GEN_2330; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2526 = 4'h4 == state ? plru1_19 : _GEN_2331; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2527 = 4'h4 == state ? plru1_20 : _GEN_2332; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2528 = 4'h4 == state ? plru1_21 : _GEN_2333; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2529 = 4'h4 == state ? plru1_22 : _GEN_2334; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2530 = 4'h4 == state ? plru1_23 : _GEN_2335; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2531 = 4'h4 == state ? plru1_24 : _GEN_2336; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2532 = 4'h4 == state ? plru1_25 : _GEN_2337; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2533 = 4'h4 == state ? plru1_26 : _GEN_2338; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2534 = 4'h4 == state ? plru1_27 : _GEN_2339; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2535 = 4'h4 == state ? plru1_28 : _GEN_2340; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2536 = 4'h4 == state ? plru1_29 : _GEN_2341; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2537 = 4'h4 == state ? plru1_30 : _GEN_2342; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2538 = 4'h4 == state ? plru1_31 : _GEN_2343; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2539 = 4'h4 == state ? plru1_32 : _GEN_2344; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2540 = 4'h4 == state ? plru1_33 : _GEN_2345; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2541 = 4'h4 == state ? plru1_34 : _GEN_2346; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2542 = 4'h4 == state ? plru1_35 : _GEN_2347; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2543 = 4'h4 == state ? plru1_36 : _GEN_2348; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2544 = 4'h4 == state ? plru1_37 : _GEN_2349; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2545 = 4'h4 == state ? plru1_38 : _GEN_2350; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2546 = 4'h4 == state ? plru1_39 : _GEN_2351; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2547 = 4'h4 == state ? plru1_40 : _GEN_2352; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2548 = 4'h4 == state ? plru1_41 : _GEN_2353; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2549 = 4'h4 == state ? plru1_42 : _GEN_2354; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2550 = 4'h4 == state ? plru1_43 : _GEN_2355; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2551 = 4'h4 == state ? plru1_44 : _GEN_2356; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2552 = 4'h4 == state ? plru1_45 : _GEN_2357; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2553 = 4'h4 == state ? plru1_46 : _GEN_2358; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2554 = 4'h4 == state ? plru1_47 : _GEN_2359; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2555 = 4'h4 == state ? plru1_48 : _GEN_2360; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2556 = 4'h4 == state ? plru1_49 : _GEN_2361; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2557 = 4'h4 == state ? plru1_50 : _GEN_2362; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2558 = 4'h4 == state ? plru1_51 : _GEN_2363; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2559 = 4'h4 == state ? plru1_52 : _GEN_2364; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2560 = 4'h4 == state ? plru1_53 : _GEN_2365; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2561 = 4'h4 == state ? plru1_54 : _GEN_2366; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2562 = 4'h4 == state ? plru1_55 : _GEN_2367; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2563 = 4'h4 == state ? plru1_56 : _GEN_2368; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2564 = 4'h4 == state ? plru1_57 : _GEN_2369; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2565 = 4'h4 == state ? plru1_58 : _GEN_2370; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2566 = 4'h4 == state ? plru1_59 : _GEN_2371; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2567 = 4'h4 == state ? plru1_60 : _GEN_2372; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2568 = 4'h4 == state ? plru1_61 : _GEN_2373; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2569 = 4'h4 == state ? plru1_62 : _GEN_2374; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2570 = 4'h4 == state ? plru1_63 : _GEN_2375; // @[Cache.scala 318:18 131:22]
  wire  _GEN_2571 = 4'h4 == state ? plru2_0 : _GEN_2376; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2572 = 4'h4 == state ? plru2_1 : _GEN_2377; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2573 = 4'h4 == state ? plru2_2 : _GEN_2378; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2574 = 4'h4 == state ? plru2_3 : _GEN_2379; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2575 = 4'h4 == state ? plru2_4 : _GEN_2380; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2576 = 4'h4 == state ? plru2_5 : _GEN_2381; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2577 = 4'h4 == state ? plru2_6 : _GEN_2382; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2578 = 4'h4 == state ? plru2_7 : _GEN_2383; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2579 = 4'h4 == state ? plru2_8 : _GEN_2384; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2580 = 4'h4 == state ? plru2_9 : _GEN_2385; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2581 = 4'h4 == state ? plru2_10 : _GEN_2386; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2582 = 4'h4 == state ? plru2_11 : _GEN_2387; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2583 = 4'h4 == state ? plru2_12 : _GEN_2388; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2584 = 4'h4 == state ? plru2_13 : _GEN_2389; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2585 = 4'h4 == state ? plru2_14 : _GEN_2390; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2586 = 4'h4 == state ? plru2_15 : _GEN_2391; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2587 = 4'h4 == state ? plru2_16 : _GEN_2392; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2588 = 4'h4 == state ? plru2_17 : _GEN_2393; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2589 = 4'h4 == state ? plru2_18 : _GEN_2394; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2590 = 4'h4 == state ? plru2_19 : _GEN_2395; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2591 = 4'h4 == state ? plru2_20 : _GEN_2396; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2592 = 4'h4 == state ? plru2_21 : _GEN_2397; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2593 = 4'h4 == state ? plru2_22 : _GEN_2398; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2594 = 4'h4 == state ? plru2_23 : _GEN_2399; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2595 = 4'h4 == state ? plru2_24 : _GEN_2400; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2596 = 4'h4 == state ? plru2_25 : _GEN_2401; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2597 = 4'h4 == state ? plru2_26 : _GEN_2402; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2598 = 4'h4 == state ? plru2_27 : _GEN_2403; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2599 = 4'h4 == state ? plru2_28 : _GEN_2404; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2600 = 4'h4 == state ? plru2_29 : _GEN_2405; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2601 = 4'h4 == state ? plru2_30 : _GEN_2406; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2602 = 4'h4 == state ? plru2_31 : _GEN_2407; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2603 = 4'h4 == state ? plru2_32 : _GEN_2408; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2604 = 4'h4 == state ? plru2_33 : _GEN_2409; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2605 = 4'h4 == state ? plru2_34 : _GEN_2410; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2606 = 4'h4 == state ? plru2_35 : _GEN_2411; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2607 = 4'h4 == state ? plru2_36 : _GEN_2412; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2608 = 4'h4 == state ? plru2_37 : _GEN_2413; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2609 = 4'h4 == state ? plru2_38 : _GEN_2414; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2610 = 4'h4 == state ? plru2_39 : _GEN_2415; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2611 = 4'h4 == state ? plru2_40 : _GEN_2416; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2612 = 4'h4 == state ? plru2_41 : _GEN_2417; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2613 = 4'h4 == state ? plru2_42 : _GEN_2418; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2614 = 4'h4 == state ? plru2_43 : _GEN_2419; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2615 = 4'h4 == state ? plru2_44 : _GEN_2420; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2616 = 4'h4 == state ? plru2_45 : _GEN_2421; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2617 = 4'h4 == state ? plru2_46 : _GEN_2422; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2618 = 4'h4 == state ? plru2_47 : _GEN_2423; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2619 = 4'h4 == state ? plru2_48 : _GEN_2424; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2620 = 4'h4 == state ? plru2_49 : _GEN_2425; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2621 = 4'h4 == state ? plru2_50 : _GEN_2426; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2622 = 4'h4 == state ? plru2_51 : _GEN_2427; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2623 = 4'h4 == state ? plru2_52 : _GEN_2428; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2624 = 4'h4 == state ? plru2_53 : _GEN_2429; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2625 = 4'h4 == state ? plru2_54 : _GEN_2430; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2626 = 4'h4 == state ? plru2_55 : _GEN_2431; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2627 = 4'h4 == state ? plru2_56 : _GEN_2432; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2628 = 4'h4 == state ? plru2_57 : _GEN_2433; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2629 = 4'h4 == state ? plru2_58 : _GEN_2434; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2630 = 4'h4 == state ? plru2_59 : _GEN_2435; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2631 = 4'h4 == state ? plru2_60 : _GEN_2436; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2632 = 4'h4 == state ? plru2_61 : _GEN_2437; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2633 = 4'h4 == state ? plru2_62 : _GEN_2438; // @[Cache.scala 318:18 133:22]
  wire  _GEN_2634 = 4'h4 == state ? plru2_63 : _GEN_2439; // @[Cache.scala 318:18 133:22]
  wire [63:0] _GEN_2635 = 4'h4 == state ? 64'h0 : _GEN_2440; // @[Cache.scala 318:18 289:22]
  wire  _GEN_2636 = 4'h3 == state ? _GEN_993 : pipeline_ready; // @[Cache.scala 318:18]
  wire [5:0] _GEN_2638 = 4'h3 == state ? _GEN_995 : _GEN_3; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2639 = 4'h3 == state ? _GEN_996 : 128'h0; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2640 = 4'h3 == state ? _GEN_997 : 21'h0; // @[Cache.scala 114:16 318:18]
  wire  _GEN_2642 = 4'h3 == state ? _GEN_1000 : pipeline_ready; // @[Cache.scala 318:18]
  wire [5:0] _GEN_2644 = 4'h3 == state ? _GEN_1002 : _GEN_3; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2645 = 4'h3 == state ? _GEN_1003 : 128'h0; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2646 = 4'h3 == state ? _GEN_1004 : 21'h0; // @[Cache.scala 114:16 318:18]
  wire  _GEN_2648 = 4'h3 == state ? _GEN_1007 : pipeline_ready; // @[Cache.scala 318:18]
  wire [5:0] _GEN_2650 = 4'h3 == state ? _GEN_1009 : _GEN_3; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2651 = 4'h3 == state ? _GEN_1010 : 128'h0; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2652 = 4'h3 == state ? _GEN_1011 : 21'h0; // @[Cache.scala 114:16 318:18]
  wire  _GEN_2654 = 4'h3 == state ? _GEN_1014 : pipeline_ready; // @[Cache.scala 318:18]
  wire [5:0] _GEN_2656 = 4'h3 == state ? _GEN_1016 : _GEN_3; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2657 = 4'h3 == state ? _GEN_1017 : 128'h0; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2658 = 4'h3 == state ? _GEN_1018 : 21'h0; // @[Cache.scala 114:16 318:18]
  wire [3:0] _GEN_2660 = 4'h3 == state ? _GEN_1340 : _GEN_2441; // @[Cache.scala 318:18]
  wire  _GEN_2661 = 4'h3 == state ? _GEN_1341 : _GEN_2443; // @[Cache.scala 318:18]
  wire  _GEN_2662 = 4'h3 == state ? _GEN_1342 : _GEN_2444; // @[Cache.scala 318:18]
  wire  _GEN_2663 = 4'h3 == state ? _GEN_1343 : _GEN_2445; // @[Cache.scala 318:18]
  wire  _GEN_2664 = 4'h3 == state ? _GEN_1344 : _GEN_2446; // @[Cache.scala 318:18]
  wire  _GEN_2665 = 4'h3 == state ? _GEN_1345 : _GEN_2447; // @[Cache.scala 318:18]
  wire  _GEN_2666 = 4'h3 == state ? _GEN_1346 : _GEN_2448; // @[Cache.scala 318:18]
  wire  _GEN_2667 = 4'h3 == state ? _GEN_1347 : _GEN_2449; // @[Cache.scala 318:18]
  wire  _GEN_2668 = 4'h3 == state ? _GEN_1348 : _GEN_2450; // @[Cache.scala 318:18]
  wire  _GEN_2669 = 4'h3 == state ? _GEN_1349 : _GEN_2451; // @[Cache.scala 318:18]
  wire  _GEN_2670 = 4'h3 == state ? _GEN_1350 : _GEN_2452; // @[Cache.scala 318:18]
  wire  _GEN_2671 = 4'h3 == state ? _GEN_1351 : _GEN_2453; // @[Cache.scala 318:18]
  wire  _GEN_2672 = 4'h3 == state ? _GEN_1352 : _GEN_2454; // @[Cache.scala 318:18]
  wire  _GEN_2673 = 4'h3 == state ? _GEN_1353 : _GEN_2455; // @[Cache.scala 318:18]
  wire  _GEN_2674 = 4'h3 == state ? _GEN_1354 : _GEN_2456; // @[Cache.scala 318:18]
  wire  _GEN_2675 = 4'h3 == state ? _GEN_1355 : _GEN_2457; // @[Cache.scala 318:18]
  wire  _GEN_2676 = 4'h3 == state ? _GEN_1356 : _GEN_2458; // @[Cache.scala 318:18]
  wire  _GEN_2677 = 4'h3 == state ? _GEN_1357 : _GEN_2459; // @[Cache.scala 318:18]
  wire  _GEN_2678 = 4'h3 == state ? _GEN_1358 : _GEN_2460; // @[Cache.scala 318:18]
  wire  _GEN_2679 = 4'h3 == state ? _GEN_1359 : _GEN_2461; // @[Cache.scala 318:18]
  wire  _GEN_2680 = 4'h3 == state ? _GEN_1360 : _GEN_2462; // @[Cache.scala 318:18]
  wire  _GEN_2681 = 4'h3 == state ? _GEN_1361 : _GEN_2463; // @[Cache.scala 318:18]
  wire  _GEN_2682 = 4'h3 == state ? _GEN_1362 : _GEN_2464; // @[Cache.scala 318:18]
  wire  _GEN_2683 = 4'h3 == state ? _GEN_1363 : _GEN_2465; // @[Cache.scala 318:18]
  wire  _GEN_2684 = 4'h3 == state ? _GEN_1364 : _GEN_2466; // @[Cache.scala 318:18]
  wire  _GEN_2685 = 4'h3 == state ? _GEN_1365 : _GEN_2467; // @[Cache.scala 318:18]
  wire  _GEN_2686 = 4'h3 == state ? _GEN_1366 : _GEN_2468; // @[Cache.scala 318:18]
  wire  _GEN_2687 = 4'h3 == state ? _GEN_1367 : _GEN_2469; // @[Cache.scala 318:18]
  wire  _GEN_2688 = 4'h3 == state ? _GEN_1368 : _GEN_2470; // @[Cache.scala 318:18]
  wire  _GEN_2689 = 4'h3 == state ? _GEN_1369 : _GEN_2471; // @[Cache.scala 318:18]
  wire  _GEN_2690 = 4'h3 == state ? _GEN_1370 : _GEN_2472; // @[Cache.scala 318:18]
  wire  _GEN_2691 = 4'h3 == state ? _GEN_1371 : _GEN_2473; // @[Cache.scala 318:18]
  wire  _GEN_2692 = 4'h3 == state ? _GEN_1372 : _GEN_2474; // @[Cache.scala 318:18]
  wire  _GEN_2693 = 4'h3 == state ? _GEN_1373 : _GEN_2475; // @[Cache.scala 318:18]
  wire  _GEN_2694 = 4'h3 == state ? _GEN_1374 : _GEN_2476; // @[Cache.scala 318:18]
  wire  _GEN_2695 = 4'h3 == state ? _GEN_1375 : _GEN_2477; // @[Cache.scala 318:18]
  wire  _GEN_2696 = 4'h3 == state ? _GEN_1376 : _GEN_2478; // @[Cache.scala 318:18]
  wire  _GEN_2697 = 4'h3 == state ? _GEN_1377 : _GEN_2479; // @[Cache.scala 318:18]
  wire  _GEN_2698 = 4'h3 == state ? _GEN_1378 : _GEN_2480; // @[Cache.scala 318:18]
  wire  _GEN_2699 = 4'h3 == state ? _GEN_1379 : _GEN_2481; // @[Cache.scala 318:18]
  wire  _GEN_2700 = 4'h3 == state ? _GEN_1380 : _GEN_2482; // @[Cache.scala 318:18]
  wire  _GEN_2701 = 4'h3 == state ? _GEN_1381 : _GEN_2483; // @[Cache.scala 318:18]
  wire  _GEN_2702 = 4'h3 == state ? _GEN_1382 : _GEN_2484; // @[Cache.scala 318:18]
  wire  _GEN_2703 = 4'h3 == state ? _GEN_1383 : _GEN_2485; // @[Cache.scala 318:18]
  wire  _GEN_2704 = 4'h3 == state ? _GEN_1384 : _GEN_2486; // @[Cache.scala 318:18]
  wire  _GEN_2705 = 4'h3 == state ? _GEN_1385 : _GEN_2487; // @[Cache.scala 318:18]
  wire  _GEN_2706 = 4'h3 == state ? _GEN_1386 : _GEN_2488; // @[Cache.scala 318:18]
  wire  _GEN_2707 = 4'h3 == state ? _GEN_1387 : _GEN_2489; // @[Cache.scala 318:18]
  wire  _GEN_2708 = 4'h3 == state ? _GEN_1388 : _GEN_2490; // @[Cache.scala 318:18]
  wire  _GEN_2709 = 4'h3 == state ? _GEN_1389 : _GEN_2491; // @[Cache.scala 318:18]
  wire  _GEN_2710 = 4'h3 == state ? _GEN_1390 : _GEN_2492; // @[Cache.scala 318:18]
  wire  _GEN_2711 = 4'h3 == state ? _GEN_1391 : _GEN_2493; // @[Cache.scala 318:18]
  wire  _GEN_2712 = 4'h3 == state ? _GEN_1392 : _GEN_2494; // @[Cache.scala 318:18]
  wire  _GEN_2713 = 4'h3 == state ? _GEN_1393 : _GEN_2495; // @[Cache.scala 318:18]
  wire  _GEN_2714 = 4'h3 == state ? _GEN_1394 : _GEN_2496; // @[Cache.scala 318:18]
  wire  _GEN_2715 = 4'h3 == state ? _GEN_1395 : _GEN_2497; // @[Cache.scala 318:18]
  wire  _GEN_2716 = 4'h3 == state ? _GEN_1396 : _GEN_2498; // @[Cache.scala 318:18]
  wire  _GEN_2717 = 4'h3 == state ? _GEN_1397 : _GEN_2499; // @[Cache.scala 318:18]
  wire  _GEN_2718 = 4'h3 == state ? _GEN_1398 : _GEN_2500; // @[Cache.scala 318:18]
  wire  _GEN_2719 = 4'h3 == state ? _GEN_1399 : _GEN_2501; // @[Cache.scala 318:18]
  wire  _GEN_2720 = 4'h3 == state ? _GEN_1400 : _GEN_2502; // @[Cache.scala 318:18]
  wire  _GEN_2721 = 4'h3 == state ? _GEN_1401 : _GEN_2503; // @[Cache.scala 318:18]
  wire  _GEN_2722 = 4'h3 == state ? _GEN_1402 : _GEN_2504; // @[Cache.scala 318:18]
  wire  _GEN_2723 = 4'h3 == state ? _GEN_1403 : _GEN_2505; // @[Cache.scala 318:18]
  wire  _GEN_2724 = 4'h3 == state ? _GEN_1404 : _GEN_2506; // @[Cache.scala 318:18]
  wire  _GEN_2725 = 4'h3 == state ? _GEN_1405 : _GEN_2507; // @[Cache.scala 318:18]
  wire  _GEN_2726 = 4'h3 == state ? _GEN_1406 : _GEN_2508; // @[Cache.scala 318:18]
  wire  _GEN_2727 = 4'h3 == state ? _GEN_1407 : _GEN_2509; // @[Cache.scala 318:18]
  wire  _GEN_2728 = 4'h3 == state ? _GEN_1408 : _GEN_2510; // @[Cache.scala 318:18]
  wire  _GEN_2729 = 4'h3 == state ? _GEN_1409 : _GEN_2511; // @[Cache.scala 318:18]
  wire  _GEN_2730 = 4'h3 == state ? _GEN_1410 : _GEN_2512; // @[Cache.scala 318:18]
  wire  _GEN_2731 = 4'h3 == state ? _GEN_1411 : _GEN_2513; // @[Cache.scala 318:18]
  wire  _GEN_2732 = 4'h3 == state ? _GEN_1412 : _GEN_2514; // @[Cache.scala 318:18]
  wire  _GEN_2733 = 4'h3 == state ? _GEN_1413 : _GEN_2515; // @[Cache.scala 318:18]
  wire  _GEN_2734 = 4'h3 == state ? _GEN_1414 : _GEN_2516; // @[Cache.scala 318:18]
  wire  _GEN_2735 = 4'h3 == state ? _GEN_1415 : _GEN_2517; // @[Cache.scala 318:18]
  wire  _GEN_2736 = 4'h3 == state ? _GEN_1416 : _GEN_2518; // @[Cache.scala 318:18]
  wire  _GEN_2737 = 4'h3 == state ? _GEN_1417 : _GEN_2519; // @[Cache.scala 318:18]
  wire  _GEN_2738 = 4'h3 == state ? _GEN_1418 : _GEN_2520; // @[Cache.scala 318:18]
  wire  _GEN_2739 = 4'h3 == state ? _GEN_1419 : _GEN_2521; // @[Cache.scala 318:18]
  wire  _GEN_2740 = 4'h3 == state ? _GEN_1420 : _GEN_2522; // @[Cache.scala 318:18]
  wire  _GEN_2741 = 4'h3 == state ? _GEN_1421 : _GEN_2523; // @[Cache.scala 318:18]
  wire  _GEN_2742 = 4'h3 == state ? _GEN_1422 : _GEN_2524; // @[Cache.scala 318:18]
  wire  _GEN_2743 = 4'h3 == state ? _GEN_1423 : _GEN_2525; // @[Cache.scala 318:18]
  wire  _GEN_2744 = 4'h3 == state ? _GEN_1424 : _GEN_2526; // @[Cache.scala 318:18]
  wire  _GEN_2745 = 4'h3 == state ? _GEN_1425 : _GEN_2527; // @[Cache.scala 318:18]
  wire  _GEN_2746 = 4'h3 == state ? _GEN_1426 : _GEN_2528; // @[Cache.scala 318:18]
  wire  _GEN_2747 = 4'h3 == state ? _GEN_1427 : _GEN_2529; // @[Cache.scala 318:18]
  wire  _GEN_2748 = 4'h3 == state ? _GEN_1428 : _GEN_2530; // @[Cache.scala 318:18]
  wire  _GEN_2749 = 4'h3 == state ? _GEN_1429 : _GEN_2531; // @[Cache.scala 318:18]
  wire  _GEN_2750 = 4'h3 == state ? _GEN_1430 : _GEN_2532; // @[Cache.scala 318:18]
  wire  _GEN_2751 = 4'h3 == state ? _GEN_1431 : _GEN_2533; // @[Cache.scala 318:18]
  wire  _GEN_2752 = 4'h3 == state ? _GEN_1432 : _GEN_2534; // @[Cache.scala 318:18]
  wire  _GEN_2753 = 4'h3 == state ? _GEN_1433 : _GEN_2535; // @[Cache.scala 318:18]
  wire  _GEN_2754 = 4'h3 == state ? _GEN_1434 : _GEN_2536; // @[Cache.scala 318:18]
  wire  _GEN_2755 = 4'h3 == state ? _GEN_1435 : _GEN_2537; // @[Cache.scala 318:18]
  wire  _GEN_2756 = 4'h3 == state ? _GEN_1436 : _GEN_2538; // @[Cache.scala 318:18]
  wire  _GEN_2757 = 4'h3 == state ? _GEN_1437 : _GEN_2539; // @[Cache.scala 318:18]
  wire  _GEN_2758 = 4'h3 == state ? _GEN_1438 : _GEN_2540; // @[Cache.scala 318:18]
  wire  _GEN_2759 = 4'h3 == state ? _GEN_1439 : _GEN_2541; // @[Cache.scala 318:18]
  wire  _GEN_2760 = 4'h3 == state ? _GEN_1440 : _GEN_2542; // @[Cache.scala 318:18]
  wire  _GEN_2761 = 4'h3 == state ? _GEN_1441 : _GEN_2543; // @[Cache.scala 318:18]
  wire  _GEN_2762 = 4'h3 == state ? _GEN_1442 : _GEN_2544; // @[Cache.scala 318:18]
  wire  _GEN_2763 = 4'h3 == state ? _GEN_1443 : _GEN_2545; // @[Cache.scala 318:18]
  wire  _GEN_2764 = 4'h3 == state ? _GEN_1444 : _GEN_2546; // @[Cache.scala 318:18]
  wire  _GEN_2765 = 4'h3 == state ? _GEN_1445 : _GEN_2547; // @[Cache.scala 318:18]
  wire  _GEN_2766 = 4'h3 == state ? _GEN_1446 : _GEN_2548; // @[Cache.scala 318:18]
  wire  _GEN_2767 = 4'h3 == state ? _GEN_1447 : _GEN_2549; // @[Cache.scala 318:18]
  wire  _GEN_2768 = 4'h3 == state ? _GEN_1448 : _GEN_2550; // @[Cache.scala 318:18]
  wire  _GEN_2769 = 4'h3 == state ? _GEN_1449 : _GEN_2551; // @[Cache.scala 318:18]
  wire  _GEN_2770 = 4'h3 == state ? _GEN_1450 : _GEN_2552; // @[Cache.scala 318:18]
  wire  _GEN_2771 = 4'h3 == state ? _GEN_1451 : _GEN_2553; // @[Cache.scala 318:18]
  wire  _GEN_2772 = 4'h3 == state ? _GEN_1452 : _GEN_2554; // @[Cache.scala 318:18]
  wire  _GEN_2773 = 4'h3 == state ? _GEN_1453 : _GEN_2555; // @[Cache.scala 318:18]
  wire  _GEN_2774 = 4'h3 == state ? _GEN_1454 : _GEN_2556; // @[Cache.scala 318:18]
  wire  _GEN_2775 = 4'h3 == state ? _GEN_1455 : _GEN_2557; // @[Cache.scala 318:18]
  wire  _GEN_2776 = 4'h3 == state ? _GEN_1456 : _GEN_2558; // @[Cache.scala 318:18]
  wire  _GEN_2777 = 4'h3 == state ? _GEN_1457 : _GEN_2559; // @[Cache.scala 318:18]
  wire  _GEN_2778 = 4'h3 == state ? _GEN_1458 : _GEN_2560; // @[Cache.scala 318:18]
  wire  _GEN_2779 = 4'h3 == state ? _GEN_1459 : _GEN_2561; // @[Cache.scala 318:18]
  wire  _GEN_2780 = 4'h3 == state ? _GEN_1460 : _GEN_2562; // @[Cache.scala 318:18]
  wire  _GEN_2781 = 4'h3 == state ? _GEN_1461 : _GEN_2563; // @[Cache.scala 318:18]
  wire  _GEN_2782 = 4'h3 == state ? _GEN_1462 : _GEN_2564; // @[Cache.scala 318:18]
  wire  _GEN_2783 = 4'h3 == state ? _GEN_1463 : _GEN_2565; // @[Cache.scala 318:18]
  wire  _GEN_2784 = 4'h3 == state ? _GEN_1464 : _GEN_2566; // @[Cache.scala 318:18]
  wire  _GEN_2785 = 4'h3 == state ? _GEN_1465 : _GEN_2567; // @[Cache.scala 318:18]
  wire  _GEN_2786 = 4'h3 == state ? _GEN_1466 : _GEN_2568; // @[Cache.scala 318:18]
  wire  _GEN_2787 = 4'h3 == state ? _GEN_1467 : _GEN_2569; // @[Cache.scala 318:18]
  wire  _GEN_2788 = 4'h3 == state ? _GEN_1468 : _GEN_2570; // @[Cache.scala 318:18]
  wire  _GEN_2789 = 4'h3 == state ? _GEN_1469 : _GEN_2571; // @[Cache.scala 318:18]
  wire  _GEN_2790 = 4'h3 == state ? _GEN_1470 : _GEN_2572; // @[Cache.scala 318:18]
  wire  _GEN_2791 = 4'h3 == state ? _GEN_1471 : _GEN_2573; // @[Cache.scala 318:18]
  wire  _GEN_2792 = 4'h3 == state ? _GEN_1472 : _GEN_2574; // @[Cache.scala 318:18]
  wire  _GEN_2793 = 4'h3 == state ? _GEN_1473 : _GEN_2575; // @[Cache.scala 318:18]
  wire  _GEN_2794 = 4'h3 == state ? _GEN_1474 : _GEN_2576; // @[Cache.scala 318:18]
  wire  _GEN_2795 = 4'h3 == state ? _GEN_1475 : _GEN_2577; // @[Cache.scala 318:18]
  wire  _GEN_2796 = 4'h3 == state ? _GEN_1476 : _GEN_2578; // @[Cache.scala 318:18]
  wire  _GEN_2797 = 4'h3 == state ? _GEN_1477 : _GEN_2579; // @[Cache.scala 318:18]
  wire  _GEN_2798 = 4'h3 == state ? _GEN_1478 : _GEN_2580; // @[Cache.scala 318:18]
  wire  _GEN_2799 = 4'h3 == state ? _GEN_1479 : _GEN_2581; // @[Cache.scala 318:18]
  wire  _GEN_2800 = 4'h3 == state ? _GEN_1480 : _GEN_2582; // @[Cache.scala 318:18]
  wire  _GEN_2801 = 4'h3 == state ? _GEN_1481 : _GEN_2583; // @[Cache.scala 318:18]
  wire  _GEN_2802 = 4'h3 == state ? _GEN_1482 : _GEN_2584; // @[Cache.scala 318:18]
  wire  _GEN_2803 = 4'h3 == state ? _GEN_1483 : _GEN_2585; // @[Cache.scala 318:18]
  wire  _GEN_2804 = 4'h3 == state ? _GEN_1484 : _GEN_2586; // @[Cache.scala 318:18]
  wire  _GEN_2805 = 4'h3 == state ? _GEN_1485 : _GEN_2587; // @[Cache.scala 318:18]
  wire  _GEN_2806 = 4'h3 == state ? _GEN_1486 : _GEN_2588; // @[Cache.scala 318:18]
  wire  _GEN_2807 = 4'h3 == state ? _GEN_1487 : _GEN_2589; // @[Cache.scala 318:18]
  wire  _GEN_2808 = 4'h3 == state ? _GEN_1488 : _GEN_2590; // @[Cache.scala 318:18]
  wire  _GEN_2809 = 4'h3 == state ? _GEN_1489 : _GEN_2591; // @[Cache.scala 318:18]
  wire  _GEN_2810 = 4'h3 == state ? _GEN_1490 : _GEN_2592; // @[Cache.scala 318:18]
  wire  _GEN_2811 = 4'h3 == state ? _GEN_1491 : _GEN_2593; // @[Cache.scala 318:18]
  wire  _GEN_2812 = 4'h3 == state ? _GEN_1492 : _GEN_2594; // @[Cache.scala 318:18]
  wire  _GEN_2813 = 4'h3 == state ? _GEN_1493 : _GEN_2595; // @[Cache.scala 318:18]
  wire  _GEN_2814 = 4'h3 == state ? _GEN_1494 : _GEN_2596; // @[Cache.scala 318:18]
  wire  _GEN_2815 = 4'h3 == state ? _GEN_1495 : _GEN_2597; // @[Cache.scala 318:18]
  wire  _GEN_2816 = 4'h3 == state ? _GEN_1496 : _GEN_2598; // @[Cache.scala 318:18]
  wire  _GEN_2817 = 4'h3 == state ? _GEN_1497 : _GEN_2599; // @[Cache.scala 318:18]
  wire  _GEN_2818 = 4'h3 == state ? _GEN_1498 : _GEN_2600; // @[Cache.scala 318:18]
  wire  _GEN_2819 = 4'h3 == state ? _GEN_1499 : _GEN_2601; // @[Cache.scala 318:18]
  wire  _GEN_2820 = 4'h3 == state ? _GEN_1500 : _GEN_2602; // @[Cache.scala 318:18]
  wire  _GEN_2821 = 4'h3 == state ? _GEN_1501 : _GEN_2603; // @[Cache.scala 318:18]
  wire  _GEN_2822 = 4'h3 == state ? _GEN_1502 : _GEN_2604; // @[Cache.scala 318:18]
  wire  _GEN_2823 = 4'h3 == state ? _GEN_1503 : _GEN_2605; // @[Cache.scala 318:18]
  wire  _GEN_2824 = 4'h3 == state ? _GEN_1504 : _GEN_2606; // @[Cache.scala 318:18]
  wire  _GEN_2825 = 4'h3 == state ? _GEN_1505 : _GEN_2607; // @[Cache.scala 318:18]
  wire  _GEN_2826 = 4'h3 == state ? _GEN_1506 : _GEN_2608; // @[Cache.scala 318:18]
  wire  _GEN_2827 = 4'h3 == state ? _GEN_1507 : _GEN_2609; // @[Cache.scala 318:18]
  wire  _GEN_2828 = 4'h3 == state ? _GEN_1508 : _GEN_2610; // @[Cache.scala 318:18]
  wire  _GEN_2829 = 4'h3 == state ? _GEN_1509 : _GEN_2611; // @[Cache.scala 318:18]
  wire  _GEN_2830 = 4'h3 == state ? _GEN_1510 : _GEN_2612; // @[Cache.scala 318:18]
  wire  _GEN_2831 = 4'h3 == state ? _GEN_1511 : _GEN_2613; // @[Cache.scala 318:18]
  wire  _GEN_2832 = 4'h3 == state ? _GEN_1512 : _GEN_2614; // @[Cache.scala 318:18]
  wire  _GEN_2833 = 4'h3 == state ? _GEN_1513 : _GEN_2615; // @[Cache.scala 318:18]
  wire  _GEN_2834 = 4'h3 == state ? _GEN_1514 : _GEN_2616; // @[Cache.scala 318:18]
  wire  _GEN_2835 = 4'h3 == state ? _GEN_1515 : _GEN_2617; // @[Cache.scala 318:18]
  wire  _GEN_2836 = 4'h3 == state ? _GEN_1516 : _GEN_2618; // @[Cache.scala 318:18]
  wire  _GEN_2837 = 4'h3 == state ? _GEN_1517 : _GEN_2619; // @[Cache.scala 318:18]
  wire  _GEN_2838 = 4'h3 == state ? _GEN_1518 : _GEN_2620; // @[Cache.scala 318:18]
  wire  _GEN_2839 = 4'h3 == state ? _GEN_1519 : _GEN_2621; // @[Cache.scala 318:18]
  wire  _GEN_2840 = 4'h3 == state ? _GEN_1520 : _GEN_2622; // @[Cache.scala 318:18]
  wire  _GEN_2841 = 4'h3 == state ? _GEN_1521 : _GEN_2623; // @[Cache.scala 318:18]
  wire  _GEN_2842 = 4'h3 == state ? _GEN_1522 : _GEN_2624; // @[Cache.scala 318:18]
  wire  _GEN_2843 = 4'h3 == state ? _GEN_1523 : _GEN_2625; // @[Cache.scala 318:18]
  wire  _GEN_2844 = 4'h3 == state ? _GEN_1524 : _GEN_2626; // @[Cache.scala 318:18]
  wire  _GEN_2845 = 4'h3 == state ? _GEN_1525 : _GEN_2627; // @[Cache.scala 318:18]
  wire  _GEN_2846 = 4'h3 == state ? _GEN_1526 : _GEN_2628; // @[Cache.scala 318:18]
  wire  _GEN_2847 = 4'h3 == state ? _GEN_1527 : _GEN_2629; // @[Cache.scala 318:18]
  wire  _GEN_2848 = 4'h3 == state ? _GEN_1528 : _GEN_2630; // @[Cache.scala 318:18]
  wire  _GEN_2849 = 4'h3 == state ? _GEN_1529 : _GEN_2631; // @[Cache.scala 318:18]
  wire  _GEN_2850 = 4'h3 == state ? _GEN_1530 : _GEN_2632; // @[Cache.scala 318:18]
  wire  _GEN_2851 = 4'h3 == state ? _GEN_1531 : _GEN_2633; // @[Cache.scala 318:18]
  wire  _GEN_2852 = 4'h3 == state ? _GEN_1532 : _GEN_2634; // @[Cache.scala 318:18]
  wire  _GEN_2853 = 4'h3 == state ? _GEN_27 : _GEN_2442; // @[Cache.scala 318:18]
  wire [63:0] _GEN_2854 = 4'h3 == state ? 64'h0 : _GEN_2635; // @[Cache.scala 318:18 289:22]
  wire [3:0] _GEN_2857 = 4'h2 == state ? _GEN_991 : _GEN_2660; // @[Cache.scala 318:18]
  wire  _GEN_2858 = 4'h2 == state ? pipeline_ready : _GEN_2636; // @[Cache.scala 318:18]
  wire  _GEN_2859 = 4'h2 == state ? 1'h0 : 4'h3 == state & _T_325; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_2860 = 4'h2 == state ? _GEN_3 : _GEN_2638; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2861 = 4'h2 == state ? 128'h0 : _GEN_2639; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2862 = 4'h2 == state ? 21'h0 : _GEN_2640; // @[Cache.scala 114:16 318:18]
  wire  _GEN_2863 = 4'h2 == state ? 1'h0 : 4'h3 == state & _GEN_998; // @[Cache.scala 116:18 318:18]
  wire  _GEN_2864 = 4'h2 == state ? pipeline_ready : _GEN_2642; // @[Cache.scala 318:18]
  wire  _GEN_2865 = 4'h2 == state ? 1'h0 : 4'h3 == state & _T_389; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_2866 = 4'h2 == state ? _GEN_3 : _GEN_2644; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2867 = 4'h2 == state ? 128'h0 : _GEN_2645; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2868 = 4'h2 == state ? 21'h0 : _GEN_2646; // @[Cache.scala 114:16 318:18]
  wire  _GEN_2869 = 4'h2 == state ? 1'h0 : 4'h3 == state & _GEN_1005; // @[Cache.scala 116:18 318:18]
  wire  _GEN_2870 = 4'h2 == state ? pipeline_ready : _GEN_2648; // @[Cache.scala 318:18]
  wire  _GEN_2871 = 4'h2 == state ? 1'h0 : 4'h3 == state & _T_453; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_2872 = 4'h2 == state ? _GEN_3 : _GEN_2650; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2873 = 4'h2 == state ? 128'h0 : _GEN_2651; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2874 = 4'h2 == state ? 21'h0 : _GEN_2652; // @[Cache.scala 114:16 318:18]
  wire  _GEN_2875 = 4'h2 == state ? 1'h0 : 4'h3 == state & _GEN_1012; // @[Cache.scala 116:18 318:18]
  wire  _GEN_2876 = 4'h2 == state ? pipeline_ready : _GEN_2654; // @[Cache.scala 318:18]
  wire  _GEN_2877 = 4'h2 == state ? 1'h0 : 4'h3 == state & _T_517; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_2878 = 4'h2 == state ? _GEN_3 : _GEN_2656; // @[Cache.scala 318:18]
  wire [127:0] _GEN_2879 = 4'h2 == state ? 128'h0 : _GEN_2657; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_2880 = 4'h2 == state ? 21'h0 : _GEN_2658; // @[Cache.scala 114:16 318:18]
  wire  _GEN_2881 = 4'h2 == state ? 1'h0 : 4'h3 == state & _GEN_1019; // @[Cache.scala 116:18 318:18]
  wire [63:0] _GEN_3075 = 4'h2 == state ? 64'h0 : _GEN_2854; // @[Cache.scala 318:18 289:22]
  wire [3:0] _GEN_3076 = 4'h1 == state ? _GEN_985 : _GEN_2857; // @[Cache.scala 318:18]
  wire  _GEN_3079 = 4'h1 == state ? pipeline_ready : _GEN_2858; // @[Cache.scala 318:18]
  wire  _GEN_3080 = 4'h1 == state ? 1'h0 : _GEN_2859; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_3081 = 4'h1 == state ? _GEN_3 : _GEN_2860; // @[Cache.scala 318:18]
  wire [127:0] _GEN_3082 = 4'h1 == state ? 128'h0 : _GEN_2861; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_3083 = 4'h1 == state ? 21'h0 : _GEN_2862; // @[Cache.scala 114:16 318:18]
  wire  _GEN_3084 = 4'h1 == state ? 1'h0 : _GEN_2863; // @[Cache.scala 116:18 318:18]
  wire  _GEN_3085 = 4'h1 == state ? pipeline_ready : _GEN_2864; // @[Cache.scala 318:18]
  wire  _GEN_3086 = 4'h1 == state ? 1'h0 : _GEN_2865; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_3087 = 4'h1 == state ? _GEN_3 : _GEN_2866; // @[Cache.scala 318:18]
  wire [127:0] _GEN_3088 = 4'h1 == state ? 128'h0 : _GEN_2867; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_3089 = 4'h1 == state ? 21'h0 : _GEN_2868; // @[Cache.scala 114:16 318:18]
  wire  _GEN_3090 = 4'h1 == state ? 1'h0 : _GEN_2869; // @[Cache.scala 116:18 318:18]
  wire  _GEN_3091 = 4'h1 == state ? pipeline_ready : _GEN_2870; // @[Cache.scala 318:18]
  wire  _GEN_3092 = 4'h1 == state ? 1'h0 : _GEN_2871; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_3093 = 4'h1 == state ? _GEN_3 : _GEN_2872; // @[Cache.scala 318:18]
  wire [127:0] _GEN_3094 = 4'h1 == state ? 128'h0 : _GEN_2873; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_3095 = 4'h1 == state ? 21'h0 : _GEN_2874; // @[Cache.scala 114:16 318:18]
  wire  _GEN_3096 = 4'h1 == state ? 1'h0 : _GEN_2875; // @[Cache.scala 116:18 318:18]
  wire  _GEN_3097 = 4'h1 == state ? pipeline_ready : _GEN_2876; // @[Cache.scala 318:18]
  wire  _GEN_3098 = 4'h1 == state ? 1'h0 : _GEN_2877; // @[Cache.scala 108:14 318:18]
  wire [5:0] _GEN_3099 = 4'h1 == state ? _GEN_3 : _GEN_2878; // @[Cache.scala 318:18]
  wire [127:0] _GEN_3100 = 4'h1 == state ? 128'h0 : _GEN_2879; // @[Cache.scala 110:16 318:18]
  wire [20:0] _GEN_3101 = 4'h1 == state ? 21'h0 : _GEN_2880; // @[Cache.scala 114:16 318:18]
  wire  _GEN_3102 = 4'h1 == state ? 1'h0 : _GEN_2881; // @[Cache.scala 116:18 318:18]
  wire [63:0] _GEN_3296 = 4'h1 == state ? 64'h0 : _GEN_3075; // @[Cache.scala 318:18 289:22]
  wire  _GEN_3490 = 4'h0 == state ? _GEN_968 : _GEN_3079; // @[Cache.scala 318:18]
  wire [5:0] _GEN_3492 = 4'h0 == state ? _GEN_970 : _GEN_3081; // @[Cache.scala 318:18]
  wire  _GEN_3495 = 4'h0 == state ? _GEN_972 : _GEN_3085; // @[Cache.scala 318:18]
  wire [5:0] _GEN_3497 = 4'h0 == state ? _GEN_974 : _GEN_3087; // @[Cache.scala 318:18]
  wire  _GEN_3500 = 4'h0 == state ? _GEN_976 : _GEN_3091; // @[Cache.scala 318:18]
  wire [5:0] _GEN_3502 = 4'h0 == state ? _GEN_978 : _GEN_3093; // @[Cache.scala 318:18]
  wire  _GEN_3505 = 4'h0 == state ? _GEN_980 : _GEN_3097; // @[Cache.scala 318:18]
  wire [5:0] _GEN_3507 = 4'h0 == state ? _GEN_982 : _GEN_3099; // @[Cache.scala 318:18]
  reg [7:0] fi_counter; // @[Cache.scala 438:27]
  wire [1:0] fi_sram_idx = fi_counter[7:6]; // @[Cache.scala 439:31]
  wire [5:0] fi_line_idx = fi_counter[5:0]; // @[Cache.scala 440:31]
  wire  _T_608 = fi_state == 3'h2; // @[Cache.scala 443:29]
  wire  _T_609 = fi_state == 3'h1; // @[Cache.scala 443:65]
  reg  REG_13; // @[Cache.scala 443:55]
  wire  fi_update = fi_state == 3'h2 & REG_13; // @[Cache.scala 443:44]
  reg [127:0] r; // @[Reg.scala 27:20]
  wire [127:0] _GEN_3524 = 2'h1 == fi_sram_idx ? sram_out_1 : sram_out_0; // @[Reg.scala 28:{23,23}]
  wire [127:0] _GEN_3525 = 2'h2 == fi_sram_idx ? sram_out_2 : _GEN_3524; // @[Reg.scala 28:{23,23}]
  wire [127:0] _GEN_3526 = 2'h3 == fi_sram_idx ? sram_out_3 : _GEN_3525; // @[Reg.scala 28:{23,23}]
  wire [127:0] _GEN_3527 = fi_update ? _GEN_3526 : r; // @[Reg.scala 28:19 27:20 28:23]
  reg [20:0] r_1; // @[Reg.scala 27:20]
  wire [20:0] _GEN_3529 = 2'h1 == fi_sram_idx ? tag_out_1 : tag_out_0; // @[Reg.scala 28:{23,23}]
  wire [20:0] _GEN_3530 = 2'h2 == fi_sram_idx ? tag_out_2 : _GEN_3529; // @[Reg.scala 28:{23,23}]
  wire [20:0] _GEN_3531 = 2'h3 == fi_sram_idx ? tag_out_3 : _GEN_3530; // @[Reg.scala 28:{23,23}]
  wire [20:0] _GEN_3532 = fi_update ? _GEN_3531 : r_1; // @[Reg.scala 28:19 27:20 28:23]
  wire [7:0] _T_611 = fi_counter + 8'h1; // @[Cache.scala 471:38]
  wire [5:0] _GEN_3535 = _T_609 ? fi_line_idx : _GEN_3492; // @[Cache.scala 473:40 476:19]
  wire [5:0] _GEN_3537 = _T_609 ? fi_line_idx : _GEN_3497; // @[Cache.scala 473:40 476:19]
  wire [5:0] _GEN_3539 = _T_609 ? fi_line_idx : _GEN_3502; // @[Cache.scala 473:40 476:19]
  wire [5:0] _GEN_3541 = _T_609 ? fi_line_idx : _GEN_3507; // @[Cache.scala 473:40 476:19]
  wire [5:0] _GEN_3544 = fi_sram_idx == 2'h0 ? fi_line_idx : _GEN_3535; // @[Cache.scala 493:38 494:28]
  wire [5:0] _GEN_3546 = fi_sram_idx == 2'h1 ? fi_line_idx : _GEN_3537; // @[Cache.scala 493:38 494:28]
  wire  _GEN_3547 = fi_sram_idx == 2'h1 ? meta_1_io_valid_r_async & meta_1_io_dirty_r_async : fi_sram_idx == 2'h0 & (
    meta_0_io_valid_r_async & meta_0_io_dirty_r_async); // @[Cache.scala 493:38 495:22]
  wire [5:0] _GEN_3548 = fi_sram_idx == 2'h2 ? fi_line_idx : _GEN_3539; // @[Cache.scala 493:38 494:28]
  wire  _GEN_3549 = fi_sram_idx == 2'h2 ? meta_2_io_valid_r_async & meta_2_io_dirty_r_async : _GEN_3547; // @[Cache.scala 493:38 495:22]
  wire [5:0] _GEN_3550 = fi_sram_idx == 2'h3 ? fi_line_idx : _GEN_3541; // @[Cache.scala 493:38 494:28]
  wire  _GEN_3551 = fi_sram_idx == 2'h3 ? meta_3_io_valid_r_async & meta_3_io_dirty_r_async : _GEN_3549; // @[Cache.scala 493:38 495:22]
  wire  _T_623 = _T_611 == 8'h0; // @[Cache.scala 502:33]
  wire [2:0] _GEN_3552 = _T_611 == 8'h0 ? 3'h5 : fi_state; // @[Cache.scala 502:42 503:22 435:25]
  wire [2:0] _GEN_3555 = _T_320 ? 3'h3 : fi_state; // @[Cache.scala 508:31 509:20 435:25]
  wire [2:0] _GEN_3556 = _T_320 ? 3'h4 : fi_state; // @[Cache.scala 513:31 514:20 435:25]
  wire [2:0] _GEN_3557 = _T_623 ? 3'h5 : 3'h1; // @[Cache.scala 520:42 521:22 523:22]
  wire [7:0] _GEN_3558 = _T_322 ? _T_611 : fi_counter; // @[Cache.scala 518:32 519:22 438:27]
  wire [2:0] _GEN_3559 = _T_322 ? _GEN_3557 : fi_state; // @[Cache.scala 435:25 518:32]
  wire [2:0] _GEN_3561 = 3'h5 == fi_state ? 3'h0 : fi_state; // @[Cache.scala 483:23 529:18 435:25]
  wire [7:0] _GEN_3562 = 3'h4 == fi_state ? _GEN_3558 : fi_counter; // @[Cache.scala 483:23 438:27]
  wire [2:0] _GEN_3563 = 3'h4 == fi_state ? _GEN_3559 : _GEN_3561; // @[Cache.scala 483:23]
  wire [2:0] _GEN_3565 = 3'h3 == fi_state ? _GEN_3556 : _GEN_3563; // @[Cache.scala 483:23]
  wire [7:0] _GEN_3566 = 3'h3 == fi_state ? fi_counter : _GEN_3562; // @[Cache.scala 483:23 438:27]
  wire [5:0] _GEN_3571 = 3'h1 == fi_state ? _GEN_3544 : _GEN_3535; // @[Cache.scala 483:23]
  wire [5:0] _GEN_3572 = 3'h1 == fi_state ? _GEN_3546 : _GEN_3537; // @[Cache.scala 483:23]
  wire [5:0] _GEN_3573 = 3'h1 == fi_state ? _GEN_3548 : _GEN_3539; // @[Cache.scala 483:23]
  wire [5:0] _GEN_3574 = 3'h1 == fi_state ? _GEN_3550 : _GEN_3541; // @[Cache.scala 483:23]
  wire  _T_632 = state == 4'h1; // @[Cache.scala 540:27]
  wire  _T_633 = state == 4'h4; // @[Cache.scala 541:27]
  wire  _T_634 = state == 4'h1 | _T_633; // @[Cache.scala 540:45]
  wire  _T_635 = state == 4'h5; // @[Cache.scala 542:27]
  wire  _T_636 = _T_634 | _T_635; // @[Cache.scala 541:46]
  wire  _T_638 = _T_636 | _T_608; // @[Cache.scala 542:46]
  wire  _T_639 = fi_state == 3'h3; // @[Cache.scala 544:30]
  wire [31:0] _T_644 = {s2_addr[31:4],4'h0}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3585 = _T_632 ? _T_644 : 32'h0; // @[Cache.scala 546:21 547:33 548:23]
  wire [31:0] _T_647 = {1'h1,s2_reg_tag_r,s2_idx,4'h0}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_3586 = _T_633 ? _T_647 : _GEN_3585; // @[Cache.scala 550:34 553:23]
  wire [31:0] _T_650 = {1'h1,_GEN_3532,fi_line_idx,4'h0}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_3588 = _T_633 ? s2_reg_dat_w[63:0] : 64'h0; // @[Cache.scala 561:22 562:34 563:24]
  wire [63:0] _GEN_3589 = _T_635 ? s2_reg_dat_w[127:64] : _GEN_3588; // @[Cache.scala 565:34 566:24]
  wire [63:0] _GEN_3590 = _T_608 ? _GEN_3527[63:0] : _GEN_3589; // @[Cache.scala 568:33 569:24]
  wire  _T_669 = _T_633 | _T_635; // @[Cache.scala 577:49]
  wire  _T_671 = _T_669 | _T_608; // @[Cache.scala 578:49]
  wire  _T_675 = state == 4'h6; // @[Cache.scala 584:28]
  wire  _T_676 = state == 4'h2 | _T_675; // @[Cache.scala 583:47]
  wire  _T_677 = fi_state == 3'h4; // @[Cache.scala 585:31]
  ysyx_210128_Sram sram_0 ( // @[Cache.scala 89:22]
    .clock(sram_0_clock),
    .io_en(sram_0_io_en),
    .io_wen(sram_0_io_wen),
    .io_addr(sram_0_io_addr),
    .io_wdata(sram_0_io_wdata),
    .io_rdata(sram_0_io_rdata)
  );
  ysyx_210128_Sram sram_1 ( // @[Cache.scala 89:22]
    .clock(sram_1_clock),
    .io_en(sram_1_io_en),
    .io_wen(sram_1_io_wen),
    .io_addr(sram_1_io_addr),
    .io_wdata(sram_1_io_wdata),
    .io_rdata(sram_1_io_rdata)
  );
  ysyx_210128_Sram sram_2 ( // @[Cache.scala 89:22]
    .clock(sram_2_clock),
    .io_en(sram_2_io_en),
    .io_wen(sram_2_io_wen),
    .io_addr(sram_2_io_addr),
    .io_wdata(sram_2_io_wdata),
    .io_rdata(sram_2_io_rdata)
  );
  ysyx_210128_Sram sram_3 ( // @[Cache.scala 89:22]
    .clock(sram_3_clock),
    .io_en(sram_3_io_en),
    .io_wen(sram_3_io_wen),
    .io_addr(sram_3_io_addr),
    .io_wdata(sram_3_io_wdata),
    .io_rdata(sram_3_io_rdata)
  );
  ysyx_210128_Meta meta_0 ( // @[Cache.scala 97:22]
    .clock(meta_0_clock),
    .reset(meta_0_reset),
    .io_idx(meta_0_io_idx),
    .io_tag_r(meta_0_io_tag_r),
    .io_tag_w(meta_0_io_tag_w),
    .io_tag_wen(meta_0_io_tag_wen),
    .io_dirty_r_async(meta_0_io_dirty_r_async),
    .io_dirty_w(meta_0_io_dirty_w),
    .io_dirty_wen(meta_0_io_dirty_wen),
    .io_valid_r_async(meta_0_io_valid_r_async),
    .io_invalidate(meta_0_io_invalidate)
  );
  ysyx_210128_Meta meta_1 ( // @[Cache.scala 97:22]
    .clock(meta_1_clock),
    .reset(meta_1_reset),
    .io_idx(meta_1_io_idx),
    .io_tag_r(meta_1_io_tag_r),
    .io_tag_w(meta_1_io_tag_w),
    .io_tag_wen(meta_1_io_tag_wen),
    .io_dirty_r_async(meta_1_io_dirty_r_async),
    .io_dirty_w(meta_1_io_dirty_w),
    .io_dirty_wen(meta_1_io_dirty_wen),
    .io_valid_r_async(meta_1_io_valid_r_async),
    .io_invalidate(meta_1_io_invalidate)
  );
  ysyx_210128_Meta meta_2 ( // @[Cache.scala 97:22]
    .clock(meta_2_clock),
    .reset(meta_2_reset),
    .io_idx(meta_2_io_idx),
    .io_tag_r(meta_2_io_tag_r),
    .io_tag_w(meta_2_io_tag_w),
    .io_tag_wen(meta_2_io_tag_wen),
    .io_dirty_r_async(meta_2_io_dirty_r_async),
    .io_dirty_w(meta_2_io_dirty_w),
    .io_dirty_wen(meta_2_io_dirty_wen),
    .io_valid_r_async(meta_2_io_valid_r_async),
    .io_invalidate(meta_2_io_invalidate)
  );
  ysyx_210128_Meta meta_3 ( // @[Cache.scala 97:22]
    .clock(meta_3_clock),
    .reset(meta_3_reset),
    .io_idx(meta_3_io_idx),
    .io_tag_r(meta_3_io_tag_r),
    .io_tag_w(meta_3_io_tag_w),
    .io_tag_wen(meta_3_io_tag_wen),
    .io_dirty_r_async(meta_3_io_dirty_r_async),
    .io_dirty_w(meta_3_io_dirty_w),
    .io_dirty_wen(meta_3_io_dirty_wen),
    .io_valid_r_async(meta_3_io_valid_r_async),
    .io_invalidate(meta_3_io_invalidate)
  );
  assign io_in_req_ready = pipeline_ready & ~fi_valid; // @[Cache.scala 287:34]
  assign io_in_resp_valid = s2_hit_real & ~s2_wen & state != 4'h8 | _T_18; // @[Cache.scala 288:71]
  assign io_in_resp_bits_id = s2_id; // @[Cache.scala 294:19]
  assign io_in_resp_bits_rdata = 4'h0 == state ? _GEN_229 : _GEN_3296; // @[Cache.scala 318:18]
  assign io_out_req_valid = _T_638 | _T_639; // @[Cache.scala 543:45]
  assign io_out_req_bits_addr = _T_608 ? _T_650 : _GEN_3586; // @[Cache.scala 555:33 556:23]
  assign io_out_req_bits_aen = _T_634 | _T_608; // @[Cache.scala 559:49]
  assign io_out_req_bits_wdata = _T_639 ? _GEN_3527[127:64] : _GEN_3590; // @[Cache.scala 571:33 572:24]
  assign io_out_req_bits_wlast = _T_635 | _T_639; // @[Cache.scala 575:51]
  assign io_out_req_bits_wen = _T_671 | _T_639; // @[Cache.scala 579:48]
  assign io_out_resp_ready = _T_676 | _T_677; // @[Cache.scala 584:47]
  assign _WIRE_10_0 = 3'h0 == fi_state ? 1'h0 : _GEN_3577; // @[Cache.scala 483:23]
  assign sram_0_clock = clock;
  assign sram_0_io_en = _T_609 | _GEN_3490; // @[Cache.scala 473:40 475:17]
  assign sram_0_io_wen = 4'h0 == state ? _GEN_969 : _GEN_3080; // @[Cache.scala 318:18]
  assign sram_0_io_addr = _T_609 ? fi_line_idx : _GEN_3492; // @[Cache.scala 473:40 476:19]
  assign sram_0_io_wdata = 4'h0 == state ? _GEN_971 : _GEN_3082; // @[Cache.scala 318:18]
  assign sram_1_clock = clock;
  assign sram_1_io_en = _T_609 | _GEN_3495; // @[Cache.scala 473:40 475:17]
  assign sram_1_io_wen = 4'h0 == state ? _GEN_973 : _GEN_3086; // @[Cache.scala 318:18]
  assign sram_1_io_addr = _T_609 ? fi_line_idx : _GEN_3497; // @[Cache.scala 473:40 476:19]
  assign sram_1_io_wdata = 4'h0 == state ? _GEN_975 : _GEN_3088; // @[Cache.scala 318:18]
  assign sram_2_clock = clock;
  assign sram_2_io_en = _T_609 | _GEN_3500; // @[Cache.scala 473:40 475:17]
  assign sram_2_io_wen = 4'h0 == state ? _GEN_977 : _GEN_3092; // @[Cache.scala 318:18]
  assign sram_2_io_addr = _T_609 ? fi_line_idx : _GEN_3502; // @[Cache.scala 473:40 476:19]
  assign sram_2_io_wdata = 4'h0 == state ? _GEN_979 : _GEN_3094; // @[Cache.scala 318:18]
  assign sram_3_clock = clock;
  assign sram_3_io_en = _T_609 | _GEN_3505; // @[Cache.scala 473:40 475:17]
  assign sram_3_io_wen = 4'h0 == state ? _GEN_981 : _GEN_3098; // @[Cache.scala 318:18]
  assign sram_3_io_addr = _T_609 ? fi_line_idx : _GEN_3507; // @[Cache.scala 473:40 476:19]
  assign sram_3_io_wdata = 4'h0 == state ? _GEN_983 : _GEN_3100; // @[Cache.scala 318:18]
  assign meta_0_clock = clock;
  assign meta_0_reset = reset;
  assign meta_0_io_idx = 3'h0 == fi_state ? _GEN_3535 : _GEN_3571; // @[Cache.scala 483:23]
  assign meta_0_io_tag_w = 4'h0 == state ? 21'h0 : _GEN_3083; // @[Cache.scala 114:16 318:18]
  assign meta_0_io_tag_wen = 4'h0 == state ? 1'h0 : _GEN_3080; // @[Cache.scala 115:18 318:18]
  assign meta_0_io_dirty_w = 4'h0 == state ? _GEN_969 : _GEN_3084; // @[Cache.scala 318:18]
  assign meta_0_io_dirty_wen = 4'h0 == state ? _GEN_969 : _GEN_3080; // @[Cache.scala 318:18]
  assign meta_0_io_invalidate = 3'h0 == fi_state ? 1'h0 : _GEN_3577; // @[Cache.scala 483:23]
  assign meta_1_clock = clock;
  assign meta_1_reset = reset;
  assign meta_1_io_idx = 3'h0 == fi_state ? _GEN_3537 : _GEN_3572; // @[Cache.scala 483:23]
  assign meta_1_io_tag_w = 4'h0 == state ? 21'h0 : _GEN_3089; // @[Cache.scala 114:16 318:18]
  assign meta_1_io_tag_wen = 4'h0 == state ? 1'h0 : _GEN_3086; // @[Cache.scala 115:18 318:18]
  assign meta_1_io_dirty_w = 4'h0 == state ? _GEN_973 : _GEN_3090; // @[Cache.scala 318:18]
  assign meta_1_io_dirty_wen = 4'h0 == state ? _GEN_973 : _GEN_3086; // @[Cache.scala 318:18]
  assign meta_1_io_invalidate = 3'h0 == fi_state ? 1'h0 : _GEN_3577; // @[Cache.scala 483:23]
  assign meta_2_clock = clock;
  assign meta_2_reset = reset;
  assign meta_2_io_idx = 3'h0 == fi_state ? _GEN_3539 : _GEN_3573; // @[Cache.scala 483:23]
  assign meta_2_io_tag_w = 4'h0 == state ? 21'h0 : _GEN_3095; // @[Cache.scala 114:16 318:18]
  assign meta_2_io_tag_wen = 4'h0 == state ? 1'h0 : _GEN_3092; // @[Cache.scala 115:18 318:18]
  assign meta_2_io_dirty_w = 4'h0 == state ? _GEN_977 : _GEN_3096; // @[Cache.scala 318:18]
  assign meta_2_io_dirty_wen = 4'h0 == state ? _GEN_977 : _GEN_3092; // @[Cache.scala 318:18]
  assign meta_2_io_invalidate = 3'h0 == fi_state ? 1'h0 : _GEN_3577; // @[Cache.scala 483:23]
  assign meta_3_clock = clock;
  assign meta_3_reset = reset;
  assign meta_3_io_idx = 3'h0 == fi_state ? _GEN_3541 : _GEN_3574; // @[Cache.scala 483:23]
  assign meta_3_io_tag_w = 4'h0 == state ? 21'h0 : _GEN_3101; // @[Cache.scala 114:16 318:18]
  assign meta_3_io_tag_wen = 4'h0 == state ? 1'h0 : _GEN_3098; // @[Cache.scala 115:18 318:18]
  assign meta_3_io_dirty_w = 4'h0 == state ? _GEN_981 : _GEN_3102; // @[Cache.scala 318:18]
  assign meta_3_io_dirty_wen = 4'h0 == state ? _GEN_981 : _GEN_3098; // @[Cache.scala 318:18]
  assign meta_3_io_invalidate = 3'h0 == fi_state ? 1'h0 : _GEN_3577; // @[Cache.scala 483:23]
  always @(posedge clock) begin
    REG <= meta_0_io_valid_r_async; // @[Cache.scala 123:59]
    REG_1 <= meta_1_io_valid_r_async; // @[Cache.scala 123:59]
    REG_2 <= meta_2_io_valid_r_async; // @[Cache.scala 123:59]
    REG_3 <= meta_3_io_valid_r_async; // @[Cache.scala 123:59]
    REG_4 <= meta_0_io_dirty_r_async; // @[Cache.scala 124:59]
    REG_5 <= meta_1_io_dirty_r_async; // @[Cache.scala 124:59]
    REG_6 <= meta_2_io_dirty_r_async; // @[Cache.scala 124:59]
    REG_7 <= meta_3_io_dirty_r_async; // @[Cache.scala 124:59]
    if (reset) begin // @[Cache.scala 129:22]
      plru0_0 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_0 <= _GEN_230;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_0 <= _GEN_2661;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_1 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_1 <= _GEN_231;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_1 <= _GEN_2662;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_2 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_2 <= _GEN_232;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_2 <= _GEN_2663;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_3 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_3 <= _GEN_233;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_3 <= _GEN_2664;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_4 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_4 <= _GEN_234;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_4 <= _GEN_2665;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_5 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_5 <= _GEN_235;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_5 <= _GEN_2666;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_6 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_6 <= _GEN_236;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_6 <= _GEN_2667;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_7 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_7 <= _GEN_237;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_7 <= _GEN_2668;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_8 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_8 <= _GEN_238;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_8 <= _GEN_2669;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_9 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_9 <= _GEN_239;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_9 <= _GEN_2670;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_10 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_10 <= _GEN_240;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_10 <= _GEN_2671;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_11 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_11 <= _GEN_241;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_11 <= _GEN_2672;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_12 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_12 <= _GEN_242;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_12 <= _GEN_2673;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_13 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_13 <= _GEN_243;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_13 <= _GEN_2674;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_14 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_14 <= _GEN_244;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_14 <= _GEN_2675;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_15 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_15 <= _GEN_245;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_15 <= _GEN_2676;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_16 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_16 <= _GEN_246;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_16 <= _GEN_2677;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_17 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_17 <= _GEN_247;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_17 <= _GEN_2678;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_18 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_18 <= _GEN_248;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_18 <= _GEN_2679;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_19 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_19 <= _GEN_249;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_19 <= _GEN_2680;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_20 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_20 <= _GEN_250;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_20 <= _GEN_2681;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_21 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_21 <= _GEN_251;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_21 <= _GEN_2682;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_22 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_22 <= _GEN_252;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_22 <= _GEN_2683;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_23 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_23 <= _GEN_253;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_23 <= _GEN_2684;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_24 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_24 <= _GEN_254;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_24 <= _GEN_2685;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_25 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_25 <= _GEN_255;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_25 <= _GEN_2686;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_26 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_26 <= _GEN_256;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_26 <= _GEN_2687;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_27 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_27 <= _GEN_257;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_27 <= _GEN_2688;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_28 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_28 <= _GEN_258;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_28 <= _GEN_2689;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_29 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_29 <= _GEN_259;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_29 <= _GEN_2690;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_30 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_30 <= _GEN_260;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_30 <= _GEN_2691;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_31 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_31 <= _GEN_261;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_31 <= _GEN_2692;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_32 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_32 <= _GEN_262;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_32 <= _GEN_2693;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_33 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_33 <= _GEN_263;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_33 <= _GEN_2694;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_34 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_34 <= _GEN_264;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_34 <= _GEN_2695;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_35 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_35 <= _GEN_265;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_35 <= _GEN_2696;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_36 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_36 <= _GEN_266;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_36 <= _GEN_2697;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_37 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_37 <= _GEN_267;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_37 <= _GEN_2698;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_38 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_38 <= _GEN_268;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_38 <= _GEN_2699;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_39 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_39 <= _GEN_269;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_39 <= _GEN_2700;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_40 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_40 <= _GEN_270;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_40 <= _GEN_2701;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_41 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_41 <= _GEN_271;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_41 <= _GEN_2702;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_42 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_42 <= _GEN_272;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_42 <= _GEN_2703;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_43 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_43 <= _GEN_273;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_43 <= _GEN_2704;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_44 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_44 <= _GEN_274;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_44 <= _GEN_2705;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_45 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_45 <= _GEN_275;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_45 <= _GEN_2706;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_46 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_46 <= _GEN_276;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_46 <= _GEN_2707;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_47 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_47 <= _GEN_277;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_47 <= _GEN_2708;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_48 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_48 <= _GEN_278;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_48 <= _GEN_2709;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_49 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_49 <= _GEN_279;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_49 <= _GEN_2710;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_50 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_50 <= _GEN_280;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_50 <= _GEN_2711;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_51 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_51 <= _GEN_281;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_51 <= _GEN_2712;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_52 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_52 <= _GEN_282;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_52 <= _GEN_2713;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_53 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_53 <= _GEN_283;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_53 <= _GEN_2714;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_54 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_54 <= _GEN_284;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_54 <= _GEN_2715;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_55 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_55 <= _GEN_285;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_55 <= _GEN_2716;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_56 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_56 <= _GEN_286;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_56 <= _GEN_2717;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_57 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_57 <= _GEN_287;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_57 <= _GEN_2718;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_58 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_58 <= _GEN_288;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_58 <= _GEN_2719;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_59 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_59 <= _GEN_289;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_59 <= _GEN_2720;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_60 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_60 <= _GEN_290;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_60 <= _GEN_2721;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_61 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_61 <= _GEN_291;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_61 <= _GEN_2722;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_62 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_62 <= _GEN_292;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_62 <= _GEN_2723;
      end
    end
    if (reset) begin // @[Cache.scala 129:22]
      plru0_63 <= 1'h0; // @[Cache.scala 129:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru0_63 <= _GEN_293;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru0_63 <= _GEN_2724;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_0 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_0 <= _GEN_422;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_0 <= _GEN_2725;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_1 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_1 <= _GEN_423;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_1 <= _GEN_2726;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_2 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_2 <= _GEN_424;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_2 <= _GEN_2727;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_3 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_3 <= _GEN_425;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_3 <= _GEN_2728;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_4 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_4 <= _GEN_426;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_4 <= _GEN_2729;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_5 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_5 <= _GEN_427;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_5 <= _GEN_2730;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_6 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_6 <= _GEN_428;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_6 <= _GEN_2731;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_7 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_7 <= _GEN_429;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_7 <= _GEN_2732;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_8 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_8 <= _GEN_430;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_8 <= _GEN_2733;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_9 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_9 <= _GEN_431;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_9 <= _GEN_2734;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_10 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_10 <= _GEN_432;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_10 <= _GEN_2735;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_11 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_11 <= _GEN_433;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_11 <= _GEN_2736;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_12 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_12 <= _GEN_434;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_12 <= _GEN_2737;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_13 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_13 <= _GEN_435;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_13 <= _GEN_2738;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_14 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_14 <= _GEN_436;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_14 <= _GEN_2739;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_15 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_15 <= _GEN_437;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_15 <= _GEN_2740;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_16 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_16 <= _GEN_438;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_16 <= _GEN_2741;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_17 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_17 <= _GEN_439;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_17 <= _GEN_2742;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_18 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_18 <= _GEN_440;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_18 <= _GEN_2743;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_19 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_19 <= _GEN_441;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_19 <= _GEN_2744;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_20 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_20 <= _GEN_442;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_20 <= _GEN_2745;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_21 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_21 <= _GEN_443;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_21 <= _GEN_2746;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_22 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_22 <= _GEN_444;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_22 <= _GEN_2747;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_23 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_23 <= _GEN_445;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_23 <= _GEN_2748;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_24 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_24 <= _GEN_446;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_24 <= _GEN_2749;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_25 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_25 <= _GEN_447;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_25 <= _GEN_2750;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_26 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_26 <= _GEN_448;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_26 <= _GEN_2751;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_27 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_27 <= _GEN_449;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_27 <= _GEN_2752;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_28 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_28 <= _GEN_450;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_28 <= _GEN_2753;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_29 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_29 <= _GEN_451;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_29 <= _GEN_2754;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_30 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_30 <= _GEN_452;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_30 <= _GEN_2755;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_31 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_31 <= _GEN_453;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_31 <= _GEN_2756;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_32 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_32 <= _GEN_454;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_32 <= _GEN_2757;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_33 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_33 <= _GEN_455;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_33 <= _GEN_2758;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_34 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_34 <= _GEN_456;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_34 <= _GEN_2759;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_35 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_35 <= _GEN_457;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_35 <= _GEN_2760;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_36 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_36 <= _GEN_458;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_36 <= _GEN_2761;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_37 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_37 <= _GEN_459;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_37 <= _GEN_2762;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_38 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_38 <= _GEN_460;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_38 <= _GEN_2763;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_39 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_39 <= _GEN_461;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_39 <= _GEN_2764;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_40 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_40 <= _GEN_462;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_40 <= _GEN_2765;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_41 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_41 <= _GEN_463;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_41 <= _GEN_2766;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_42 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_42 <= _GEN_464;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_42 <= _GEN_2767;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_43 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_43 <= _GEN_465;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_43 <= _GEN_2768;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_44 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_44 <= _GEN_466;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_44 <= _GEN_2769;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_45 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_45 <= _GEN_467;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_45 <= _GEN_2770;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_46 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_46 <= _GEN_468;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_46 <= _GEN_2771;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_47 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_47 <= _GEN_469;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_47 <= _GEN_2772;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_48 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_48 <= _GEN_470;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_48 <= _GEN_2773;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_49 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_49 <= _GEN_471;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_49 <= _GEN_2774;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_50 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_50 <= _GEN_472;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_50 <= _GEN_2775;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_51 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_51 <= _GEN_473;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_51 <= _GEN_2776;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_52 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_52 <= _GEN_474;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_52 <= _GEN_2777;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_53 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_53 <= _GEN_475;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_53 <= _GEN_2778;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_54 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_54 <= _GEN_476;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_54 <= _GEN_2779;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_55 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_55 <= _GEN_477;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_55 <= _GEN_2780;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_56 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_56 <= _GEN_478;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_56 <= _GEN_2781;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_57 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_57 <= _GEN_479;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_57 <= _GEN_2782;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_58 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_58 <= _GEN_480;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_58 <= _GEN_2783;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_59 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_59 <= _GEN_481;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_59 <= _GEN_2784;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_60 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_60 <= _GEN_482;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_60 <= _GEN_2785;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_61 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_61 <= _GEN_483;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_61 <= _GEN_2786;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_62 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_62 <= _GEN_484;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_62 <= _GEN_2787;
      end
    end
    if (reset) begin // @[Cache.scala 131:22]
      plru1_63 <= 1'h0; // @[Cache.scala 131:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru1_63 <= _GEN_485;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru1_63 <= _GEN_2788;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_0 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_0 <= _GEN_486;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_0 <= _GEN_2789;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_1 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_1 <= _GEN_487;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_1 <= _GEN_2790;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_2 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_2 <= _GEN_488;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_2 <= _GEN_2791;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_3 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_3 <= _GEN_489;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_3 <= _GEN_2792;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_4 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_4 <= _GEN_490;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_4 <= _GEN_2793;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_5 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_5 <= _GEN_491;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_5 <= _GEN_2794;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_6 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_6 <= _GEN_492;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_6 <= _GEN_2795;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_7 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_7 <= _GEN_493;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_7 <= _GEN_2796;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_8 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_8 <= _GEN_494;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_8 <= _GEN_2797;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_9 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_9 <= _GEN_495;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_9 <= _GEN_2798;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_10 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_10 <= _GEN_496;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_10 <= _GEN_2799;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_11 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_11 <= _GEN_497;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_11 <= _GEN_2800;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_12 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_12 <= _GEN_498;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_12 <= _GEN_2801;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_13 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_13 <= _GEN_499;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_13 <= _GEN_2802;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_14 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_14 <= _GEN_500;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_14 <= _GEN_2803;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_15 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_15 <= _GEN_501;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_15 <= _GEN_2804;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_16 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_16 <= _GEN_502;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_16 <= _GEN_2805;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_17 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_17 <= _GEN_503;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_17 <= _GEN_2806;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_18 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_18 <= _GEN_504;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_18 <= _GEN_2807;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_19 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_19 <= _GEN_505;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_19 <= _GEN_2808;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_20 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_20 <= _GEN_506;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_20 <= _GEN_2809;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_21 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_21 <= _GEN_507;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_21 <= _GEN_2810;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_22 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_22 <= _GEN_508;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_22 <= _GEN_2811;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_23 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_23 <= _GEN_509;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_23 <= _GEN_2812;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_24 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_24 <= _GEN_510;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_24 <= _GEN_2813;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_25 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_25 <= _GEN_511;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_25 <= _GEN_2814;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_26 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_26 <= _GEN_512;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_26 <= _GEN_2815;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_27 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_27 <= _GEN_513;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_27 <= _GEN_2816;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_28 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_28 <= _GEN_514;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_28 <= _GEN_2817;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_29 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_29 <= _GEN_515;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_29 <= _GEN_2818;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_30 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_30 <= _GEN_516;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_30 <= _GEN_2819;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_31 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_31 <= _GEN_517;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_31 <= _GEN_2820;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_32 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_32 <= _GEN_518;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_32 <= _GEN_2821;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_33 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_33 <= _GEN_519;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_33 <= _GEN_2822;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_34 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_34 <= _GEN_520;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_34 <= _GEN_2823;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_35 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_35 <= _GEN_521;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_35 <= _GEN_2824;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_36 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_36 <= _GEN_522;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_36 <= _GEN_2825;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_37 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_37 <= _GEN_523;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_37 <= _GEN_2826;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_38 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_38 <= _GEN_524;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_38 <= _GEN_2827;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_39 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_39 <= _GEN_525;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_39 <= _GEN_2828;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_40 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_40 <= _GEN_526;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_40 <= _GEN_2829;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_41 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_41 <= _GEN_527;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_41 <= _GEN_2830;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_42 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_42 <= _GEN_528;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_42 <= _GEN_2831;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_43 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_43 <= _GEN_529;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_43 <= _GEN_2832;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_44 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_44 <= _GEN_530;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_44 <= _GEN_2833;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_45 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_45 <= _GEN_531;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_45 <= _GEN_2834;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_46 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_46 <= _GEN_532;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_46 <= _GEN_2835;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_47 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_47 <= _GEN_533;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_47 <= _GEN_2836;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_48 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_48 <= _GEN_534;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_48 <= _GEN_2837;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_49 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_49 <= _GEN_535;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_49 <= _GEN_2838;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_50 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_50 <= _GEN_536;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_50 <= _GEN_2839;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_51 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_51 <= _GEN_537;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_51 <= _GEN_2840;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_52 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_52 <= _GEN_538;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_52 <= _GEN_2841;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_53 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_53 <= _GEN_539;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_53 <= _GEN_2842;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_54 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_54 <= _GEN_540;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_54 <= _GEN_2843;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_55 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_55 <= _GEN_541;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_55 <= _GEN_2844;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_56 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_56 <= _GEN_542;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_56 <= _GEN_2845;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_57 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_57 <= _GEN_543;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_57 <= _GEN_2846;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_58 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_58 <= _GEN_544;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_58 <= _GEN_2847;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_59 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_59 <= _GEN_545;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_59 <= _GEN_2848;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_60 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_60 <= _GEN_546;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_60 <= _GEN_2849;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_61 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_61 <= _GEN_547;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_61 <= _GEN_2850;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_62 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_62 <= _GEN_548;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_62 <= _GEN_2851;
      end
    end
    if (reset) begin // @[Cache.scala 133:22]
      plru2_63 <= 1'h0; // @[Cache.scala 133:22]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      if (REG_11) begin // @[Cache.scala 325:37]
        if (s2_hit) begin // @[Cache.scala 326:23]
          plru2_63 <= _GEN_549;
        end
      end
    end else if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h2 == state)) begin // @[Cache.scala 318:18]
        plru2_63 <= _GEN_2852;
      end
    end
    REG_9 <= (hit_ready | _T_18) & io_in_resp_ready | invalid_ready; // @[Cache.scala 282:66]
    if (reset) begin // @[Cache.scala 215:25]
      s2_addr <= 32'h0; // @[Cache.scala 215:25]
    end else if (pipeline_ready) begin // @[Cache.scala 246:24]
      s2_addr <= io_in_req_bits_addr; // @[Cache.scala 248:14]
    end
    if (reset) begin // @[Cache.scala 239:27]
      s2_reg_hit <= 1'h0; // @[Cache.scala 239:27]
    end else if (!(pipeline_ready)) begin // @[Cache.scala 246:24]
      if (~pipeline_ready & REG_8) begin // @[Cache.scala 256:58]
        s2_reg_hit <= s2_hit; // @[Cache.scala 259:18]
      end
    end
    if (reset) begin // @[Cache.scala 219:25]
      s2_wen <= 1'h0; // @[Cache.scala 219:25]
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      s2_wen <= _GEN_27;
    end else if (4'h1 == state) begin // @[Cache.scala 318:18]
      s2_wen <= _GEN_27;
    end else if (4'h2 == state) begin // @[Cache.scala 318:18]
      s2_wen <= _GEN_27;
    end else begin
      s2_wen <= _GEN_2853;
    end
    if (reset) begin // @[Cache.scala 213:22]
      state <= 4'h8; // @[Cache.scala 213:22]
    end else if (fi_fire) begin // @[Cache.scala 447:18]
      state <= 4'h8; // @[Cache.scala 448:11]
    end else if (pipeline_ready) begin // @[Cache.scala 417:24]
      if (io_in_req_valid) begin // @[Cache.scala 418:17]
        state <= 4'h0;
      end else begin
        state <= 4'h8;
      end
    end else if (4'h0 == state) begin // @[Cache.scala 318:18]
      state <= _GEN_984;
    end else begin
      state <= _GEN_3076;
    end
    if (reset) begin // @[Utils.scala 34:20]
      fi_valid <= 1'h0; // @[Utils.scala 34:20]
    end else if (fi_finish) begin // @[Utils.scala 41:19]
      fi_valid <= 1'h0; // @[Utils.scala 41:23]
    end else begin
      fi_valid <= _GEN_0;
    end
    if (reset) begin // @[Cache.scala 435:25]
      fi_state <= 3'h0; // @[Cache.scala 435:25]
    end else if (3'h0 == fi_state) begin // @[Cache.scala 483:23]
      if (fi_fire) begin // @[Cache.scala 485:24]
        fi_state <= 3'h1; // @[Cache.scala 487:20]
      end
    end else if (3'h1 == fi_state) begin // @[Cache.scala 483:23]
      if (_GEN_3551) begin // @[Cache.scala 498:25]
        fi_state <= 3'h2; // @[Cache.scala 499:20]
      end else begin
        fi_state <= _GEN_3552;
      end
    end else if (3'h2 == fi_state) begin // @[Cache.scala 483:23]
      fi_state <= _GEN_3555;
    end else begin
      fi_state <= _GEN_3565;
    end
    if (reset) begin // @[Cache.scala 220:25]
      s2_wdata <= 64'h0; // @[Cache.scala 220:25]
    end else if (pipeline_ready) begin // @[Cache.scala 246:24]
      s2_wdata <= io_in_req_bits_wdata; // @[Cache.scala 250:14]
    end
    if (reset) begin // @[Cache.scala 221:25]
      s2_wmask <= 8'h0; // @[Cache.scala 221:25]
    end else if (pipeline_ready) begin // @[Cache.scala 246:24]
      s2_wmask <= io_in_req_bits_wmask; // @[Cache.scala 251:14]
    end
    if (reset) begin // @[Cache.scala 223:25]
      s2_id <= 4'h0; // @[Cache.scala 223:25]
    end else if (pipeline_ready) begin // @[Cache.scala 246:24]
      s2_id <= io_in_req_bits_id; // @[Cache.scala 255:14]
    end
    if (reset) begin // @[Cache.scala 241:29]
      s2_reg_rdata <= 128'h0; // @[Cache.scala 241:29]
    end else if (!(pipeline_ready)) begin // @[Cache.scala 246:24]
      if (~pipeline_ready & REG_8) begin // @[Cache.scala 256:58]
        if (2'h3 == s2_way) begin // @[Cache.scala 261:18]
          s2_reg_rdata <= sram_out_3; // @[Cache.scala 261:18]
        end else begin
          s2_reg_rdata <= _GEN_6;
        end
      end
    end
    if (reset) begin // @[Cache.scala 242:29]
      s2_reg_dirty <= 1'h0; // @[Cache.scala 242:29]
    end else if (!(pipeline_ready)) begin // @[Cache.scala 246:24]
      if (~pipeline_ready & REG_8) begin // @[Cache.scala 256:58]
        if (2'h3 == replace_way) begin // @[Cache.scala 262:18]
          s2_reg_dirty <= REG_7; // @[Cache.scala 262:18]
        end else begin
          s2_reg_dirty <= _GEN_10;
        end
      end
    end
    if (reset) begin // @[Cache.scala 243:29]
      s2_reg_tag_r <= 21'h0; // @[Cache.scala 243:29]
    end else if (!(pipeline_ready)) begin // @[Cache.scala 246:24]
      if (~pipeline_ready & REG_8) begin // @[Cache.scala 256:58]
        if (2'h3 == replace_way) begin // @[Cache.scala 263:18]
          s2_reg_tag_r <= tag_out_3; // @[Cache.scala 263:18]
        end else begin
          s2_reg_tag_r <= _GEN_14;
        end
      end
    end
    if (reset) begin // @[Cache.scala 244:29]
      s2_reg_dat_w <= 128'h0; // @[Cache.scala 244:29]
    end else if (!(pipeline_ready)) begin // @[Cache.scala 246:24]
      if (~pipeline_ready & REG_8) begin // @[Cache.scala 256:58]
        if (2'h3 == replace_way) begin // @[Cache.scala 264:18]
          s2_reg_dat_w <= sram_out_3; // @[Cache.scala 264:18]
        end else begin
          s2_reg_dat_w <= _GEN_18;
        end
      end
    end
    REG_8 <= (hit_ready | _T_18) & io_in_resp_ready | invalid_ready; // @[Cache.scala 282:66]
    if (reset) begin // @[Cache.scala 270:23]
      wdata1 <= 64'h0; // @[Cache.scala 270:23]
    end else if (!(4'h0 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
        if (4'h2 == state) begin // @[Cache.scala 318:18]
          wdata1 <= _GEN_989;
        end
      end
    end
    if (reset) begin // @[Cache.scala 271:23]
      wdata2 <= 64'h0; // @[Cache.scala 271:23]
    end else if (!(4'h0 == state)) begin // @[Cache.scala 318:18]
      if (!(4'h1 == state)) begin // @[Cache.scala 318:18]
        if (4'h2 == state) begin // @[Cache.scala 318:18]
          wdata2 <= _GEN_990;
        end
      end
    end
    REG_10 <= (hit_ready | _T_18) & io_in_resp_ready | invalid_ready; // @[Cache.scala 282:66]
    REG_11 <= (hit_ready | _T_18) & io_in_resp_ready | invalid_ready; // @[Cache.scala 282:66]
    if (s2_offs) begin // @[Cache.scala 410:40]
      REG_12 <= wdata2;
    end else begin
      REG_12 <= wdata1;
    end
    if (reset) begin // @[Cache.scala 438:27]
      fi_counter <= 8'h0; // @[Cache.scala 438:27]
    end else if (3'h0 == fi_state) begin // @[Cache.scala 483:23]
      if (fi_fire) begin // @[Cache.scala 485:24]
        fi_counter <= 8'h0; // @[Cache.scala 486:22]
      end
    end else if (3'h1 == fi_state) begin // @[Cache.scala 483:23]
      if (!(_GEN_3551)) begin // @[Cache.scala 498:25]
        fi_counter <= _T_611; // @[Cache.scala 501:22]
      end
    end else if (!(3'h2 == fi_state)) begin // @[Cache.scala 483:23]
      fi_counter <= _GEN_3566;
    end
    REG_13 <= fi_state == 3'h1; // @[Cache.scala 443:65]
    if (reset) begin // @[Reg.scala 27:20]
      r <= 128'h0; // @[Reg.scala 27:20]
    end else if (fi_update) begin // @[Reg.scala 28:19]
      if (2'h3 == fi_sram_idx) begin // @[Reg.scala 28:23]
        r <= sram_out_3; // @[Reg.scala 28:23]
      end else if (2'h2 == fi_sram_idx) begin // @[Reg.scala 28:23]
        r <= sram_out_2; // @[Reg.scala 28:23]
      end else begin
        r <= _GEN_3524;
      end
    end
    if (reset) begin // @[Reg.scala 27:20]
      r_1 <= 21'h0; // @[Reg.scala 27:20]
    end else if (fi_update) begin // @[Reg.scala 28:19]
      if (2'h3 == fi_sram_idx) begin // @[Reg.scala 28:23]
        r_1 <= tag_out_3; // @[Reg.scala 28:23]
      end else if (2'h2 == fi_sram_idx) begin // @[Reg.scala 28:23]
        r_1 <= tag_out_2; // @[Reg.scala 28:23]
      end else begin
        r_1 <= _GEN_3529;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  REG_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  REG_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  REG_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  REG_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  REG_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  REG_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  plru0_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  plru0_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  plru0_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  plru0_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  plru0_4 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  plru0_5 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  plru0_6 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  plru0_7 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  plru0_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  plru0_9 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  plru0_10 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  plru0_11 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  plru0_12 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  plru0_13 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  plru0_14 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  plru0_15 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  plru0_16 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  plru0_17 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  plru0_18 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  plru0_19 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  plru0_20 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  plru0_21 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  plru0_22 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  plru0_23 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  plru0_24 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  plru0_25 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  plru0_26 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  plru0_27 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  plru0_28 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  plru0_29 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  plru0_30 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  plru0_31 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  plru0_32 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  plru0_33 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  plru0_34 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  plru0_35 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  plru0_36 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  plru0_37 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  plru0_38 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  plru0_39 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  plru0_40 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  plru0_41 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  plru0_42 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  plru0_43 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  plru0_44 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  plru0_45 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  plru0_46 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  plru0_47 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  plru0_48 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  plru0_49 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  plru0_50 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  plru0_51 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  plru0_52 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  plru0_53 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  plru0_54 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  plru0_55 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  plru0_56 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  plru0_57 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  plru0_58 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  plru0_59 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  plru0_60 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  plru0_61 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  plru0_62 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  plru0_63 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  plru1_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  plru1_1 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  plru1_2 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  plru1_3 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  plru1_4 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  plru1_5 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  plru1_6 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  plru1_7 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  plru1_8 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  plru1_9 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  plru1_10 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  plru1_11 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  plru1_12 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  plru1_13 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  plru1_14 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  plru1_15 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  plru1_16 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  plru1_17 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  plru1_18 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  plru1_19 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  plru1_20 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  plru1_21 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  plru1_22 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  plru1_23 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  plru1_24 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  plru1_25 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  plru1_26 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  plru1_27 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  plru1_28 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  plru1_29 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  plru1_30 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  plru1_31 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  plru1_32 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  plru1_33 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  plru1_34 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  plru1_35 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  plru1_36 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  plru1_37 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  plru1_38 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  plru1_39 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  plru1_40 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  plru1_41 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  plru1_42 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  plru1_43 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  plru1_44 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  plru1_45 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  plru1_46 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  plru1_47 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  plru1_48 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  plru1_49 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  plru1_50 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  plru1_51 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  plru1_52 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  plru1_53 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  plru1_54 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  plru1_55 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  plru1_56 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  plru1_57 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  plru1_58 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  plru1_59 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  plru1_60 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  plru1_61 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  plru1_62 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  plru1_63 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  plru2_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  plru2_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  plru2_2 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  plru2_3 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  plru2_4 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  plru2_5 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  plru2_6 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  plru2_7 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  plru2_8 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  plru2_9 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  plru2_10 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  plru2_11 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  plru2_12 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  plru2_13 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  plru2_14 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  plru2_15 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  plru2_16 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  plru2_17 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  plru2_18 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  plru2_19 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  plru2_20 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  plru2_21 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  plru2_22 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  plru2_23 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  plru2_24 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  plru2_25 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  plru2_26 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  plru2_27 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  plru2_28 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  plru2_29 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  plru2_30 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  plru2_31 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  plru2_32 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  plru2_33 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  plru2_34 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  plru2_35 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  plru2_36 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  plru2_37 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  plru2_38 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  plru2_39 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  plru2_40 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  plru2_41 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  plru2_42 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  plru2_43 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  plru2_44 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  plru2_45 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  plru2_46 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  plru2_47 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  plru2_48 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  plru2_49 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  plru2_50 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  plru2_51 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  plru2_52 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  plru2_53 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  plru2_54 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  plru2_55 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  plru2_56 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  plru2_57 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  plru2_58 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  plru2_59 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  plru2_60 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  plru2_61 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  plru2_62 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  plru2_63 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  REG_9 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  s2_addr = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  s2_reg_hit = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  s2_wen = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  state = _RAND_204[3:0];
  _RAND_205 = {1{`RANDOM}};
  fi_valid = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  fi_state = _RAND_206[2:0];
  _RAND_207 = {2{`RANDOM}};
  s2_wdata = _RAND_207[63:0];
  _RAND_208 = {1{`RANDOM}};
  s2_wmask = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  s2_id = _RAND_209[3:0];
  _RAND_210 = {4{`RANDOM}};
  s2_reg_rdata = _RAND_210[127:0];
  _RAND_211 = {1{`RANDOM}};
  s2_reg_dirty = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  s2_reg_tag_r = _RAND_212[20:0];
  _RAND_213 = {4{`RANDOM}};
  s2_reg_dat_w = _RAND_213[127:0];
  _RAND_214 = {1{`RANDOM}};
  REG_8 = _RAND_214[0:0];
  _RAND_215 = {2{`RANDOM}};
  wdata1 = _RAND_215[63:0];
  _RAND_216 = {2{`RANDOM}};
  wdata2 = _RAND_216[63:0];
  _RAND_217 = {1{`RANDOM}};
  REG_10 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  REG_11 = _RAND_218[0:0];
  _RAND_219 = {2{`RANDOM}};
  REG_12 = _RAND_219[63:0];
  _RAND_220 = {1{`RANDOM}};
  fi_counter = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  REG_13 = _RAND_221[0:0];
  _RAND_222 = {4{`RANDOM}};
  r = _RAND_222[127:0];
  _RAND_223 = {1{`RANDOM}};
  r_1 = _RAND_223[20:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_Uncache_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [3:0]  io_in_req_bits_id,
  input  [31:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input  [1:0]  io_in_req_bits_size,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_id,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [63:0] io_out_req_bits_wdata,
  output [7:0]  io_out_req_bits_wmask,
  output        io_out_req_bits_wen,
  output [1:0]  io_out_req_bits_size,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Uncache.scala 17:22]
  reg [31:0] addr; // @[Uncache.scala 20:22]
  reg [63:0] wdata; // @[Uncache.scala 21:22]
  reg [7:0] wmask; // @[Uncache.scala 22:22]
  reg  wen; // @[Uncache.scala 23:22]
  reg [1:0] size; // @[Uncache.scala 24:22]
  reg [3:0] in_id; // @[Uncache.scala 25:22]
  reg [31:0] rdata_1; // @[Uncache.scala 29:24]
  reg [31:0] rdata_2; // @[Uncache.scala 30:24]
  wire  req_split = size == 2'h3 & addr[2:0] == 3'h0; // @[Uncache.scala 34:35]
  wire  _T_5 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_10 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _T_14 = req_split ? 3'h3 : 3'h5; // @[Uncache.scala 68:21]
  wire [31:0] _GEN_10 = _T_12 ? io_out_resp_bits_rdata[31:0] : rdata_1; // @[Uncache.scala 66:30 67:17 29:24]
  wire [2:0] _GEN_11 = _T_12 ? _T_14 : state; // @[Uncache.scala 66:30 68:15 17:22]
  wire [2:0] _GEN_12 = _T_10 ? 3'h4 : state; // @[Uncache.scala 72:29 73:15 17:22]
  wire [31:0] _GEN_13 = _T_12 ? io_out_resp_bits_rdata[31:0] : rdata_2; // @[Uncache.scala 77:30 79:19 30:24]
  wire [2:0] _GEN_14 = _T_12 ? 3'h5 : state; // @[Uncache.scala 77:30 83:15 17:22]
  wire  _T_21 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_15 = _T_21 ? 3'h0 : state; // @[Uncache.scala 87:29 88:15 17:22]
  wire [2:0] _GEN_16 = 3'h5 == state ? _GEN_15 : state; // @[Uncache.scala 36:18 17:22]
  wire [31:0] _GEN_17 = 3'h4 == state ? _GEN_13 : rdata_2; // @[Uncache.scala 36:18 30:24]
  wire [2:0] _GEN_18 = 3'h4 == state ? _GEN_14 : _GEN_16; // @[Uncache.scala 36:18]
  wire [2:0] _GEN_19 = 3'h3 == state ? _GEN_12 : _GEN_18; // @[Uncache.scala 36:18]
  wire [31:0] _GEN_20 = 3'h3 == state ? rdata_2 : _GEN_17; // @[Uncache.scala 36:18 30:24]
  wire  _T_24 = state == 3'h3; // @[Uncache.scala 98:55]
  wire [31:0] _T_34 = addr + 32'h4; // @[Uncache.scala 115:70]
  assign io_in_req_ready = state == 3'h0; // @[Uncache.scala 97:34]
  assign io_in_resp_valid = state == 3'h5; // @[Uncache.scala 106:34]
  assign io_in_resp_bits_id = in_id; // @[Uncache.scala 108:24]
  assign io_in_resp_bits_rdata = {rdata_2,rdata_1}; // @[Cat.scala 30:58]
  assign io_out_req_valid = state == 3'h1 | state == 3'h3; // @[Uncache.scala 98:46]
  assign io_out_req_bits_addr = req_split & _T_24 ? _T_34 : addr; // @[Uncache.scala 115:30]
  assign io_out_req_bits_wdata = wdata; // @[Uncache.scala 116:24]
  assign io_out_req_bits_wmask = wmask; // @[Uncache.scala 117:24]
  assign io_out_req_bits_wen = wen; // @[Uncache.scala 102:24]
  assign io_out_req_bits_size = req_split ? 2'h2 : size; // @[Uncache.scala 118:30]
  assign io_out_resp_ready = state == 3'h2 | state == 3'h4; // @[Uncache.scala 105:47]
  always @(posedge clock) begin
    if (reset) begin // @[Uncache.scala 17:22]
      state <= 3'h0; // @[Uncache.scala 17:22]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        if (~io_in_req_bits_addr[2]) begin // @[Uncache.scala 52:21]
          state <= 3'h1;
        end else begin
          state <= 3'h3;
        end
      end
    end else if (3'h1 == state) begin // @[Uncache.scala 36:18]
      if (_T_10) begin // @[Uncache.scala 61:29]
        state <= 3'h2; // @[Uncache.scala 62:15]
      end
    end else if (3'h2 == state) begin // @[Uncache.scala 36:18]
      state <= _GEN_11;
    end else begin
      state <= _GEN_19;
    end
    if (reset) begin // @[Uncache.scala 20:22]
      addr <= 32'h0; // @[Uncache.scala 20:22]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        addr <= io_in_req_bits_addr; // @[Uncache.scala 39:15]
      end
    end
    if (reset) begin // @[Uncache.scala 21:22]
      wdata <= 64'h0; // @[Uncache.scala 21:22]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        wdata <= io_in_req_bits_wdata; // @[Uncache.scala 40:15]
      end
    end
    if (reset) begin // @[Uncache.scala 22:22]
      wmask <= 8'h0; // @[Uncache.scala 22:22]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        wmask <= io_in_req_bits_wmask; // @[Uncache.scala 41:15]
      end
    end
    if (reset) begin // @[Uncache.scala 23:22]
      wen <= 1'h0; // @[Uncache.scala 23:22]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        wen <= io_in_req_bits_wen; // @[Uncache.scala 42:15]
      end
    end
    if (reset) begin // @[Uncache.scala 24:22]
      size <= 2'h0; // @[Uncache.scala 24:22]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        size <= io_in_req_bits_size; // @[Uncache.scala 43:15]
      end
    end
    if (reset) begin // @[Uncache.scala 25:22]
      in_id <= 4'h0; // @[Uncache.scala 25:22]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        in_id <= io_in_req_bits_id; // @[Uncache.scala 44:15]
      end
    end
    if (reset) begin // @[Uncache.scala 29:24]
      rdata_1 <= 32'h0; // @[Uncache.scala 29:24]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        rdata_1 <= 32'h0; // @[Uncache.scala 50:17]
      end
    end else if (!(3'h1 == state)) begin // @[Uncache.scala 36:18]
      if (3'h2 == state) begin // @[Uncache.scala 36:18]
        rdata_1 <= _GEN_10;
      end
    end
    if (reset) begin // @[Uncache.scala 30:24]
      rdata_2 <= 32'h0; // @[Uncache.scala 30:24]
    end else if (3'h0 == state) begin // @[Uncache.scala 36:18]
      if (_T_5) begin // @[Uncache.scala 38:28]
        rdata_2 <= 32'h0; // @[Uncache.scala 51:17]
      end
    end else if (!(3'h1 == state)) begin // @[Uncache.scala 36:18]
      if (!(3'h2 == state)) begin // @[Uncache.scala 36:18]
        rdata_2 <= _GEN_20;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  addr = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  wdata = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  wmask = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  wen = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  size = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  in_id = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  rdata_1 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  rdata_2 = _RAND_8[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_CacheController_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [3:0]  io_in_req_bits_id,
  input  [31:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input  [1:0]  io_in_req_bits_size,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_id,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_cache_req_ready,
  output        io_out_cache_req_valid,
  output [31:0] io_out_cache_req_bits_addr,
  output        io_out_cache_req_bits_aen,
  output [63:0] io_out_cache_req_bits_wdata,
  output        io_out_cache_req_bits_wlast,
  output        io_out_cache_req_bits_wen,
  output        io_out_cache_resp_ready,
  input         io_out_cache_resp_valid,
  input  [63:0] io_out_cache_resp_bits_rdata,
  input         io_out_cache_resp_bits_rlast,
  input         io_out_uncache_req_ready,
  output        io_out_uncache_req_valid,
  output [31:0] io_out_uncache_req_bits_addr,
  output [63:0] io_out_uncache_req_bits_wdata,
  output [7:0]  io_out_uncache_req_bits_wmask,
  output        io_out_uncache_req_bits_wen,
  output [1:0]  io_out_uncache_req_bits_size,
  output        io_out_uncache_resp_ready,
  input         io_out_uncache_resp_valid,
  input  [63:0] io_out_uncache_resp_bits_rdata,
  input         fence_i,
  output        _WIRE_10,
  input         empty
);
  wire  cache_clock; // @[CacheController.scala 14:21]
  wire  cache_reset; // @[CacheController.scala 14:21]
  wire  cache_io_in_req_ready; // @[CacheController.scala 14:21]
  wire  cache_io_in_req_valid; // @[CacheController.scala 14:21]
  wire [3:0] cache_io_in_req_bits_id; // @[CacheController.scala 14:21]
  wire [31:0] cache_io_in_req_bits_addr; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_in_req_bits_wdata; // @[CacheController.scala 14:21]
  wire [7:0] cache_io_in_req_bits_wmask; // @[CacheController.scala 14:21]
  wire  cache_io_in_req_bits_wen; // @[CacheController.scala 14:21]
  wire  cache_io_in_resp_ready; // @[CacheController.scala 14:21]
  wire  cache_io_in_resp_valid; // @[CacheController.scala 14:21]
  wire [3:0] cache_io_in_resp_bits_id; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_in_resp_bits_rdata; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_ready; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_valid; // @[CacheController.scala 14:21]
  wire [31:0] cache_io_out_req_bits_addr; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_bits_aen; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_out_req_bits_wdata; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_bits_wlast; // @[CacheController.scala 14:21]
  wire  cache_io_out_req_bits_wen; // @[CacheController.scala 14:21]
  wire  cache_io_out_resp_ready; // @[CacheController.scala 14:21]
  wire  cache_io_out_resp_valid; // @[CacheController.scala 14:21]
  wire [63:0] cache_io_out_resp_bits_rdata; // @[CacheController.scala 14:21]
  wire  cache_io_out_resp_bits_rlast; // @[CacheController.scala 14:21]
  wire  cache_fence_i_0; // @[CacheController.scala 14:21]
  wire  cache__WIRE_10_0; // @[CacheController.scala 14:21]
  wire  cache_sq_empty_0; // @[CacheController.scala 14:21]
  wire  uncache_clock; // @[CacheController.scala 15:23]
  wire  uncache_reset; // @[CacheController.scala 15:23]
  wire  uncache_io_in_req_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_in_req_valid; // @[CacheController.scala 15:23]
  wire [3:0] uncache_io_in_req_bits_id; // @[CacheController.scala 15:23]
  wire [31:0] uncache_io_in_req_bits_addr; // @[CacheController.scala 15:23]
  wire [63:0] uncache_io_in_req_bits_wdata; // @[CacheController.scala 15:23]
  wire [7:0] uncache_io_in_req_bits_wmask; // @[CacheController.scala 15:23]
  wire  uncache_io_in_req_bits_wen; // @[CacheController.scala 15:23]
  wire [1:0] uncache_io_in_req_bits_size; // @[CacheController.scala 15:23]
  wire  uncache_io_in_resp_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_in_resp_valid; // @[CacheController.scala 15:23]
  wire [3:0] uncache_io_in_resp_bits_id; // @[CacheController.scala 15:23]
  wire [63:0] uncache_io_in_resp_bits_rdata; // @[CacheController.scala 15:23]
  wire  uncache_io_out_req_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_out_req_valid; // @[CacheController.scala 15:23]
  wire [31:0] uncache_io_out_req_bits_addr; // @[CacheController.scala 15:23]
  wire [63:0] uncache_io_out_req_bits_wdata; // @[CacheController.scala 15:23]
  wire [7:0] uncache_io_out_req_bits_wmask; // @[CacheController.scala 15:23]
  wire  uncache_io_out_req_bits_wen; // @[CacheController.scala 15:23]
  wire [1:0] uncache_io_out_req_bits_size; // @[CacheController.scala 15:23]
  wire  uncache_io_out_resp_ready; // @[CacheController.scala 15:23]
  wire  uncache_io_out_resp_valid; // @[CacheController.scala 15:23]
  wire [63:0] uncache_io_out_resp_bits_rdata; // @[CacheController.scala 15:23]
  wire  crossbar1to2_clock; // @[CacheController.scala 17:28]
  wire  crossbar1to2_reset; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_req_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_req_valid; // @[CacheController.scala 17:28]
  wire [3:0] crossbar1to2_io_in_req_bits_id; // @[CacheController.scala 17:28]
  wire [31:0] crossbar1to2_io_in_req_bits_addr; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_in_req_bits_wdata; // @[CacheController.scala 17:28]
  wire [7:0] crossbar1to2_io_in_req_bits_wmask; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_req_bits_wen; // @[CacheController.scala 17:28]
  wire [1:0] crossbar1to2_io_in_req_bits_size; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_resp_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_in_resp_valid; // @[CacheController.scala 17:28]
  wire [3:0] crossbar1to2_io_in_resp_bits_id; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_in_resp_bits_rdata; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_req_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_req_valid; // @[CacheController.scala 17:28]
  wire [3:0] crossbar1to2_io_out_0_req_bits_id; // @[CacheController.scala 17:28]
  wire [31:0] crossbar1to2_io_out_0_req_bits_addr; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_out_0_req_bits_wdata; // @[CacheController.scala 17:28]
  wire [7:0] crossbar1to2_io_out_0_req_bits_wmask; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_req_bits_wen; // @[CacheController.scala 17:28]
  wire [1:0] crossbar1to2_io_out_0_req_bits_size; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_resp_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_0_resp_valid; // @[CacheController.scala 17:28]
  wire [3:0] crossbar1to2_io_out_0_resp_bits_id; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_out_0_resp_bits_rdata; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_req_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_req_valid; // @[CacheController.scala 17:28]
  wire [3:0] crossbar1to2_io_out_1_req_bits_id; // @[CacheController.scala 17:28]
  wire [31:0] crossbar1to2_io_out_1_req_bits_addr; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_out_1_req_bits_wdata; // @[CacheController.scala 17:28]
  wire [7:0] crossbar1to2_io_out_1_req_bits_wmask; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_req_bits_wen; // @[CacheController.scala 17:28]
  wire [1:0] crossbar1to2_io_out_1_req_bits_size; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_resp_ready; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_out_1_resp_valid; // @[CacheController.scala 17:28]
  wire [3:0] crossbar1to2_io_out_1_resp_bits_id; // @[CacheController.scala 17:28]
  wire [63:0] crossbar1to2_io_out_1_resp_bits_rdata; // @[CacheController.scala 17:28]
  wire  crossbar1to2_io_to_1; // @[CacheController.scala 17:28]
  ysyx_210128_Cache_1 cache ( // @[CacheController.scala 14:21]
    .clock(cache_clock),
    .reset(cache_reset),
    .io_in_req_ready(cache_io_in_req_ready),
    .io_in_req_valid(cache_io_in_req_valid),
    .io_in_req_bits_id(cache_io_in_req_bits_id),
    .io_in_req_bits_addr(cache_io_in_req_bits_addr),
    .io_in_req_bits_wdata(cache_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(cache_io_in_req_bits_wmask),
    .io_in_req_bits_wen(cache_io_in_req_bits_wen),
    .io_in_resp_ready(cache_io_in_resp_ready),
    .io_in_resp_valid(cache_io_in_resp_valid),
    .io_in_resp_bits_id(cache_io_in_resp_bits_id),
    .io_in_resp_bits_rdata(cache_io_in_resp_bits_rdata),
    .io_out_req_ready(cache_io_out_req_ready),
    .io_out_req_valid(cache_io_out_req_valid),
    .io_out_req_bits_addr(cache_io_out_req_bits_addr),
    .io_out_req_bits_aen(cache_io_out_req_bits_aen),
    .io_out_req_bits_wdata(cache_io_out_req_bits_wdata),
    .io_out_req_bits_wlast(cache_io_out_req_bits_wlast),
    .io_out_req_bits_wen(cache_io_out_req_bits_wen),
    .io_out_resp_ready(cache_io_out_resp_ready),
    .io_out_resp_valid(cache_io_out_resp_valid),
    .io_out_resp_bits_rdata(cache_io_out_resp_bits_rdata),
    .io_out_resp_bits_rlast(cache_io_out_resp_bits_rlast),
    .fence_i_0(cache_fence_i_0),
    ._WIRE_10_0(cache__WIRE_10_0),
    .sq_empty_0(cache_sq_empty_0)
  );
  ysyx_210128_Uncache_1 uncache ( // @[CacheController.scala 15:23]
    .clock(uncache_clock),
    .reset(uncache_reset),
    .io_in_req_ready(uncache_io_in_req_ready),
    .io_in_req_valid(uncache_io_in_req_valid),
    .io_in_req_bits_id(uncache_io_in_req_bits_id),
    .io_in_req_bits_addr(uncache_io_in_req_bits_addr),
    .io_in_req_bits_wdata(uncache_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(uncache_io_in_req_bits_wmask),
    .io_in_req_bits_wen(uncache_io_in_req_bits_wen),
    .io_in_req_bits_size(uncache_io_in_req_bits_size),
    .io_in_resp_ready(uncache_io_in_resp_ready),
    .io_in_resp_valid(uncache_io_in_resp_valid),
    .io_in_resp_bits_id(uncache_io_in_resp_bits_id),
    .io_in_resp_bits_rdata(uncache_io_in_resp_bits_rdata),
    .io_out_req_ready(uncache_io_out_req_ready),
    .io_out_req_valid(uncache_io_out_req_valid),
    .io_out_req_bits_addr(uncache_io_out_req_bits_addr),
    .io_out_req_bits_wdata(uncache_io_out_req_bits_wdata),
    .io_out_req_bits_wmask(uncache_io_out_req_bits_wmask),
    .io_out_req_bits_wen(uncache_io_out_req_bits_wen),
    .io_out_req_bits_size(uncache_io_out_req_bits_size),
    .io_out_resp_ready(uncache_io_out_resp_ready),
    .io_out_resp_valid(uncache_io_out_resp_valid),
    .io_out_resp_bits_rdata(uncache_io_out_resp_bits_rdata)
  );
  ysyx_210128_CacheBusCrossbar1to2_1 crossbar1to2 ( // @[CacheController.scala 17:28]
    .clock(crossbar1to2_clock),
    .reset(crossbar1to2_reset),
    .io_in_req_ready(crossbar1to2_io_in_req_ready),
    .io_in_req_valid(crossbar1to2_io_in_req_valid),
    .io_in_req_bits_id(crossbar1to2_io_in_req_bits_id),
    .io_in_req_bits_addr(crossbar1to2_io_in_req_bits_addr),
    .io_in_req_bits_wdata(crossbar1to2_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(crossbar1to2_io_in_req_bits_wmask),
    .io_in_req_bits_wen(crossbar1to2_io_in_req_bits_wen),
    .io_in_req_bits_size(crossbar1to2_io_in_req_bits_size),
    .io_in_resp_ready(crossbar1to2_io_in_resp_ready),
    .io_in_resp_valid(crossbar1to2_io_in_resp_valid),
    .io_in_resp_bits_id(crossbar1to2_io_in_resp_bits_id),
    .io_in_resp_bits_rdata(crossbar1to2_io_in_resp_bits_rdata),
    .io_out_0_req_ready(crossbar1to2_io_out_0_req_ready),
    .io_out_0_req_valid(crossbar1to2_io_out_0_req_valid),
    .io_out_0_req_bits_id(crossbar1to2_io_out_0_req_bits_id),
    .io_out_0_req_bits_addr(crossbar1to2_io_out_0_req_bits_addr),
    .io_out_0_req_bits_wdata(crossbar1to2_io_out_0_req_bits_wdata),
    .io_out_0_req_bits_wmask(crossbar1to2_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wen(crossbar1to2_io_out_0_req_bits_wen),
    .io_out_0_req_bits_size(crossbar1to2_io_out_0_req_bits_size),
    .io_out_0_resp_ready(crossbar1to2_io_out_0_resp_ready),
    .io_out_0_resp_valid(crossbar1to2_io_out_0_resp_valid),
    .io_out_0_resp_bits_id(crossbar1to2_io_out_0_resp_bits_id),
    .io_out_0_resp_bits_rdata(crossbar1to2_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(crossbar1to2_io_out_1_req_ready),
    .io_out_1_req_valid(crossbar1to2_io_out_1_req_valid),
    .io_out_1_req_bits_id(crossbar1to2_io_out_1_req_bits_id),
    .io_out_1_req_bits_addr(crossbar1to2_io_out_1_req_bits_addr),
    .io_out_1_req_bits_wdata(crossbar1to2_io_out_1_req_bits_wdata),
    .io_out_1_req_bits_wmask(crossbar1to2_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wen(crossbar1to2_io_out_1_req_bits_wen),
    .io_out_1_req_bits_size(crossbar1to2_io_out_1_req_bits_size),
    .io_out_1_resp_ready(crossbar1to2_io_out_1_resp_ready),
    .io_out_1_resp_valid(crossbar1to2_io_out_1_resp_valid),
    .io_out_1_resp_bits_id(crossbar1to2_io_out_1_resp_bits_id),
    .io_out_1_resp_bits_rdata(crossbar1to2_io_out_1_resp_bits_rdata),
    .io_to_1(crossbar1to2_io_to_1)
  );
  assign io_in_req_ready = crossbar1to2_io_in_req_ready; // @[CacheController.scala 19:22]
  assign io_in_resp_valid = crossbar1to2_io_in_resp_valid; // @[CacheController.scala 19:22]
  assign io_in_resp_bits_id = crossbar1to2_io_in_resp_bits_id; // @[CacheController.scala 19:22]
  assign io_in_resp_bits_rdata = crossbar1to2_io_in_resp_bits_rdata; // @[CacheController.scala 19:22]
  assign io_out_cache_req_valid = cache_io_out_req_valid; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_addr = cache_io_out_req_bits_addr; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_aen = cache_io_out_req_bits_aen; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_wdata = cache_io_out_req_bits_wdata; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_wlast = cache_io_out_req_bits_wlast; // @[CacheController.scala 23:16]
  assign io_out_cache_req_bits_wen = cache_io_out_req_bits_wen; // @[CacheController.scala 23:16]
  assign io_out_cache_resp_ready = cache_io_out_resp_ready; // @[CacheController.scala 23:16]
  assign io_out_uncache_req_valid = uncache_io_out_req_valid; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_addr = uncache_io_out_req_bits_addr; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_wdata = uncache_io_out_req_bits_wdata; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_wmask = uncache_io_out_req_bits_wmask; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_wen = uncache_io_out_req_bits_wen; // @[CacheController.scala 24:18]
  assign io_out_uncache_req_bits_size = uncache_io_out_req_bits_size; // @[CacheController.scala 24:18]
  assign io_out_uncache_resp_ready = uncache_io_out_resp_ready; // @[CacheController.scala 24:18]
  assign _WIRE_10 = cache__WIRE_10_0;
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_io_in_req_valid = crossbar1to2_io_out_0_req_valid; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_id = crossbar1to2_io_out_0_req_bits_id; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_addr = crossbar1to2_io_out_0_req_bits_addr; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_wdata = crossbar1to2_io_out_0_req_bits_wdata; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_wmask = crossbar1to2_io_out_0_req_bits_wmask; // @[CacheController.scala 20:26]
  assign cache_io_in_req_bits_wen = crossbar1to2_io_out_0_req_bits_wen; // @[CacheController.scala 20:26]
  assign cache_io_in_resp_ready = crossbar1to2_io_out_0_resp_ready; // @[CacheController.scala 20:26]
  assign cache_io_out_req_ready = io_out_cache_req_ready; // @[CacheController.scala 23:16]
  assign cache_io_out_resp_valid = io_out_cache_resp_valid; // @[CacheController.scala 23:16]
  assign cache_io_out_resp_bits_rdata = io_out_cache_resp_bits_rdata; // @[CacheController.scala 23:16]
  assign cache_io_out_resp_bits_rlast = io_out_cache_resp_bits_rlast; // @[CacheController.scala 23:16]
  assign cache_fence_i_0 = fence_i;
  assign cache_sq_empty_0 = empty;
  assign uncache_clock = clock;
  assign uncache_reset = reset;
  assign uncache_io_in_req_valid = crossbar1to2_io_out_1_req_valid; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_id = crossbar1to2_io_out_1_req_bits_id; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_addr = crossbar1to2_io_out_1_req_bits_addr; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_wdata = crossbar1to2_io_out_1_req_bits_wdata; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_wmask = crossbar1to2_io_out_1_req_bits_wmask; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_wen = crossbar1to2_io_out_1_req_bits_wen; // @[CacheController.scala 21:26]
  assign uncache_io_in_req_bits_size = crossbar1to2_io_out_1_req_bits_size; // @[CacheController.scala 21:26]
  assign uncache_io_in_resp_ready = crossbar1to2_io_out_1_resp_ready; // @[CacheController.scala 21:26]
  assign uncache_io_out_req_ready = io_out_uncache_req_ready; // @[CacheController.scala 24:18]
  assign uncache_io_out_resp_valid = io_out_uncache_resp_valid; // @[CacheController.scala 24:18]
  assign uncache_io_out_resp_bits_rdata = io_out_uncache_resp_bits_rdata; // @[CacheController.scala 24:18]
  assign crossbar1to2_clock = clock;
  assign crossbar1to2_reset = reset;
  assign crossbar1to2_io_in_req_valid = io_in_req_valid; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_id = io_in_req_bits_id; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_addr = io_in_req_bits_addr; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_wdata = io_in_req_bits_wdata; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_wmask = io_in_req_bits_wmask; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_wen = io_in_req_bits_wen; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_req_bits_size = io_in_req_bits_size; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_in_resp_ready = io_in_resp_ready; // @[CacheController.scala 19:22]
  assign crossbar1to2_io_out_0_req_ready = cache_io_in_req_ready; // @[CacheController.scala 20:26]
  assign crossbar1to2_io_out_0_resp_valid = cache_io_in_resp_valid; // @[CacheController.scala 20:26]
  assign crossbar1to2_io_out_0_resp_bits_id = cache_io_in_resp_bits_id; // @[CacheController.scala 20:26]
  assign crossbar1to2_io_out_0_resp_bits_rdata = cache_io_in_resp_bits_rdata; // @[CacheController.scala 20:26]
  assign crossbar1to2_io_out_1_req_ready = uncache_io_in_req_ready; // @[CacheController.scala 21:26]
  assign crossbar1to2_io_out_1_resp_valid = uncache_io_in_resp_valid; // @[CacheController.scala 21:26]
  assign crossbar1to2_io_out_1_resp_bits_id = uncache_io_in_resp_bits_id; // @[CacheController.scala 21:26]
  assign crossbar1to2_io_out_1_resp_bits_rdata = uncache_io_in_resp_bits_rdata; // @[CacheController.scala 21:26]
  assign crossbar1to2_io_to_1 = ~io_in_req_bits_addr[31]; // @[CacheController.scala 13:45]
endmodule
module ysyx_210128_Clint(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [3:0]  io_in_req_bits_id,
  input  [31:0] io_in_req_bits_addr,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wen,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_id,
  output [63:0] io_in_resp_bits_rdata,
  output        mtip_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime; // @[Clint.scala 12:22]
  reg [63:0] mtimecmp; // @[Clint.scala 13:25]
  reg [63:0] clint_freq; // @[Clint.scala 17:27]
  reg [63:0] clint_step; // @[Clint.scala 18:27]
  reg [63:0] counter; // @[Clint.scala 20:24]
  wire [63:0] counter_next = counter + 64'h1; // @[Clint.scala 21:30]
  wire [63:0] _T_5 = mtime + clint_step; // @[Clint.scala 24:20]
  wire [15:0] addr = io_in_req_bits_addr[15:0]; // @[Clint.scala 35:33]
  wire [7:0] _T_15 = io_in_req_bits_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_17 = io_in_req_bits_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_19 = io_in_req_bits_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_21 = io_in_req_bits_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_23 = io_in_req_bits_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_25 = io_in_req_bits_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_27 = io_in_req_bits_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_29 = io_in_req_bits_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] wmask = {_T_29,_T_27,_T_25,_T_23,_T_21,_T_19,_T_17,_T_15}; // @[Cat.scala 30:58]
  wire  _T_30 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_31 = io_in_req_bits_wen & _T_30; // @[Clint.scala 41:59]
  wire  _T_32 = addr == 16'h4000; // @[RegMap.scala 14:18]
  wire [63:0] _GEN_1 = addr == 16'h4000 ? mtimecmp : 64'h0; // @[RegMap.scala 14:25 15:15]
  wire [63:0] _T_35 = io_in_req_bits_wdata & wmask; // @[Utils.scala 20:15]
  wire [63:0] _T_36 = ~wmask; // @[Utils.scala 20:37]
  wire [63:0] _T_37 = mtimecmp & _T_36; // @[Utils.scala 20:35]
  wire [63:0] _T_38 = _T_35 | _T_37; // @[Utils.scala 20:23]
  wire  _T_39 = addr == 16'h8000; // @[RegMap.scala 14:18]
  wire [63:0] _GEN_3 = addr == 16'h8000 ? clint_freq : _GEN_1; // @[RegMap.scala 14:25 15:15]
  wire [63:0] _T_44 = clint_freq & _T_36; // @[Utils.scala 20:35]
  wire [63:0] _T_45 = _T_35 | _T_44; // @[Utils.scala 20:23]
  wire  _T_46 = addr == 16'h8008; // @[RegMap.scala 14:18]
  wire [63:0] _GEN_5 = addr == 16'h8008 ? clint_step : _GEN_3; // @[RegMap.scala 14:25 15:15]
  wire [63:0] _T_51 = clint_step & _T_36; // @[Utils.scala 20:35]
  wire [63:0] _T_52 = _T_35 | _T_51; // @[Utils.scala 20:23]
  wire  _T_53 = addr == 16'hbff8; // @[RegMap.scala 14:18]
  wire [63:0] rdata = addr == 16'hbff8 ? mtime : _GEN_5; // @[RegMap.scala 14:25 15:15]
  wire [63:0] _T_58 = mtime & _T_36; // @[Utils.scala 20:35]
  wire [63:0] _T_59 = _T_35 | _T_58; // @[Utils.scala 20:23]
  reg [63:0] reg_rdata; // @[Clint.scala 43:26]
  reg [3:0] reg_id; // @[Clint.scala 44:23]
  reg  state; // @[Clint.scala 48:22]
  wire  _GEN_13 = _T_30 | state; // @[Clint.scala 52:31 59:15 48:22]
  wire  _T_63 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 40:37]
  wire  mtip = mtime >= mtimecmp; // @[Clint.scala 75:18]
  assign io_in_req_ready = ~state; // @[Clint.scala 69:29]
  assign io_in_resp_valid = state; // @[Clint.scala 70:30]
  assign io_in_resp_bits_id = reg_id; // @[Clint.scala 72:22]
  assign io_in_resp_bits_rdata = reg_rdata; // @[Clint.scala 71:25]
  assign mtip_1 = mtip;
  always @(posedge clock) begin
    if (reset) begin // @[Clint.scala 12:22]
      mtime <= 64'h0; // @[Clint.scala 12:22]
    end else if (_T_53 & _T_31) begin // @[RegMap.scala 18:34]
      mtime <= _T_59; // @[RegMap.scala 19:13]
    end else if (counter_next == clint_freq) begin // @[Clint.scala 23:38]
      mtime <= _T_5; // @[Clint.scala 24:11]
    end
    if (reset) begin // @[Clint.scala 13:25]
      mtimecmp <= 64'h0; // @[Clint.scala 13:25]
    end else if (_T_32 & _T_31) begin // @[RegMap.scala 18:34]
      mtimecmp <= _T_38; // @[RegMap.scala 19:13]
    end
    if (reset) begin // @[Clint.scala 17:27]
      clint_freq <= 64'h1; // @[Clint.scala 17:27]
    end else if (_T_39 & _T_31) begin // @[RegMap.scala 18:34]
      clint_freq <= _T_45; // @[RegMap.scala 19:13]
    end
    if (reset) begin // @[Clint.scala 18:27]
      clint_step <= 64'h1; // @[Clint.scala 18:27]
    end else if (_T_46 & _T_31) begin // @[RegMap.scala 18:34]
      clint_step <= _T_52; // @[RegMap.scala 19:13]
    end
    if (reset) begin // @[Clint.scala 20:24]
      counter <= 64'h0; // @[Clint.scala 20:24]
    end else if (counter_next < clint_freq) begin // @[Clint.scala 22:17]
      counter <= counter_next;
    end else begin
      counter <= 64'h0;
    end
    if (reset) begin // @[Clint.scala 43:26]
      reg_rdata <= 64'h0; // @[Clint.scala 43:26]
    end else if (~state) begin // @[Clint.scala 50:18]
      if (_T_30) begin // @[Clint.scala 52:31]
        if (!(io_in_req_bits_wen)) begin // @[Clint.scala 53:20]
          reg_rdata <= rdata; // @[Clint.scala 56:21]
        end
      end
    end
    if (reset) begin // @[Clint.scala 44:23]
      reg_id <= 4'h0; // @[Clint.scala 44:23]
    end else if (~state) begin // @[Clint.scala 50:18]
      if (_T_30) begin // @[Clint.scala 52:31]
        reg_id <= io_in_req_bits_id;
      end
    end
    if (reset) begin // @[Clint.scala 48:22]
      state <= 1'h0; // @[Clint.scala 48:22]
    end else if (~state) begin // @[Clint.scala 50:18]
      state <= _GEN_13;
    end else if (state) begin // @[Clint.scala 50:18]
      if (_T_63) begin // @[Clint.scala 63:32]
        state <= 1'h0; // @[Clint.scala 64:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  clint_freq = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  clint_step = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  counter = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  reg_rdata = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  reg_id = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_Core(
  input         clock,
  input         reset,
  input         io_core_bus_0_req_ready,
  output        io_core_bus_0_req_valid,
  output [31:0] io_core_bus_0_req_bits_addr,
  output        io_core_bus_0_req_bits_aen,
  output [63:0] io_core_bus_0_req_bits_wdata,
  output        io_core_bus_0_req_bits_wlast,
  output        io_core_bus_0_req_bits_wen,
  output        io_core_bus_0_resp_ready,
  input         io_core_bus_0_resp_valid,
  input  [63:0] io_core_bus_0_resp_bits_rdata,
  input         io_core_bus_0_resp_bits_rlast,
  input         io_core_bus_1_req_ready,
  output        io_core_bus_1_req_valid,
  output [31:0] io_core_bus_1_req_bits_addr,
  output        io_core_bus_1_req_bits_aen,
  output [63:0] io_core_bus_1_req_bits_wdata,
  output        io_core_bus_1_req_bits_wlast,
  output        io_core_bus_1_req_bits_wen,
  output        io_core_bus_1_resp_ready,
  input         io_core_bus_1_resp_valid,
  input  [63:0] io_core_bus_1_resp_bits_rdata,
  input         io_core_bus_1_resp_bits_rlast,
  input         io_core_bus_2_req_ready,
  output        io_core_bus_2_req_valid,
  output [31:0] io_core_bus_2_req_bits_addr,
  output [1:0]  io_core_bus_2_req_bits_size,
  output        io_core_bus_2_resp_ready,
  input         io_core_bus_2_resp_valid,
  input  [63:0] io_core_bus_2_resp_bits_rdata,
  input         io_core_bus_3_req_ready,
  output        io_core_bus_3_req_valid,
  output [31:0] io_core_bus_3_req_bits_addr,
  output [63:0] io_core_bus_3_req_bits_wdata,
  output [7:0]  io_core_bus_3_req_bits_wmask,
  output        io_core_bus_3_req_bits_wen,
  output [1:0]  io_core_bus_3_req_bits_size,
  output        io_core_bus_3_resp_ready,
  input         io_core_bus_3_resp_valid,
  input  [63:0] io_core_bus_3_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  fetch_clock; // @[Core.scala 17:21]
  wire  fetch_reset; // @[Core.scala 17:21]
  wire  fetch_io_imem_req_ready; // @[Core.scala 17:21]
  wire  fetch_io_imem_req_valid; // @[Core.scala 17:21]
  wire [31:0] fetch_io_imem_req_bits_addr; // @[Core.scala 17:21]
  wire [67:0] fetch_io_imem_req_bits_user; // @[Core.scala 17:21]
  wire  fetch_io_imem_resp_ready; // @[Core.scala 17:21]
  wire  fetch_io_imem_resp_valid; // @[Core.scala 17:21]
  wire [63:0] fetch_io_imem_resp_bits_rdata; // @[Core.scala 17:21]
  wire [67:0] fetch_io_imem_resp_bits_user; // @[Core.scala 17:21]
  wire  fetch_io_jmp_packet_valid; // @[Core.scala 17:21]
  wire [31:0] fetch_io_jmp_packet_inst_pc; // @[Core.scala 17:21]
  wire  fetch_io_jmp_packet_jmp; // @[Core.scala 17:21]
  wire [31:0] fetch_io_jmp_packet_jmp_pc; // @[Core.scala 17:21]
  wire  fetch_io_jmp_packet_mis; // @[Core.scala 17:21]
  wire  fetch_io_jmp_packet_sys; // @[Core.scala 17:21]
  wire  fetch_io_out_ready; // @[Core.scala 17:21]
  wire  fetch_io_out_valid; // @[Core.scala 17:21]
  wire [31:0] fetch_io_out_bits_vec_0_pc; // @[Core.scala 17:21]
  wire [31:0] fetch_io_out_bits_vec_0_inst; // @[Core.scala 17:21]
  wire  fetch_io_out_bits_vec_0_pred_br; // @[Core.scala 17:21]
  wire [31:0] fetch_io_out_bits_vec_0_pred_bpc; // @[Core.scala 17:21]
  wire  fetch_io_out_bits_vec_0_valid; // @[Core.scala 17:21]
  wire [31:0] fetch_io_out_bits_vec_1_pc; // @[Core.scala 17:21]
  wire [31:0] fetch_io_out_bits_vec_1_inst; // @[Core.scala 17:21]
  wire  fetch_io_out_bits_vec_1_pred_br; // @[Core.scala 17:21]
  wire [31:0] fetch_io_out_bits_vec_1_pred_bpc; // @[Core.scala 17:21]
  wire  fetch_io_out_bits_vec_1_valid; // @[Core.scala 17:21]
  wire  icache_clock; // @[Core.scala 19:22]
  wire  icache_reset; // @[Core.scala 19:22]
  wire  icache_io_in_req_ready; // @[Core.scala 19:22]
  wire  icache_io_in_req_valid; // @[Core.scala 19:22]
  wire [31:0] icache_io_in_req_bits_addr; // @[Core.scala 19:22]
  wire [67:0] icache_io_in_req_bits_user; // @[Core.scala 19:22]
  wire  icache_io_in_resp_ready; // @[Core.scala 19:22]
  wire  icache_io_in_resp_valid; // @[Core.scala 19:22]
  wire [63:0] icache_io_in_resp_bits_rdata; // @[Core.scala 19:22]
  wire [67:0] icache_io_in_resp_bits_user; // @[Core.scala 19:22]
  wire  icache_io_out_cache_req_ready; // @[Core.scala 19:22]
  wire  icache_io_out_cache_req_valid; // @[Core.scala 19:22]
  wire [31:0] icache_io_out_cache_req_bits_addr; // @[Core.scala 19:22]
  wire  icache_io_out_cache_req_bits_aen; // @[Core.scala 19:22]
  wire [63:0] icache_io_out_cache_req_bits_wdata; // @[Core.scala 19:22]
  wire  icache_io_out_cache_req_bits_wlast; // @[Core.scala 19:22]
  wire  icache_io_out_cache_req_bits_wen; // @[Core.scala 19:22]
  wire  icache_io_out_cache_resp_ready; // @[Core.scala 19:22]
  wire  icache_io_out_cache_resp_valid; // @[Core.scala 19:22]
  wire [63:0] icache_io_out_cache_resp_bits_rdata; // @[Core.scala 19:22]
  wire  icache_io_out_cache_resp_bits_rlast; // @[Core.scala 19:22]
  wire  icache_io_out_uncache_req_ready; // @[Core.scala 19:22]
  wire  icache_io_out_uncache_req_valid; // @[Core.scala 19:22]
  wire [31:0] icache_io_out_uncache_req_bits_addr; // @[Core.scala 19:22]
  wire [1:0] icache_io_out_uncache_req_bits_size; // @[Core.scala 19:22]
  wire  icache_io_out_uncache_resp_ready; // @[Core.scala 19:22]
  wire  icache_io_out_uncache_resp_valid; // @[Core.scala 19:22]
  wire [63:0] icache_io_out_uncache_resp_bits_rdata; // @[Core.scala 19:22]
  wire  icache_fence_i; // @[Core.scala 19:22]
  wire  icache__WIRE_10; // @[Core.scala 19:22]
  wire  icache_empty; // @[Core.scala 19:22]
  wire  ibuf_clock; // @[Core.scala 26:20]
  wire  ibuf_reset; // @[Core.scala 26:20]
  wire  ibuf_io_in_ready; // @[Core.scala 26:20]
  wire  ibuf_io_in_valid; // @[Core.scala 26:20]
  wire [31:0] ibuf_io_in_bits_vec_0_pc; // @[Core.scala 26:20]
  wire [31:0] ibuf_io_in_bits_vec_0_inst; // @[Core.scala 26:20]
  wire  ibuf_io_in_bits_vec_0_pred_br; // @[Core.scala 26:20]
  wire [31:0] ibuf_io_in_bits_vec_0_pred_bpc; // @[Core.scala 26:20]
  wire  ibuf_io_in_bits_vec_0_valid; // @[Core.scala 26:20]
  wire [31:0] ibuf_io_in_bits_vec_1_pc; // @[Core.scala 26:20]
  wire [31:0] ibuf_io_in_bits_vec_1_inst; // @[Core.scala 26:20]
  wire  ibuf_io_in_bits_vec_1_pred_br; // @[Core.scala 26:20]
  wire [31:0] ibuf_io_in_bits_vec_1_pred_bpc; // @[Core.scala 26:20]
  wire  ibuf_io_in_bits_vec_1_valid; // @[Core.scala 26:20]
  wire  ibuf_io_out_ready; // @[Core.scala 26:20]
  wire  ibuf_io_out_valid; // @[Core.scala 26:20]
  wire [31:0] ibuf_io_out_bits_vec_0_pc; // @[Core.scala 26:20]
  wire [31:0] ibuf_io_out_bits_vec_0_inst; // @[Core.scala 26:20]
  wire  ibuf_io_out_bits_vec_0_pred_br; // @[Core.scala 26:20]
  wire [31:0] ibuf_io_out_bits_vec_0_pred_bpc; // @[Core.scala 26:20]
  wire  ibuf_io_out_bits_vec_0_valid; // @[Core.scala 26:20]
  wire [31:0] ibuf_io_out_bits_vec_1_pc; // @[Core.scala 26:20]
  wire [31:0] ibuf_io_out_bits_vec_1_inst; // @[Core.scala 26:20]
  wire  ibuf_io_out_bits_vec_1_pred_br; // @[Core.scala 26:20]
  wire [31:0] ibuf_io_out_bits_vec_1_pred_bpc; // @[Core.scala 26:20]
  wire  ibuf_io_out_bits_vec_1_valid; // @[Core.scala 26:20]
  wire  ibuf_io_flush; // @[Core.scala 26:20]
  wire  decode_clock; // @[Core.scala 32:22]
  wire  decode_reset; // @[Core.scala 32:22]
  wire  decode_io_in_ready; // @[Core.scala 32:22]
  wire  decode_io_in_valid; // @[Core.scala 32:22]
  wire [31:0] decode_io_in_bits_vec_0_pc; // @[Core.scala 32:22]
  wire [31:0] decode_io_in_bits_vec_0_inst; // @[Core.scala 32:22]
  wire  decode_io_in_bits_vec_0_pred_br; // @[Core.scala 32:22]
  wire [31:0] decode_io_in_bits_vec_0_pred_bpc; // @[Core.scala 32:22]
  wire  decode_io_in_bits_vec_0_valid; // @[Core.scala 32:22]
  wire [31:0] decode_io_in_bits_vec_1_pc; // @[Core.scala 32:22]
  wire [31:0] decode_io_in_bits_vec_1_inst; // @[Core.scala 32:22]
  wire  decode_io_in_bits_vec_1_pred_br; // @[Core.scala 32:22]
  wire [31:0] decode_io_in_bits_vec_1_pred_bpc; // @[Core.scala 32:22]
  wire  decode_io_in_bits_vec_1_valid; // @[Core.scala 32:22]
  wire  decode_io_out_ready; // @[Core.scala 32:22]
  wire  decode_io_out_valid; // @[Core.scala 32:22]
  wire  decode_io_out_bits_vec_0_valid; // @[Core.scala 32:22]
  wire [31:0] decode_io_out_bits_vec_0_pc; // @[Core.scala 32:22]
  wire [31:0] decode_io_out_bits_vec_0_npc; // @[Core.scala 32:22]
  wire [31:0] decode_io_out_bits_vec_0_inst; // @[Core.scala 32:22]
  wire [2:0] decode_io_out_bits_vec_0_fu_code; // @[Core.scala 32:22]
  wire [3:0] decode_io_out_bits_vec_0_alu_code; // @[Core.scala 32:22]
  wire [3:0] decode_io_out_bits_vec_0_jmp_code; // @[Core.scala 32:22]
  wire [1:0] decode_io_out_bits_vec_0_mem_code; // @[Core.scala 32:22]
  wire [1:0] decode_io_out_bits_vec_0_mem_size; // @[Core.scala 32:22]
  wire [2:0] decode_io_out_bits_vec_0_sys_code; // @[Core.scala 32:22]
  wire  decode_io_out_bits_vec_0_w_type; // @[Core.scala 32:22]
  wire [1:0] decode_io_out_bits_vec_0_rs1_src; // @[Core.scala 32:22]
  wire [1:0] decode_io_out_bits_vec_0_rs2_src; // @[Core.scala 32:22]
  wire [4:0] decode_io_out_bits_vec_0_rs1_addr; // @[Core.scala 32:22]
  wire [4:0] decode_io_out_bits_vec_0_rs2_addr; // @[Core.scala 32:22]
  wire [4:0] decode_io_out_bits_vec_0_rd_addr; // @[Core.scala 32:22]
  wire  decode_io_out_bits_vec_0_rd_en; // @[Core.scala 32:22]
  wire [31:0] decode_io_out_bits_vec_0_imm; // @[Core.scala 32:22]
  wire  decode_io_out_bits_vec_0_pred_br; // @[Core.scala 32:22]
  wire [31:0] decode_io_out_bits_vec_0_pred_bpc; // @[Core.scala 32:22]
  wire  decode_io_out_bits_vec_1_valid; // @[Core.scala 32:22]
  wire [31:0] decode_io_out_bits_vec_1_pc; // @[Core.scala 32:22]
  wire [31:0] decode_io_out_bits_vec_1_npc; // @[Core.scala 32:22]
  wire [31:0] decode_io_out_bits_vec_1_inst; // @[Core.scala 32:22]
  wire [2:0] decode_io_out_bits_vec_1_fu_code; // @[Core.scala 32:22]
  wire [3:0] decode_io_out_bits_vec_1_alu_code; // @[Core.scala 32:22]
  wire [3:0] decode_io_out_bits_vec_1_jmp_code; // @[Core.scala 32:22]
  wire [1:0] decode_io_out_bits_vec_1_mem_code; // @[Core.scala 32:22]
  wire [1:0] decode_io_out_bits_vec_1_mem_size; // @[Core.scala 32:22]
  wire [2:0] decode_io_out_bits_vec_1_sys_code; // @[Core.scala 32:22]
  wire  decode_io_out_bits_vec_1_w_type; // @[Core.scala 32:22]
  wire [1:0] decode_io_out_bits_vec_1_rs1_src; // @[Core.scala 32:22]
  wire [1:0] decode_io_out_bits_vec_1_rs2_src; // @[Core.scala 32:22]
  wire [4:0] decode_io_out_bits_vec_1_rs1_addr; // @[Core.scala 32:22]
  wire [4:0] decode_io_out_bits_vec_1_rs2_addr; // @[Core.scala 32:22]
  wire [4:0] decode_io_out_bits_vec_1_rd_addr; // @[Core.scala 32:22]
  wire  decode_io_out_bits_vec_1_rd_en; // @[Core.scala 32:22]
  wire [31:0] decode_io_out_bits_vec_1_imm; // @[Core.scala 32:22]
  wire  decode_io_out_bits_vec_1_pred_br; // @[Core.scala 32:22]
  wire [31:0] decode_io_out_bits_vec_1_pred_bpc; // @[Core.scala 32:22]
  wire  decode_io_flush; // @[Core.scala 32:22]
  wire  rename_clock; // @[Core.scala 36:22]
  wire  rename_reset; // @[Core.scala 36:22]
  wire  rename_io_in_ready; // @[Core.scala 36:22]
  wire  rename_io_in_valid; // @[Core.scala 36:22]
  wire  rename_io_in_bits_vec_0_valid; // @[Core.scala 36:22]
  wire [31:0] rename_io_in_bits_vec_0_pc; // @[Core.scala 36:22]
  wire [31:0] rename_io_in_bits_vec_0_npc; // @[Core.scala 36:22]
  wire [31:0] rename_io_in_bits_vec_0_inst; // @[Core.scala 36:22]
  wire [2:0] rename_io_in_bits_vec_0_fu_code; // @[Core.scala 36:22]
  wire [3:0] rename_io_in_bits_vec_0_alu_code; // @[Core.scala 36:22]
  wire [3:0] rename_io_in_bits_vec_0_jmp_code; // @[Core.scala 36:22]
  wire [1:0] rename_io_in_bits_vec_0_mem_code; // @[Core.scala 36:22]
  wire [1:0] rename_io_in_bits_vec_0_mem_size; // @[Core.scala 36:22]
  wire [2:0] rename_io_in_bits_vec_0_sys_code; // @[Core.scala 36:22]
  wire  rename_io_in_bits_vec_0_w_type; // @[Core.scala 36:22]
  wire [1:0] rename_io_in_bits_vec_0_rs1_src; // @[Core.scala 36:22]
  wire [1:0] rename_io_in_bits_vec_0_rs2_src; // @[Core.scala 36:22]
  wire [4:0] rename_io_in_bits_vec_0_rs1_addr; // @[Core.scala 36:22]
  wire [4:0] rename_io_in_bits_vec_0_rs2_addr; // @[Core.scala 36:22]
  wire [4:0] rename_io_in_bits_vec_0_rd_addr; // @[Core.scala 36:22]
  wire  rename_io_in_bits_vec_0_rd_en; // @[Core.scala 36:22]
  wire [31:0] rename_io_in_bits_vec_0_imm; // @[Core.scala 36:22]
  wire  rename_io_in_bits_vec_0_pred_br; // @[Core.scala 36:22]
  wire [31:0] rename_io_in_bits_vec_0_pred_bpc; // @[Core.scala 36:22]
  wire  rename_io_in_bits_vec_1_valid; // @[Core.scala 36:22]
  wire [31:0] rename_io_in_bits_vec_1_pc; // @[Core.scala 36:22]
  wire [31:0] rename_io_in_bits_vec_1_npc; // @[Core.scala 36:22]
  wire [31:0] rename_io_in_bits_vec_1_inst; // @[Core.scala 36:22]
  wire [2:0] rename_io_in_bits_vec_1_fu_code; // @[Core.scala 36:22]
  wire [3:0] rename_io_in_bits_vec_1_alu_code; // @[Core.scala 36:22]
  wire [3:0] rename_io_in_bits_vec_1_jmp_code; // @[Core.scala 36:22]
  wire [1:0] rename_io_in_bits_vec_1_mem_code; // @[Core.scala 36:22]
  wire [1:0] rename_io_in_bits_vec_1_mem_size; // @[Core.scala 36:22]
  wire [2:0] rename_io_in_bits_vec_1_sys_code; // @[Core.scala 36:22]
  wire  rename_io_in_bits_vec_1_w_type; // @[Core.scala 36:22]
  wire [1:0] rename_io_in_bits_vec_1_rs1_src; // @[Core.scala 36:22]
  wire [1:0] rename_io_in_bits_vec_1_rs2_src; // @[Core.scala 36:22]
  wire [4:0] rename_io_in_bits_vec_1_rs1_addr; // @[Core.scala 36:22]
  wire [4:0] rename_io_in_bits_vec_1_rs2_addr; // @[Core.scala 36:22]
  wire [4:0] rename_io_in_bits_vec_1_rd_addr; // @[Core.scala 36:22]
  wire  rename_io_in_bits_vec_1_rd_en; // @[Core.scala 36:22]
  wire [31:0] rename_io_in_bits_vec_1_imm; // @[Core.scala 36:22]
  wire  rename_io_in_bits_vec_1_pred_br; // @[Core.scala 36:22]
  wire [31:0] rename_io_in_bits_vec_1_pred_bpc; // @[Core.scala 36:22]
  wire  rename_io_out_ready; // @[Core.scala 36:22]
  wire  rename_io_out_valid; // @[Core.scala 36:22]
  wire  rename_io_out_bits_vec_0_valid; // @[Core.scala 36:22]
  wire [31:0] rename_io_out_bits_vec_0_pc; // @[Core.scala 36:22]
  wire [31:0] rename_io_out_bits_vec_0_npc; // @[Core.scala 36:22]
  wire [31:0] rename_io_out_bits_vec_0_inst; // @[Core.scala 36:22]
  wire [2:0] rename_io_out_bits_vec_0_fu_code; // @[Core.scala 36:22]
  wire [3:0] rename_io_out_bits_vec_0_alu_code; // @[Core.scala 36:22]
  wire [3:0] rename_io_out_bits_vec_0_jmp_code; // @[Core.scala 36:22]
  wire [1:0] rename_io_out_bits_vec_0_mem_code; // @[Core.scala 36:22]
  wire [1:0] rename_io_out_bits_vec_0_mem_size; // @[Core.scala 36:22]
  wire [2:0] rename_io_out_bits_vec_0_sys_code; // @[Core.scala 36:22]
  wire  rename_io_out_bits_vec_0_w_type; // @[Core.scala 36:22]
  wire [1:0] rename_io_out_bits_vec_0_rs1_src; // @[Core.scala 36:22]
  wire [1:0] rename_io_out_bits_vec_0_rs2_src; // @[Core.scala 36:22]
  wire [4:0] rename_io_out_bits_vec_0_rd_addr; // @[Core.scala 36:22]
  wire  rename_io_out_bits_vec_0_rd_en; // @[Core.scala 36:22]
  wire [31:0] rename_io_out_bits_vec_0_imm; // @[Core.scala 36:22]
  wire  rename_io_out_bits_vec_0_pred_br; // @[Core.scala 36:22]
  wire [31:0] rename_io_out_bits_vec_0_pred_bpc; // @[Core.scala 36:22]
  wire [5:0] rename_io_out_bits_vec_0_rs1_paddr; // @[Core.scala 36:22]
  wire [5:0] rename_io_out_bits_vec_0_rs2_paddr; // @[Core.scala 36:22]
  wire [5:0] rename_io_out_bits_vec_0_rd_paddr; // @[Core.scala 36:22]
  wire [5:0] rename_io_out_bits_vec_0_rd_ppaddr; // @[Core.scala 36:22]
  wire  rename_io_out_bits_vec_1_valid; // @[Core.scala 36:22]
  wire [31:0] rename_io_out_bits_vec_1_pc; // @[Core.scala 36:22]
  wire [31:0] rename_io_out_bits_vec_1_npc; // @[Core.scala 36:22]
  wire [31:0] rename_io_out_bits_vec_1_inst; // @[Core.scala 36:22]
  wire [2:0] rename_io_out_bits_vec_1_fu_code; // @[Core.scala 36:22]
  wire [3:0] rename_io_out_bits_vec_1_alu_code; // @[Core.scala 36:22]
  wire [3:0] rename_io_out_bits_vec_1_jmp_code; // @[Core.scala 36:22]
  wire [1:0] rename_io_out_bits_vec_1_mem_code; // @[Core.scala 36:22]
  wire [1:0] rename_io_out_bits_vec_1_mem_size; // @[Core.scala 36:22]
  wire [2:0] rename_io_out_bits_vec_1_sys_code; // @[Core.scala 36:22]
  wire  rename_io_out_bits_vec_1_w_type; // @[Core.scala 36:22]
  wire [1:0] rename_io_out_bits_vec_1_rs1_src; // @[Core.scala 36:22]
  wire [1:0] rename_io_out_bits_vec_1_rs2_src; // @[Core.scala 36:22]
  wire [4:0] rename_io_out_bits_vec_1_rd_addr; // @[Core.scala 36:22]
  wire  rename_io_out_bits_vec_1_rd_en; // @[Core.scala 36:22]
  wire [31:0] rename_io_out_bits_vec_1_imm; // @[Core.scala 36:22]
  wire  rename_io_out_bits_vec_1_pred_br; // @[Core.scala 36:22]
  wire [31:0] rename_io_out_bits_vec_1_pred_bpc; // @[Core.scala 36:22]
  wire [5:0] rename_io_out_bits_vec_1_rs1_paddr; // @[Core.scala 36:22]
  wire [5:0] rename_io_out_bits_vec_1_rs2_paddr; // @[Core.scala 36:22]
  wire [5:0] rename_io_out_bits_vec_1_rd_paddr; // @[Core.scala 36:22]
  wire [5:0] rename_io_out_bits_vec_1_rd_ppaddr; // @[Core.scala 36:22]
  wire [63:0] rename_io_avail_list; // @[Core.scala 36:22]
  wire  rename_io_flush; // @[Core.scala 36:22]
  wire  rename_io_exe_0_valid; // @[Core.scala 36:22]
  wire  rename_io_exe_0_rd_en; // @[Core.scala 36:22]
  wire [5:0] rename_io_exe_0_rd_paddr; // @[Core.scala 36:22]
  wire  rename_io_exe_1_valid; // @[Core.scala 36:22]
  wire  rename_io_exe_1_rd_en; // @[Core.scala 36:22]
  wire [5:0] rename_io_exe_1_rd_paddr; // @[Core.scala 36:22]
  wire  rename_io_exe_2_valid; // @[Core.scala 36:22]
  wire  rename_io_exe_2_rd_en; // @[Core.scala 36:22]
  wire [5:0] rename_io_exe_2_rd_paddr; // @[Core.scala 36:22]
  wire  rename_io_cm_recover; // @[Core.scala 36:22]
  wire  rename_io_cm_0_valid; // @[Core.scala 36:22]
  wire [4:0] rename_io_cm_0_rd_addr; // @[Core.scala 36:22]
  wire  rename_io_cm_0_rd_en; // @[Core.scala 36:22]
  wire [5:0] rename_io_cm_0_rd_paddr; // @[Core.scala 36:22]
  wire [5:0] rename_io_cm_0_rd_ppaddr; // @[Core.scala 36:22]
  wire  rename_io_cm_1_valid; // @[Core.scala 36:22]
  wire [4:0] rename_io_cm_1_rd_addr; // @[Core.scala 36:22]
  wire  rename_io_cm_1_rd_en; // @[Core.scala 36:22]
  wire [5:0] rename_io_cm_1_rd_paddr; // @[Core.scala 36:22]
  wire [5:0] rename_io_cm_1_rd_ppaddr; // @[Core.scala 36:22]
  wire  stall_reg_clock; // @[Core.scala 42:25]
  wire  stall_reg_reset; // @[Core.scala 42:25]
  wire  stall_reg_io_flush; // @[Core.scala 42:25]
  wire  stall_reg_io_in_ready; // @[Core.scala 42:25]
  wire  stall_reg_io_in_valid; // @[Core.scala 42:25]
  wire  stall_reg_io_in_bits_vec_0_valid; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_in_bits_vec_0_pc; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_in_bits_vec_0_npc; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_in_bits_vec_0_inst; // @[Core.scala 42:25]
  wire [2:0] stall_reg_io_in_bits_vec_0_fu_code; // @[Core.scala 42:25]
  wire [3:0] stall_reg_io_in_bits_vec_0_alu_code; // @[Core.scala 42:25]
  wire [3:0] stall_reg_io_in_bits_vec_0_jmp_code; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_in_bits_vec_0_mem_code; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_in_bits_vec_0_mem_size; // @[Core.scala 42:25]
  wire [2:0] stall_reg_io_in_bits_vec_0_sys_code; // @[Core.scala 42:25]
  wire  stall_reg_io_in_bits_vec_0_w_type; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_in_bits_vec_0_rs1_src; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_in_bits_vec_0_rs2_src; // @[Core.scala 42:25]
  wire [4:0] stall_reg_io_in_bits_vec_0_rd_addr; // @[Core.scala 42:25]
  wire  stall_reg_io_in_bits_vec_0_rd_en; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_in_bits_vec_0_imm; // @[Core.scala 42:25]
  wire  stall_reg_io_in_bits_vec_0_pred_br; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_in_bits_vec_0_pred_bpc; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_in_bits_vec_0_rs1_paddr; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_in_bits_vec_0_rs2_paddr; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_in_bits_vec_0_rd_paddr; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_in_bits_vec_0_rd_ppaddr; // @[Core.scala 42:25]
  wire  stall_reg_io_in_bits_vec_1_valid; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_in_bits_vec_1_pc; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_in_bits_vec_1_npc; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_in_bits_vec_1_inst; // @[Core.scala 42:25]
  wire [2:0] stall_reg_io_in_bits_vec_1_fu_code; // @[Core.scala 42:25]
  wire [3:0] stall_reg_io_in_bits_vec_1_alu_code; // @[Core.scala 42:25]
  wire [3:0] stall_reg_io_in_bits_vec_1_jmp_code; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_in_bits_vec_1_mem_code; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_in_bits_vec_1_mem_size; // @[Core.scala 42:25]
  wire [2:0] stall_reg_io_in_bits_vec_1_sys_code; // @[Core.scala 42:25]
  wire  stall_reg_io_in_bits_vec_1_w_type; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_in_bits_vec_1_rs1_src; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_in_bits_vec_1_rs2_src; // @[Core.scala 42:25]
  wire [4:0] stall_reg_io_in_bits_vec_1_rd_addr; // @[Core.scala 42:25]
  wire  stall_reg_io_in_bits_vec_1_rd_en; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_in_bits_vec_1_imm; // @[Core.scala 42:25]
  wire  stall_reg_io_in_bits_vec_1_pred_br; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_in_bits_vec_1_pred_bpc; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_in_bits_vec_1_rs1_paddr; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_in_bits_vec_1_rs2_paddr; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_in_bits_vec_1_rd_paddr; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_in_bits_vec_1_rd_ppaddr; // @[Core.scala 42:25]
  wire  stall_reg_io_out_ready; // @[Core.scala 42:25]
  wire  stall_reg_io_out_valid; // @[Core.scala 42:25]
  wire  stall_reg_io_out_bits_vec_0_valid; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_out_bits_vec_0_pc; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_out_bits_vec_0_npc; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_out_bits_vec_0_inst; // @[Core.scala 42:25]
  wire [2:0] stall_reg_io_out_bits_vec_0_fu_code; // @[Core.scala 42:25]
  wire [3:0] stall_reg_io_out_bits_vec_0_alu_code; // @[Core.scala 42:25]
  wire [3:0] stall_reg_io_out_bits_vec_0_jmp_code; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_out_bits_vec_0_mem_code; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_out_bits_vec_0_mem_size; // @[Core.scala 42:25]
  wire [2:0] stall_reg_io_out_bits_vec_0_sys_code; // @[Core.scala 42:25]
  wire  stall_reg_io_out_bits_vec_0_w_type; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_out_bits_vec_0_rs1_src; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_out_bits_vec_0_rs2_src; // @[Core.scala 42:25]
  wire [4:0] stall_reg_io_out_bits_vec_0_rd_addr; // @[Core.scala 42:25]
  wire  stall_reg_io_out_bits_vec_0_rd_en; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_out_bits_vec_0_imm; // @[Core.scala 42:25]
  wire  stall_reg_io_out_bits_vec_0_pred_br; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_out_bits_vec_0_pred_bpc; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_out_bits_vec_0_rs1_paddr; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_out_bits_vec_0_rs2_paddr; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_out_bits_vec_0_rd_paddr; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_out_bits_vec_0_rd_ppaddr; // @[Core.scala 42:25]
  wire  stall_reg_io_out_bits_vec_1_valid; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_out_bits_vec_1_pc; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_out_bits_vec_1_npc; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_out_bits_vec_1_inst; // @[Core.scala 42:25]
  wire [2:0] stall_reg_io_out_bits_vec_1_fu_code; // @[Core.scala 42:25]
  wire [3:0] stall_reg_io_out_bits_vec_1_alu_code; // @[Core.scala 42:25]
  wire [3:0] stall_reg_io_out_bits_vec_1_jmp_code; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_out_bits_vec_1_mem_code; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_out_bits_vec_1_mem_size; // @[Core.scala 42:25]
  wire [2:0] stall_reg_io_out_bits_vec_1_sys_code; // @[Core.scala 42:25]
  wire  stall_reg_io_out_bits_vec_1_w_type; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_out_bits_vec_1_rs1_src; // @[Core.scala 42:25]
  wire [1:0] stall_reg_io_out_bits_vec_1_rs2_src; // @[Core.scala 42:25]
  wire [4:0] stall_reg_io_out_bits_vec_1_rd_addr; // @[Core.scala 42:25]
  wire  stall_reg_io_out_bits_vec_1_rd_en; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_out_bits_vec_1_imm; // @[Core.scala 42:25]
  wire  stall_reg_io_out_bits_vec_1_pred_br; // @[Core.scala 42:25]
  wire [31:0] stall_reg_io_out_bits_vec_1_pred_bpc; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_out_bits_vec_1_rs1_paddr; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_out_bits_vec_1_rs2_paddr; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_out_bits_vec_1_rd_paddr; // @[Core.scala 42:25]
  wire [5:0] stall_reg_io_out_bits_vec_1_rd_ppaddr; // @[Core.scala 42:25]
  wire  rob_clock; // @[Core.scala 46:19]
  wire  rob_reset; // @[Core.scala 46:19]
  wire  rob_io_in_ready; // @[Core.scala 46:19]
  wire  rob_io_in_valid; // @[Core.scala 46:19]
  wire  rob_io_in_bits_vec_0_valid; // @[Core.scala 46:19]
  wire [31:0] rob_io_in_bits_vec_0_pc; // @[Core.scala 46:19]
  wire [2:0] rob_io_in_bits_vec_0_fu_code; // @[Core.scala 46:19]
  wire [2:0] rob_io_in_bits_vec_0_sys_code; // @[Core.scala 46:19]
  wire [4:0] rob_io_in_bits_vec_0_rd_addr; // @[Core.scala 46:19]
  wire  rob_io_in_bits_vec_0_rd_en; // @[Core.scala 46:19]
  wire [5:0] rob_io_in_bits_vec_0_rd_paddr; // @[Core.scala 46:19]
  wire [5:0] rob_io_in_bits_vec_0_rd_ppaddr; // @[Core.scala 46:19]
  wire  rob_io_in_bits_vec_1_valid; // @[Core.scala 46:19]
  wire [31:0] rob_io_in_bits_vec_1_pc; // @[Core.scala 46:19]
  wire [2:0] rob_io_in_bits_vec_1_fu_code; // @[Core.scala 46:19]
  wire [2:0] rob_io_in_bits_vec_1_sys_code; // @[Core.scala 46:19]
  wire [4:0] rob_io_in_bits_vec_1_rd_addr; // @[Core.scala 46:19]
  wire  rob_io_in_bits_vec_1_rd_en; // @[Core.scala 46:19]
  wire [5:0] rob_io_in_bits_vec_1_rd_paddr; // @[Core.scala 46:19]
  wire [5:0] rob_io_in_bits_vec_1_rd_ppaddr; // @[Core.scala 46:19]
  wire [3:0] rob_io_rob_addr_0; // @[Core.scala 46:19]
  wire [3:0] rob_io_rob_addr_1; // @[Core.scala 46:19]
  wire  rob_io_exe_0_valid; // @[Core.scala 46:19]
  wire [3:0] rob_io_exe_0_rob_addr; // @[Core.scala 46:19]
  wire  rob_io_exe_1_valid; // @[Core.scala 46:19]
  wire [3:0] rob_io_exe_1_rob_addr; // @[Core.scala 46:19]
  wire  rob_io_exe_2_valid; // @[Core.scala 46:19]
  wire [3:0] rob_io_exe_2_rob_addr; // @[Core.scala 46:19]
  wire  rob_io_exe_ecp_0_jmp_valid; // @[Core.scala 46:19]
  wire  rob_io_exe_ecp_0_jmp; // @[Core.scala 46:19]
  wire [31:0] rob_io_exe_ecp_0_jmp_pc; // @[Core.scala 46:19]
  wire  rob_io_exe_ecp_0_mis; // @[Core.scala 46:19]
  wire  rob_io_exe_ecp_1_jmp_valid; // @[Core.scala 46:19]
  wire  rob_io_exe_ecp_1_jmp; // @[Core.scala 46:19]
  wire [31:0] rob_io_exe_ecp_1_jmp_pc; // @[Core.scala 46:19]
  wire  rob_io_exe_ecp_1_mis; // @[Core.scala 46:19]
  wire  rob_io_exe_ecp_2_store_valid; // @[Core.scala 46:19]
  wire  rob_io_cm_0_valid; // @[Core.scala 46:19]
  wire [4:0] rob_io_cm_0_rd_addr; // @[Core.scala 46:19]
  wire  rob_io_cm_0_rd_en; // @[Core.scala 46:19]
  wire [5:0] rob_io_cm_0_rd_paddr; // @[Core.scala 46:19]
  wire [5:0] rob_io_cm_0_rd_ppaddr; // @[Core.scala 46:19]
  wire  rob_io_cm_1_valid; // @[Core.scala 46:19]
  wire [4:0] rob_io_cm_1_rd_addr; // @[Core.scala 46:19]
  wire  rob_io_cm_1_rd_en; // @[Core.scala 46:19]
  wire [5:0] rob_io_cm_1_rd_paddr; // @[Core.scala 46:19]
  wire [5:0] rob_io_cm_1_rd_ppaddr; // @[Core.scala 46:19]
  wire  rob_io_jmp_packet_valid; // @[Core.scala 46:19]
  wire [31:0] rob_io_jmp_packet_inst_pc; // @[Core.scala 46:19]
  wire  rob_io_jmp_packet_jmp; // @[Core.scala 46:19]
  wire [31:0] rob_io_jmp_packet_jmp_pc; // @[Core.scala 46:19]
  wire  rob_io_jmp_packet_mis; // @[Core.scala 46:19]
  wire  rob_io_jmp_packet_sys; // @[Core.scala 46:19]
  wire  rob_io_sq_deq_req; // @[Core.scala 46:19]
  wire  rob_io_flush; // @[Core.scala 46:19]
  wire  rob_io_sys_ready; // @[Core.scala 46:19]
  wire  rob_csr_mip_mtip_intr_0; // @[Core.scala 46:19]
  wire [63:0] rob_intr_mcause_0; // @[Core.scala 46:19]
  wire [63:0] rob_intr_mstatus_0; // @[Core.scala 46:19]
  wire [29:0] rob_csr_mtvec_idx_0; // @[Core.scala 46:19]
  wire  rob_csr_mie_mtie_0; // @[Core.scala 46:19]
  wire  rob_intr_0; // @[Core.scala 46:19]
  wire [63:0] rob_csr_mstatus_0; // @[Core.scala 46:19]
  wire [63:0] rob_intr_mepc_0; // @[Core.scala 46:19]
  wire  isu_clock; // @[Core.scala 47:19]
  wire  isu_reset; // @[Core.scala 47:19]
  wire  isu_io_flush; // @[Core.scala 47:19]
  wire  isu_io_in_ready; // @[Core.scala 47:19]
  wire  isu_io_in_valid; // @[Core.scala 47:19]
  wire  isu_io_in_bits_vec_0_valid; // @[Core.scala 47:19]
  wire [31:0] isu_io_in_bits_vec_0_pc; // @[Core.scala 47:19]
  wire [31:0] isu_io_in_bits_vec_0_npc; // @[Core.scala 47:19]
  wire [31:0] isu_io_in_bits_vec_0_inst; // @[Core.scala 47:19]
  wire [2:0] isu_io_in_bits_vec_0_fu_code; // @[Core.scala 47:19]
  wire [3:0] isu_io_in_bits_vec_0_alu_code; // @[Core.scala 47:19]
  wire [3:0] isu_io_in_bits_vec_0_jmp_code; // @[Core.scala 47:19]
  wire [1:0] isu_io_in_bits_vec_0_mem_code; // @[Core.scala 47:19]
  wire [1:0] isu_io_in_bits_vec_0_mem_size; // @[Core.scala 47:19]
  wire [2:0] isu_io_in_bits_vec_0_sys_code; // @[Core.scala 47:19]
  wire  isu_io_in_bits_vec_0_w_type; // @[Core.scala 47:19]
  wire [1:0] isu_io_in_bits_vec_0_rs1_src; // @[Core.scala 47:19]
  wire [1:0] isu_io_in_bits_vec_0_rs2_src; // @[Core.scala 47:19]
  wire  isu_io_in_bits_vec_0_rd_en; // @[Core.scala 47:19]
  wire [31:0] isu_io_in_bits_vec_0_imm; // @[Core.scala 47:19]
  wire  isu_io_in_bits_vec_0_pred_br; // @[Core.scala 47:19]
  wire [31:0] isu_io_in_bits_vec_0_pred_bpc; // @[Core.scala 47:19]
  wire [5:0] isu_io_in_bits_vec_0_rs1_paddr; // @[Core.scala 47:19]
  wire [5:0] isu_io_in_bits_vec_0_rs2_paddr; // @[Core.scala 47:19]
  wire [5:0] isu_io_in_bits_vec_0_rd_paddr; // @[Core.scala 47:19]
  wire  isu_io_in_bits_vec_1_valid; // @[Core.scala 47:19]
  wire [31:0] isu_io_in_bits_vec_1_pc; // @[Core.scala 47:19]
  wire [31:0] isu_io_in_bits_vec_1_npc; // @[Core.scala 47:19]
  wire [31:0] isu_io_in_bits_vec_1_inst; // @[Core.scala 47:19]
  wire [2:0] isu_io_in_bits_vec_1_fu_code; // @[Core.scala 47:19]
  wire [3:0] isu_io_in_bits_vec_1_alu_code; // @[Core.scala 47:19]
  wire [3:0] isu_io_in_bits_vec_1_jmp_code; // @[Core.scala 47:19]
  wire [1:0] isu_io_in_bits_vec_1_mem_code; // @[Core.scala 47:19]
  wire [1:0] isu_io_in_bits_vec_1_mem_size; // @[Core.scala 47:19]
  wire [2:0] isu_io_in_bits_vec_1_sys_code; // @[Core.scala 47:19]
  wire  isu_io_in_bits_vec_1_w_type; // @[Core.scala 47:19]
  wire [1:0] isu_io_in_bits_vec_1_rs1_src; // @[Core.scala 47:19]
  wire [1:0] isu_io_in_bits_vec_1_rs2_src; // @[Core.scala 47:19]
  wire  isu_io_in_bits_vec_1_rd_en; // @[Core.scala 47:19]
  wire [31:0] isu_io_in_bits_vec_1_imm; // @[Core.scala 47:19]
  wire  isu_io_in_bits_vec_1_pred_br; // @[Core.scala 47:19]
  wire [31:0] isu_io_in_bits_vec_1_pred_bpc; // @[Core.scala 47:19]
  wire [5:0] isu_io_in_bits_vec_1_rs1_paddr; // @[Core.scala 47:19]
  wire [5:0] isu_io_in_bits_vec_1_rs2_paddr; // @[Core.scala 47:19]
  wire [5:0] isu_io_in_bits_vec_1_rd_paddr; // @[Core.scala 47:19]
  wire [3:0] isu_io_rob_addr_0; // @[Core.scala 47:19]
  wire [3:0] isu_io_rob_addr_1; // @[Core.scala 47:19]
  wire  isu_io_out_0_valid; // @[Core.scala 47:19]
  wire [31:0] isu_io_out_0_pc; // @[Core.scala 47:19]
  wire [31:0] isu_io_out_0_npc; // @[Core.scala 47:19]
  wire [31:0] isu_io_out_0_inst; // @[Core.scala 47:19]
  wire [2:0] isu_io_out_0_fu_code; // @[Core.scala 47:19]
  wire [3:0] isu_io_out_0_alu_code; // @[Core.scala 47:19]
  wire [3:0] isu_io_out_0_jmp_code; // @[Core.scala 47:19]
  wire [2:0] isu_io_out_0_sys_code; // @[Core.scala 47:19]
  wire  isu_io_out_0_w_type; // @[Core.scala 47:19]
  wire [1:0] isu_io_out_0_rs1_src; // @[Core.scala 47:19]
  wire [1:0] isu_io_out_0_rs2_src; // @[Core.scala 47:19]
  wire  isu_io_out_0_rd_en; // @[Core.scala 47:19]
  wire [31:0] isu_io_out_0_imm; // @[Core.scala 47:19]
  wire  isu_io_out_0_pred_br; // @[Core.scala 47:19]
  wire [31:0] isu_io_out_0_pred_bpc; // @[Core.scala 47:19]
  wire [5:0] isu_io_out_0_rs1_paddr; // @[Core.scala 47:19]
  wire [5:0] isu_io_out_0_rs2_paddr; // @[Core.scala 47:19]
  wire [5:0] isu_io_out_0_rd_paddr; // @[Core.scala 47:19]
  wire [3:0] isu_io_out_0_rob_addr; // @[Core.scala 47:19]
  wire  isu_io_out_1_valid; // @[Core.scala 47:19]
  wire [31:0] isu_io_out_1_pc; // @[Core.scala 47:19]
  wire [31:0] isu_io_out_1_npc; // @[Core.scala 47:19]
  wire [2:0] isu_io_out_1_fu_code; // @[Core.scala 47:19]
  wire [3:0] isu_io_out_1_alu_code; // @[Core.scala 47:19]
  wire [3:0] isu_io_out_1_jmp_code; // @[Core.scala 47:19]
  wire  isu_io_out_1_w_type; // @[Core.scala 47:19]
  wire [1:0] isu_io_out_1_rs1_src; // @[Core.scala 47:19]
  wire [1:0] isu_io_out_1_rs2_src; // @[Core.scala 47:19]
  wire  isu_io_out_1_rd_en; // @[Core.scala 47:19]
  wire [31:0] isu_io_out_1_imm; // @[Core.scala 47:19]
  wire  isu_io_out_1_pred_br; // @[Core.scala 47:19]
  wire [31:0] isu_io_out_1_pred_bpc; // @[Core.scala 47:19]
  wire [5:0] isu_io_out_1_rs1_paddr; // @[Core.scala 47:19]
  wire [5:0] isu_io_out_1_rs2_paddr; // @[Core.scala 47:19]
  wire [5:0] isu_io_out_1_rd_paddr; // @[Core.scala 47:19]
  wire [3:0] isu_io_out_1_rob_addr; // @[Core.scala 47:19]
  wire  isu_io_out_2_valid; // @[Core.scala 47:19]
  wire [31:0] isu_io_out_2_pc; // @[Core.scala 47:19]
  wire [2:0] isu_io_out_2_fu_code; // @[Core.scala 47:19]
  wire [3:0] isu_io_out_2_alu_code; // @[Core.scala 47:19]
  wire [1:0] isu_io_out_2_mem_code; // @[Core.scala 47:19]
  wire [1:0] isu_io_out_2_mem_size; // @[Core.scala 47:19]
  wire  isu_io_out_2_w_type; // @[Core.scala 47:19]
  wire [1:0] isu_io_out_2_rs1_src; // @[Core.scala 47:19]
  wire [1:0] isu_io_out_2_rs2_src; // @[Core.scala 47:19]
  wire  isu_io_out_2_rd_en; // @[Core.scala 47:19]
  wire [31:0] isu_io_out_2_imm; // @[Core.scala 47:19]
  wire [5:0] isu_io_out_2_rs1_paddr; // @[Core.scala 47:19]
  wire [5:0] isu_io_out_2_rs2_paddr; // @[Core.scala 47:19]
  wire [5:0] isu_io_out_2_rd_paddr; // @[Core.scala 47:19]
  wire [3:0] isu_io_out_2_rob_addr; // @[Core.scala 47:19]
  wire [63:0] isu_io_avail_list; // @[Core.scala 47:19]
  wire  isu_io_lsu_ready; // @[Core.scala 47:19]
  wire  isu_io_sys_ready; // @[Core.scala 47:19]
  wire  rf_clock; // @[Core.scala 70:18]
  wire  rf_reset; // @[Core.scala 70:18]
  wire  rf_io_in_0_valid; // @[Core.scala 70:18]
  wire [31:0] rf_io_in_0_pc; // @[Core.scala 70:18]
  wire [31:0] rf_io_in_0_npc; // @[Core.scala 70:18]
  wire [31:0] rf_io_in_0_inst; // @[Core.scala 70:18]
  wire [2:0] rf_io_in_0_fu_code; // @[Core.scala 70:18]
  wire [3:0] rf_io_in_0_alu_code; // @[Core.scala 70:18]
  wire [3:0] rf_io_in_0_jmp_code; // @[Core.scala 70:18]
  wire [2:0] rf_io_in_0_sys_code; // @[Core.scala 70:18]
  wire  rf_io_in_0_w_type; // @[Core.scala 70:18]
  wire [1:0] rf_io_in_0_rs1_src; // @[Core.scala 70:18]
  wire [1:0] rf_io_in_0_rs2_src; // @[Core.scala 70:18]
  wire  rf_io_in_0_rd_en; // @[Core.scala 70:18]
  wire [31:0] rf_io_in_0_imm; // @[Core.scala 70:18]
  wire  rf_io_in_0_pred_br; // @[Core.scala 70:18]
  wire [31:0] rf_io_in_0_pred_bpc; // @[Core.scala 70:18]
  wire [5:0] rf_io_in_0_rs1_paddr; // @[Core.scala 70:18]
  wire [5:0] rf_io_in_0_rs2_paddr; // @[Core.scala 70:18]
  wire [5:0] rf_io_in_0_rd_paddr; // @[Core.scala 70:18]
  wire [3:0] rf_io_in_0_rob_addr; // @[Core.scala 70:18]
  wire  rf_io_in_1_valid; // @[Core.scala 70:18]
  wire [31:0] rf_io_in_1_pc; // @[Core.scala 70:18]
  wire [31:0] rf_io_in_1_npc; // @[Core.scala 70:18]
  wire [2:0] rf_io_in_1_fu_code; // @[Core.scala 70:18]
  wire [3:0] rf_io_in_1_alu_code; // @[Core.scala 70:18]
  wire [3:0] rf_io_in_1_jmp_code; // @[Core.scala 70:18]
  wire  rf_io_in_1_w_type; // @[Core.scala 70:18]
  wire [1:0] rf_io_in_1_rs1_src; // @[Core.scala 70:18]
  wire [1:0] rf_io_in_1_rs2_src; // @[Core.scala 70:18]
  wire  rf_io_in_1_rd_en; // @[Core.scala 70:18]
  wire [31:0] rf_io_in_1_imm; // @[Core.scala 70:18]
  wire  rf_io_in_1_pred_br; // @[Core.scala 70:18]
  wire [31:0] rf_io_in_1_pred_bpc; // @[Core.scala 70:18]
  wire [5:0] rf_io_in_1_rs1_paddr; // @[Core.scala 70:18]
  wire [5:0] rf_io_in_1_rs2_paddr; // @[Core.scala 70:18]
  wire [5:0] rf_io_in_1_rd_paddr; // @[Core.scala 70:18]
  wire [3:0] rf_io_in_1_rob_addr; // @[Core.scala 70:18]
  wire  rf_io_in_2_valid; // @[Core.scala 70:18]
  wire [31:0] rf_io_in_2_pc; // @[Core.scala 70:18]
  wire [2:0] rf_io_in_2_fu_code; // @[Core.scala 70:18]
  wire [3:0] rf_io_in_2_alu_code; // @[Core.scala 70:18]
  wire [1:0] rf_io_in_2_mem_code; // @[Core.scala 70:18]
  wire [1:0] rf_io_in_2_mem_size; // @[Core.scala 70:18]
  wire  rf_io_in_2_w_type; // @[Core.scala 70:18]
  wire [1:0] rf_io_in_2_rs1_src; // @[Core.scala 70:18]
  wire [1:0] rf_io_in_2_rs2_src; // @[Core.scala 70:18]
  wire  rf_io_in_2_rd_en; // @[Core.scala 70:18]
  wire [31:0] rf_io_in_2_imm; // @[Core.scala 70:18]
  wire [5:0] rf_io_in_2_rs1_paddr; // @[Core.scala 70:18]
  wire [5:0] rf_io_in_2_rs2_paddr; // @[Core.scala 70:18]
  wire [5:0] rf_io_in_2_rd_paddr; // @[Core.scala 70:18]
  wire [3:0] rf_io_in_2_rob_addr; // @[Core.scala 70:18]
  wire  rf_io_out_0_valid; // @[Core.scala 70:18]
  wire [31:0] rf_io_out_0_pc; // @[Core.scala 70:18]
  wire [31:0] rf_io_out_0_npc; // @[Core.scala 70:18]
  wire [31:0] rf_io_out_0_inst; // @[Core.scala 70:18]
  wire [2:0] rf_io_out_0_fu_code; // @[Core.scala 70:18]
  wire [3:0] rf_io_out_0_alu_code; // @[Core.scala 70:18]
  wire [3:0] rf_io_out_0_jmp_code; // @[Core.scala 70:18]
  wire [2:0] rf_io_out_0_sys_code; // @[Core.scala 70:18]
  wire  rf_io_out_0_w_type; // @[Core.scala 70:18]
  wire [1:0] rf_io_out_0_rs1_src; // @[Core.scala 70:18]
  wire [1:0] rf_io_out_0_rs2_src; // @[Core.scala 70:18]
  wire  rf_io_out_0_rd_en; // @[Core.scala 70:18]
  wire [31:0] rf_io_out_0_imm; // @[Core.scala 70:18]
  wire  rf_io_out_0_pred_br; // @[Core.scala 70:18]
  wire [31:0] rf_io_out_0_pred_bpc; // @[Core.scala 70:18]
  wire [5:0] rf_io_out_0_rd_paddr; // @[Core.scala 70:18]
  wire [3:0] rf_io_out_0_rob_addr; // @[Core.scala 70:18]
  wire  rf_io_out_1_valid; // @[Core.scala 70:18]
  wire [31:0] rf_io_out_1_pc; // @[Core.scala 70:18]
  wire [31:0] rf_io_out_1_npc; // @[Core.scala 70:18]
  wire [2:0] rf_io_out_1_fu_code; // @[Core.scala 70:18]
  wire [3:0] rf_io_out_1_alu_code; // @[Core.scala 70:18]
  wire [3:0] rf_io_out_1_jmp_code; // @[Core.scala 70:18]
  wire  rf_io_out_1_w_type; // @[Core.scala 70:18]
  wire [1:0] rf_io_out_1_rs1_src; // @[Core.scala 70:18]
  wire [1:0] rf_io_out_1_rs2_src; // @[Core.scala 70:18]
  wire  rf_io_out_1_rd_en; // @[Core.scala 70:18]
  wire [31:0] rf_io_out_1_imm; // @[Core.scala 70:18]
  wire  rf_io_out_1_pred_br; // @[Core.scala 70:18]
  wire [31:0] rf_io_out_1_pred_bpc; // @[Core.scala 70:18]
  wire [5:0] rf_io_out_1_rd_paddr; // @[Core.scala 70:18]
  wire [3:0] rf_io_out_1_rob_addr; // @[Core.scala 70:18]
  wire  rf_io_out_2_valid; // @[Core.scala 70:18]
  wire [31:0] rf_io_out_2_pc; // @[Core.scala 70:18]
  wire [2:0] rf_io_out_2_fu_code; // @[Core.scala 70:18]
  wire [3:0] rf_io_out_2_alu_code; // @[Core.scala 70:18]
  wire [1:0] rf_io_out_2_mem_code; // @[Core.scala 70:18]
  wire [1:0] rf_io_out_2_mem_size; // @[Core.scala 70:18]
  wire  rf_io_out_2_w_type; // @[Core.scala 70:18]
  wire [1:0] rf_io_out_2_rs1_src; // @[Core.scala 70:18]
  wire [1:0] rf_io_out_2_rs2_src; // @[Core.scala 70:18]
  wire  rf_io_out_2_rd_en; // @[Core.scala 70:18]
  wire [31:0] rf_io_out_2_imm; // @[Core.scala 70:18]
  wire [5:0] rf_io_out_2_rd_paddr; // @[Core.scala 70:18]
  wire [3:0] rf_io_out_2_rob_addr; // @[Core.scala 70:18]
  wire [63:0] rf_io_rs1_data_0; // @[Core.scala 70:18]
  wire [63:0] rf_io_rs1_data_1; // @[Core.scala 70:18]
  wire [63:0] rf_io_rs1_data_2; // @[Core.scala 70:18]
  wire [63:0] rf_io_rs2_data_0; // @[Core.scala 70:18]
  wire [63:0] rf_io_rs2_data_1; // @[Core.scala 70:18]
  wire [63:0] rf_io_rs2_data_2; // @[Core.scala 70:18]
  wire  rf_io_rd_en_0; // @[Core.scala 70:18]
  wire  rf_io_rd_en_1; // @[Core.scala 70:18]
  wire  rf_io_rd_en_2; // @[Core.scala 70:18]
  wire [5:0] rf_io_rd_paddr_0; // @[Core.scala 70:18]
  wire [5:0] rf_io_rd_paddr_1; // @[Core.scala 70:18]
  wire [5:0] rf_io_rd_paddr_2; // @[Core.scala 70:18]
  wire [63:0] rf_io_rd_data_0; // @[Core.scala 70:18]
  wire [63:0] rf_io_rd_data_1; // @[Core.scala 70:18]
  wire [63:0] rf_io_rd_data_2; // @[Core.scala 70:18]
  wire  rf_io_flush; // @[Core.scala 70:18]
  wire  execution_clock; // @[Core.scala 76:25]
  wire  execution_reset; // @[Core.scala 76:25]
  wire  execution_io_in_0_valid; // @[Core.scala 76:25]
  wire [31:0] execution_io_in_0_pc; // @[Core.scala 76:25]
  wire [31:0] execution_io_in_0_npc; // @[Core.scala 76:25]
  wire [31:0] execution_io_in_0_inst; // @[Core.scala 76:25]
  wire [2:0] execution_io_in_0_fu_code; // @[Core.scala 76:25]
  wire [3:0] execution_io_in_0_alu_code; // @[Core.scala 76:25]
  wire [3:0] execution_io_in_0_jmp_code; // @[Core.scala 76:25]
  wire [2:0] execution_io_in_0_sys_code; // @[Core.scala 76:25]
  wire  execution_io_in_0_w_type; // @[Core.scala 76:25]
  wire [1:0] execution_io_in_0_rs1_src; // @[Core.scala 76:25]
  wire [1:0] execution_io_in_0_rs2_src; // @[Core.scala 76:25]
  wire  execution_io_in_0_rd_en; // @[Core.scala 76:25]
  wire [31:0] execution_io_in_0_imm; // @[Core.scala 76:25]
  wire  execution_io_in_0_pred_br; // @[Core.scala 76:25]
  wire [31:0] execution_io_in_0_pred_bpc; // @[Core.scala 76:25]
  wire [5:0] execution_io_in_0_rd_paddr; // @[Core.scala 76:25]
  wire [3:0] execution_io_in_0_rob_addr; // @[Core.scala 76:25]
  wire  execution_io_in_1_valid; // @[Core.scala 76:25]
  wire [31:0] execution_io_in_1_pc; // @[Core.scala 76:25]
  wire [31:0] execution_io_in_1_npc; // @[Core.scala 76:25]
  wire [2:0] execution_io_in_1_fu_code; // @[Core.scala 76:25]
  wire [3:0] execution_io_in_1_alu_code; // @[Core.scala 76:25]
  wire [3:0] execution_io_in_1_jmp_code; // @[Core.scala 76:25]
  wire  execution_io_in_1_w_type; // @[Core.scala 76:25]
  wire [1:0] execution_io_in_1_rs1_src; // @[Core.scala 76:25]
  wire [1:0] execution_io_in_1_rs2_src; // @[Core.scala 76:25]
  wire  execution_io_in_1_rd_en; // @[Core.scala 76:25]
  wire [31:0] execution_io_in_1_imm; // @[Core.scala 76:25]
  wire  execution_io_in_1_pred_br; // @[Core.scala 76:25]
  wire [31:0] execution_io_in_1_pred_bpc; // @[Core.scala 76:25]
  wire [5:0] execution_io_in_1_rd_paddr; // @[Core.scala 76:25]
  wire [3:0] execution_io_in_1_rob_addr; // @[Core.scala 76:25]
  wire  execution_io_in_2_valid; // @[Core.scala 76:25]
  wire [31:0] execution_io_in_2_pc; // @[Core.scala 76:25]
  wire [2:0] execution_io_in_2_fu_code; // @[Core.scala 76:25]
  wire [3:0] execution_io_in_2_alu_code; // @[Core.scala 76:25]
  wire [1:0] execution_io_in_2_mem_code; // @[Core.scala 76:25]
  wire [1:0] execution_io_in_2_mem_size; // @[Core.scala 76:25]
  wire  execution_io_in_2_w_type; // @[Core.scala 76:25]
  wire [1:0] execution_io_in_2_rs1_src; // @[Core.scala 76:25]
  wire [1:0] execution_io_in_2_rs2_src; // @[Core.scala 76:25]
  wire  execution_io_in_2_rd_en; // @[Core.scala 76:25]
  wire [31:0] execution_io_in_2_imm; // @[Core.scala 76:25]
  wire [5:0] execution_io_in_2_rd_paddr; // @[Core.scala 76:25]
  wire [3:0] execution_io_in_2_rob_addr; // @[Core.scala 76:25]
  wire [63:0] execution_io_rs1_data_0; // @[Core.scala 76:25]
  wire [63:0] execution_io_rs1_data_1; // @[Core.scala 76:25]
  wire [63:0] execution_io_rs1_data_2; // @[Core.scala 76:25]
  wire [63:0] execution_io_rs2_data_0; // @[Core.scala 76:25]
  wire [63:0] execution_io_rs2_data_1; // @[Core.scala 76:25]
  wire [63:0] execution_io_rs2_data_2; // @[Core.scala 76:25]
  wire  execution_io_out_0_valid; // @[Core.scala 76:25]
  wire [3:0] execution_io_out_0_rob_addr; // @[Core.scala 76:25]
  wire  execution_io_out_1_valid; // @[Core.scala 76:25]
  wire [3:0] execution_io_out_1_rob_addr; // @[Core.scala 76:25]
  wire  execution_io_out_2_valid; // @[Core.scala 76:25]
  wire [3:0] execution_io_out_2_rob_addr; // @[Core.scala 76:25]
  wire  execution_io_out_ecp_0_jmp_valid; // @[Core.scala 76:25]
  wire  execution_io_out_ecp_0_jmp; // @[Core.scala 76:25]
  wire [31:0] execution_io_out_ecp_0_jmp_pc; // @[Core.scala 76:25]
  wire  execution_io_out_ecp_0_mis; // @[Core.scala 76:25]
  wire  execution_io_out_ecp_1_jmp_valid; // @[Core.scala 76:25]
  wire  execution_io_out_ecp_1_jmp; // @[Core.scala 76:25]
  wire [31:0] execution_io_out_ecp_1_jmp_pc; // @[Core.scala 76:25]
  wire  execution_io_out_ecp_1_mis; // @[Core.scala 76:25]
  wire  execution_io_out_ecp_2_store_valid; // @[Core.scala 76:25]
  wire  execution_io_rd_en_0; // @[Core.scala 76:25]
  wire  execution_io_rd_en_1; // @[Core.scala 76:25]
  wire  execution_io_rd_en_2; // @[Core.scala 76:25]
  wire [5:0] execution_io_rd_paddr_0; // @[Core.scala 76:25]
  wire [5:0] execution_io_rd_paddr_1; // @[Core.scala 76:25]
  wire [5:0] execution_io_rd_paddr_2; // @[Core.scala 76:25]
  wire [63:0] execution_io_rd_data_0; // @[Core.scala 76:25]
  wire [63:0] execution_io_rd_data_1; // @[Core.scala 76:25]
  wire [63:0] execution_io_rd_data_2; // @[Core.scala 76:25]
  wire  execution_io_flush; // @[Core.scala 76:25]
  wire  execution_io_lsu_ready; // @[Core.scala 76:25]
  wire  execution_io_dmem_st_req_ready; // @[Core.scala 76:25]
  wire  execution_io_dmem_st_req_valid; // @[Core.scala 76:25]
  wire [31:0] execution_io_dmem_st_req_bits_addr; // @[Core.scala 76:25]
  wire [63:0] execution_io_dmem_st_req_bits_wdata; // @[Core.scala 76:25]
  wire [7:0] execution_io_dmem_st_req_bits_wmask; // @[Core.scala 76:25]
  wire [1:0] execution_io_dmem_st_req_bits_size; // @[Core.scala 76:25]
  wire  execution_io_dmem_st_resp_ready; // @[Core.scala 76:25]
  wire  execution_io_dmem_st_resp_valid; // @[Core.scala 76:25]
  wire  execution_io_dmem_ld_req_ready; // @[Core.scala 76:25]
  wire  execution_io_dmem_ld_req_valid; // @[Core.scala 76:25]
  wire [31:0] execution_io_dmem_ld_req_bits_addr; // @[Core.scala 76:25]
  wire [1:0] execution_io_dmem_ld_req_bits_size; // @[Core.scala 76:25]
  wire  execution_io_dmem_ld_resp_ready; // @[Core.scala 76:25]
  wire  execution_io_dmem_ld_resp_valid; // @[Core.scala 76:25]
  wire [63:0] execution_io_dmem_ld_resp_bits_rdata; // @[Core.scala 76:25]
  wire  execution_io_lsu_wakeup_uop_valid; // @[Core.scala 76:25]
  wire  execution_io_lsu_wakeup_uop_rd_en; // @[Core.scala 76:25]
  wire [5:0] execution_io_lsu_wakeup_uop_rd_paddr; // @[Core.scala 76:25]
  wire  execution_mtip; // @[Core.scala 76:25]
  wire [63:0] execution_intr_mcause; // @[Core.scala 76:25]
  wire [63:0] execution_instr_cnt; // @[Core.scala 76:25]
  wire [63:0] execution_intr_mstatus; // @[Core.scala 76:25]
  wire [29:0] execution__T_6_0; // @[Core.scala 76:25]
  wire  execution__T_5_0; // @[Core.scala 76:25]
  wire  execution_intr; // @[Core.scala 76:25]
  wire  execution_fence_i; // @[Core.scala 76:25]
  wire [63:0] execution_cycle_cnt; // @[Core.scala 76:25]
  wire [63:0] execution_mstatus; // @[Core.scala 76:25]
  wire [63:0] execution_intr_mepc; // @[Core.scala 76:25]
  wire  execution_mtip_0; // @[Core.scala 76:25]
  wire  sq_clock; // @[Core.scala 95:18]
  wire  sq_reset; // @[Core.scala 95:18]
  wire  sq_io_flush; // @[Core.scala 95:18]
  wire  sq_io_in_st_req_ready; // @[Core.scala 95:18]
  wire  sq_io_in_st_req_valid; // @[Core.scala 95:18]
  wire [31:0] sq_io_in_st_req_bits_addr; // @[Core.scala 95:18]
  wire [63:0] sq_io_in_st_req_bits_wdata; // @[Core.scala 95:18]
  wire [7:0] sq_io_in_st_req_bits_wmask; // @[Core.scala 95:18]
  wire [1:0] sq_io_in_st_req_bits_size; // @[Core.scala 95:18]
  wire  sq_io_in_st_resp_ready; // @[Core.scala 95:18]
  wire  sq_io_in_st_resp_valid; // @[Core.scala 95:18]
  wire  sq_io_in_ld_req_ready; // @[Core.scala 95:18]
  wire  sq_io_in_ld_req_valid; // @[Core.scala 95:18]
  wire [31:0] sq_io_in_ld_req_bits_addr; // @[Core.scala 95:18]
  wire [1:0] sq_io_in_ld_req_bits_size; // @[Core.scala 95:18]
  wire  sq_io_in_ld_resp_ready; // @[Core.scala 95:18]
  wire  sq_io_in_ld_resp_valid; // @[Core.scala 95:18]
  wire [63:0] sq_io_in_ld_resp_bits_rdata; // @[Core.scala 95:18]
  wire  sq_io_out_st_req_ready; // @[Core.scala 95:18]
  wire  sq_io_out_st_req_valid; // @[Core.scala 95:18]
  wire [31:0] sq_io_out_st_req_bits_addr; // @[Core.scala 95:18]
  wire [63:0] sq_io_out_st_req_bits_wdata; // @[Core.scala 95:18]
  wire [7:0] sq_io_out_st_req_bits_wmask; // @[Core.scala 95:18]
  wire [1:0] sq_io_out_st_req_bits_size; // @[Core.scala 95:18]
  wire  sq_io_out_st_resp_ready; // @[Core.scala 95:18]
  wire  sq_io_out_st_resp_valid; // @[Core.scala 95:18]
  wire  sq_io_out_ld_req_ready; // @[Core.scala 95:18]
  wire  sq_io_out_ld_req_valid; // @[Core.scala 95:18]
  wire [31:0] sq_io_out_ld_req_bits_addr; // @[Core.scala 95:18]
  wire [1:0] sq_io_out_ld_req_bits_size; // @[Core.scala 95:18]
  wire  sq_io_out_ld_resp_ready; // @[Core.scala 95:18]
  wire  sq_io_out_ld_resp_valid; // @[Core.scala 95:18]
  wire [63:0] sq_io_out_ld_resp_bits_rdata; // @[Core.scala 95:18]
  wire  sq_io_deq_req; // @[Core.scala 95:18]
  wire  sq_empty_0; // @[Core.scala 95:18]
  wire  crossbar2to1_clock; // @[Core.scala 101:28]
  wire  crossbar2to1_io_in_0_req_ready; // @[Core.scala 101:28]
  wire  crossbar2to1_io_in_0_req_valid; // @[Core.scala 101:28]
  wire [31:0] crossbar2to1_io_in_0_req_bits_addr; // @[Core.scala 101:28]
  wire [63:0] crossbar2to1_io_in_0_req_bits_wdata; // @[Core.scala 101:28]
  wire [7:0] crossbar2to1_io_in_0_req_bits_wmask; // @[Core.scala 101:28]
  wire [1:0] crossbar2to1_io_in_0_req_bits_size; // @[Core.scala 101:28]
  wire  crossbar2to1_io_in_0_resp_ready; // @[Core.scala 101:28]
  wire  crossbar2to1_io_in_0_resp_valid; // @[Core.scala 101:28]
  wire  crossbar2to1_io_in_1_req_ready; // @[Core.scala 101:28]
  wire  crossbar2to1_io_in_1_req_valid; // @[Core.scala 101:28]
  wire [31:0] crossbar2to1_io_in_1_req_bits_addr; // @[Core.scala 101:28]
  wire [1:0] crossbar2to1_io_in_1_req_bits_size; // @[Core.scala 101:28]
  wire  crossbar2to1_io_in_1_resp_ready; // @[Core.scala 101:28]
  wire  crossbar2to1_io_in_1_resp_valid; // @[Core.scala 101:28]
  wire [63:0] crossbar2to1_io_in_1_resp_bits_rdata; // @[Core.scala 101:28]
  wire  crossbar2to1_io_out_req_ready; // @[Core.scala 101:28]
  wire  crossbar2to1_io_out_req_valid; // @[Core.scala 101:28]
  wire [3:0] crossbar2to1_io_out_req_bits_id; // @[Core.scala 101:28]
  wire [31:0] crossbar2to1_io_out_req_bits_addr; // @[Core.scala 101:28]
  wire [63:0] crossbar2to1_io_out_req_bits_wdata; // @[Core.scala 101:28]
  wire [7:0] crossbar2to1_io_out_req_bits_wmask; // @[Core.scala 101:28]
  wire  crossbar2to1_io_out_req_bits_wen; // @[Core.scala 101:28]
  wire [1:0] crossbar2to1_io_out_req_bits_size; // @[Core.scala 101:28]
  wire  crossbar2to1_io_out_resp_ready; // @[Core.scala 101:28]
  wire  crossbar2to1_io_out_resp_valid; // @[Core.scala 101:28]
  wire [3:0] crossbar2to1_io_out_resp_bits_id; // @[Core.scala 101:28]
  wire [63:0] crossbar2to1_io_out_resp_bits_rdata; // @[Core.scala 101:28]
  wire  crossbar1to2_clock; // @[Core.scala 105:28]
  wire  crossbar1to2_reset; // @[Core.scala 105:28]
  wire  crossbar1to2_io_in_req_ready; // @[Core.scala 105:28]
  wire  crossbar1to2_io_in_req_valid; // @[Core.scala 105:28]
  wire [3:0] crossbar1to2_io_in_req_bits_id; // @[Core.scala 105:28]
  wire [31:0] crossbar1to2_io_in_req_bits_addr; // @[Core.scala 105:28]
  wire [63:0] crossbar1to2_io_in_req_bits_wdata; // @[Core.scala 105:28]
  wire [7:0] crossbar1to2_io_in_req_bits_wmask; // @[Core.scala 105:28]
  wire  crossbar1to2_io_in_req_bits_wen; // @[Core.scala 105:28]
  wire [1:0] crossbar1to2_io_in_req_bits_size; // @[Core.scala 105:28]
  wire  crossbar1to2_io_in_resp_ready; // @[Core.scala 105:28]
  wire  crossbar1to2_io_in_resp_valid; // @[Core.scala 105:28]
  wire [3:0] crossbar1to2_io_in_resp_bits_id; // @[Core.scala 105:28]
  wire [63:0] crossbar1to2_io_in_resp_bits_rdata; // @[Core.scala 105:28]
  wire  crossbar1to2_io_out_0_req_ready; // @[Core.scala 105:28]
  wire  crossbar1to2_io_out_0_req_valid; // @[Core.scala 105:28]
  wire [3:0] crossbar1to2_io_out_0_req_bits_id; // @[Core.scala 105:28]
  wire [31:0] crossbar1to2_io_out_0_req_bits_addr; // @[Core.scala 105:28]
  wire [63:0] crossbar1to2_io_out_0_req_bits_wdata; // @[Core.scala 105:28]
  wire [7:0] crossbar1to2_io_out_0_req_bits_wmask; // @[Core.scala 105:28]
  wire  crossbar1to2_io_out_0_req_bits_wen; // @[Core.scala 105:28]
  wire [1:0] crossbar1to2_io_out_0_req_bits_size; // @[Core.scala 105:28]
  wire  crossbar1to2_io_out_0_resp_ready; // @[Core.scala 105:28]
  wire  crossbar1to2_io_out_0_resp_valid; // @[Core.scala 105:28]
  wire [3:0] crossbar1to2_io_out_0_resp_bits_id; // @[Core.scala 105:28]
  wire [63:0] crossbar1to2_io_out_0_resp_bits_rdata; // @[Core.scala 105:28]
  wire  crossbar1to2_io_out_1_req_ready; // @[Core.scala 105:28]
  wire  crossbar1to2_io_out_1_req_valid; // @[Core.scala 105:28]
  wire [3:0] crossbar1to2_io_out_1_req_bits_id; // @[Core.scala 105:28]
  wire [31:0] crossbar1to2_io_out_1_req_bits_addr; // @[Core.scala 105:28]
  wire [63:0] crossbar1to2_io_out_1_req_bits_wdata; // @[Core.scala 105:28]
  wire [7:0] crossbar1to2_io_out_1_req_bits_wmask; // @[Core.scala 105:28]
  wire  crossbar1to2_io_out_1_req_bits_wen; // @[Core.scala 105:28]
  wire [1:0] crossbar1to2_io_out_1_req_bits_size; // @[Core.scala 105:28]
  wire  crossbar1to2_io_out_1_resp_ready; // @[Core.scala 105:28]
  wire  crossbar1to2_io_out_1_resp_valid; // @[Core.scala 105:28]
  wire [3:0] crossbar1to2_io_out_1_resp_bits_id; // @[Core.scala 105:28]
  wire [63:0] crossbar1to2_io_out_1_resp_bits_rdata; // @[Core.scala 105:28]
  wire  crossbar1to2_io_to_1; // @[Core.scala 105:28]
  wire  dcache_clock; // @[Core.scala 112:22]
  wire  dcache_reset; // @[Core.scala 112:22]
  wire  dcache_io_in_req_ready; // @[Core.scala 112:22]
  wire  dcache_io_in_req_valid; // @[Core.scala 112:22]
  wire [3:0] dcache_io_in_req_bits_id; // @[Core.scala 112:22]
  wire [31:0] dcache_io_in_req_bits_addr; // @[Core.scala 112:22]
  wire [63:0] dcache_io_in_req_bits_wdata; // @[Core.scala 112:22]
  wire [7:0] dcache_io_in_req_bits_wmask; // @[Core.scala 112:22]
  wire  dcache_io_in_req_bits_wen; // @[Core.scala 112:22]
  wire [1:0] dcache_io_in_req_bits_size; // @[Core.scala 112:22]
  wire  dcache_io_in_resp_ready; // @[Core.scala 112:22]
  wire  dcache_io_in_resp_valid; // @[Core.scala 112:22]
  wire [3:0] dcache_io_in_resp_bits_id; // @[Core.scala 112:22]
  wire [63:0] dcache_io_in_resp_bits_rdata; // @[Core.scala 112:22]
  wire  dcache_io_out_cache_req_ready; // @[Core.scala 112:22]
  wire  dcache_io_out_cache_req_valid; // @[Core.scala 112:22]
  wire [31:0] dcache_io_out_cache_req_bits_addr; // @[Core.scala 112:22]
  wire  dcache_io_out_cache_req_bits_aen; // @[Core.scala 112:22]
  wire [63:0] dcache_io_out_cache_req_bits_wdata; // @[Core.scala 112:22]
  wire  dcache_io_out_cache_req_bits_wlast; // @[Core.scala 112:22]
  wire  dcache_io_out_cache_req_bits_wen; // @[Core.scala 112:22]
  wire  dcache_io_out_cache_resp_ready; // @[Core.scala 112:22]
  wire  dcache_io_out_cache_resp_valid; // @[Core.scala 112:22]
  wire [63:0] dcache_io_out_cache_resp_bits_rdata; // @[Core.scala 112:22]
  wire  dcache_io_out_cache_resp_bits_rlast; // @[Core.scala 112:22]
  wire  dcache_io_out_uncache_req_ready; // @[Core.scala 112:22]
  wire  dcache_io_out_uncache_req_valid; // @[Core.scala 112:22]
  wire [31:0] dcache_io_out_uncache_req_bits_addr; // @[Core.scala 112:22]
  wire [63:0] dcache_io_out_uncache_req_bits_wdata; // @[Core.scala 112:22]
  wire [7:0] dcache_io_out_uncache_req_bits_wmask; // @[Core.scala 112:22]
  wire  dcache_io_out_uncache_req_bits_wen; // @[Core.scala 112:22]
  wire [1:0] dcache_io_out_uncache_req_bits_size; // @[Core.scala 112:22]
  wire  dcache_io_out_uncache_resp_ready; // @[Core.scala 112:22]
  wire  dcache_io_out_uncache_resp_valid; // @[Core.scala 112:22]
  wire [63:0] dcache_io_out_uncache_resp_bits_rdata; // @[Core.scala 112:22]
  wire  dcache_fence_i; // @[Core.scala 112:22]
  wire  dcache__WIRE_10; // @[Core.scala 112:22]
  wire  dcache_empty; // @[Core.scala 112:22]
  wire  clint_clock; // @[Core.scala 117:21]
  wire  clint_reset; // @[Core.scala 117:21]
  wire  clint_io_in_req_ready; // @[Core.scala 117:21]
  wire  clint_io_in_req_valid; // @[Core.scala 117:21]
  wire [3:0] clint_io_in_req_bits_id; // @[Core.scala 117:21]
  wire [31:0] clint_io_in_req_bits_addr; // @[Core.scala 117:21]
  wire [63:0] clint_io_in_req_bits_wdata; // @[Core.scala 117:21]
  wire [7:0] clint_io_in_req_bits_wmask; // @[Core.scala 117:21]
  wire  clint_io_in_req_bits_wen; // @[Core.scala 117:21]
  wire  clint_io_in_resp_ready; // @[Core.scala 117:21]
  wire  clint_io_in_resp_valid; // @[Core.scala 117:21]
  wire [3:0] clint_io_in_resp_bits_id; // @[Core.scala 117:21]
  wire [63:0] clint_io_in_resp_bits_rdata; // @[Core.scala 117:21]
  wire  clint_mtip_1; // @[Core.scala 117:21]
  reg  REG; // @[Core.scala 53:34]
  reg [63:0] cycle_cnt; // @[Core.scala 132:26]
  reg [63:0] instr_cnt; // @[Core.scala 133:26]
  wire [63:0] _T_8 = cycle_cnt + 64'h1; // @[Core.scala 138:26]
  wire [1:0] _T_9 = rob_io_cm_0_valid + rob_io_cm_1_valid; // @[Bitwise.scala 47:55]
  wire [63:0] _GEN_0 = {{62'd0}, _T_9}; // @[Core.scala 139:26]
  wire [63:0] _T_12 = instr_cnt + _GEN_0; // @[Core.scala 139:26]
  ysyx_210128_InstFetch fetch ( // @[Core.scala 17:21]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_imem_req_ready(fetch_io_imem_req_ready),
    .io_imem_req_valid(fetch_io_imem_req_valid),
    .io_imem_req_bits_addr(fetch_io_imem_req_bits_addr),
    .io_imem_req_bits_user(fetch_io_imem_req_bits_user),
    .io_imem_resp_ready(fetch_io_imem_resp_ready),
    .io_imem_resp_valid(fetch_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(fetch_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(fetch_io_imem_resp_bits_user),
    .io_jmp_packet_valid(fetch_io_jmp_packet_valid),
    .io_jmp_packet_inst_pc(fetch_io_jmp_packet_inst_pc),
    .io_jmp_packet_jmp(fetch_io_jmp_packet_jmp),
    .io_jmp_packet_jmp_pc(fetch_io_jmp_packet_jmp_pc),
    .io_jmp_packet_mis(fetch_io_jmp_packet_mis),
    .io_jmp_packet_sys(fetch_io_jmp_packet_sys),
    .io_out_ready(fetch_io_out_ready),
    .io_out_valid(fetch_io_out_valid),
    .io_out_bits_vec_0_pc(fetch_io_out_bits_vec_0_pc),
    .io_out_bits_vec_0_inst(fetch_io_out_bits_vec_0_inst),
    .io_out_bits_vec_0_pred_br(fetch_io_out_bits_vec_0_pred_br),
    .io_out_bits_vec_0_pred_bpc(fetch_io_out_bits_vec_0_pred_bpc),
    .io_out_bits_vec_0_valid(fetch_io_out_bits_vec_0_valid),
    .io_out_bits_vec_1_pc(fetch_io_out_bits_vec_1_pc),
    .io_out_bits_vec_1_inst(fetch_io_out_bits_vec_1_inst),
    .io_out_bits_vec_1_pred_br(fetch_io_out_bits_vec_1_pred_br),
    .io_out_bits_vec_1_pred_bpc(fetch_io_out_bits_vec_1_pred_bpc),
    .io_out_bits_vec_1_valid(fetch_io_out_bits_vec_1_valid)
  );
  ysyx_210128_CacheController icache ( // @[Core.scala 19:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_in_req_ready(icache_io_in_req_ready),
    .io_in_req_valid(icache_io_in_req_valid),
    .io_in_req_bits_addr(icache_io_in_req_bits_addr),
    .io_in_req_bits_user(icache_io_in_req_bits_user),
    .io_in_resp_ready(icache_io_in_resp_ready),
    .io_in_resp_valid(icache_io_in_resp_valid),
    .io_in_resp_bits_rdata(icache_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(icache_io_in_resp_bits_user),
    .io_out_cache_req_ready(icache_io_out_cache_req_ready),
    .io_out_cache_req_valid(icache_io_out_cache_req_valid),
    .io_out_cache_req_bits_addr(icache_io_out_cache_req_bits_addr),
    .io_out_cache_req_bits_aen(icache_io_out_cache_req_bits_aen),
    .io_out_cache_req_bits_wdata(icache_io_out_cache_req_bits_wdata),
    .io_out_cache_req_bits_wlast(icache_io_out_cache_req_bits_wlast),
    .io_out_cache_req_bits_wen(icache_io_out_cache_req_bits_wen),
    .io_out_cache_resp_ready(icache_io_out_cache_resp_ready),
    .io_out_cache_resp_valid(icache_io_out_cache_resp_valid),
    .io_out_cache_resp_bits_rdata(icache_io_out_cache_resp_bits_rdata),
    .io_out_cache_resp_bits_rlast(icache_io_out_cache_resp_bits_rlast),
    .io_out_uncache_req_ready(icache_io_out_uncache_req_ready),
    .io_out_uncache_req_valid(icache_io_out_uncache_req_valid),
    .io_out_uncache_req_bits_addr(icache_io_out_uncache_req_bits_addr),
    .io_out_uncache_req_bits_size(icache_io_out_uncache_req_bits_size),
    .io_out_uncache_resp_ready(icache_io_out_uncache_resp_ready),
    .io_out_uncache_resp_valid(icache_io_out_uncache_resp_valid),
    .io_out_uncache_resp_bits_rdata(icache_io_out_uncache_resp_bits_rdata),
    .fence_i(icache_fence_i),
    ._WIRE_10(icache__WIRE_10),
    .empty(icache_empty)
  );
  ysyx_210128_InstBuffer ibuf ( // @[Core.scala 26:20]
    .clock(ibuf_clock),
    .reset(ibuf_reset),
    .io_in_ready(ibuf_io_in_ready),
    .io_in_valid(ibuf_io_in_valid),
    .io_in_bits_vec_0_pc(ibuf_io_in_bits_vec_0_pc),
    .io_in_bits_vec_0_inst(ibuf_io_in_bits_vec_0_inst),
    .io_in_bits_vec_0_pred_br(ibuf_io_in_bits_vec_0_pred_br),
    .io_in_bits_vec_0_pred_bpc(ibuf_io_in_bits_vec_0_pred_bpc),
    .io_in_bits_vec_0_valid(ibuf_io_in_bits_vec_0_valid),
    .io_in_bits_vec_1_pc(ibuf_io_in_bits_vec_1_pc),
    .io_in_bits_vec_1_inst(ibuf_io_in_bits_vec_1_inst),
    .io_in_bits_vec_1_pred_br(ibuf_io_in_bits_vec_1_pred_br),
    .io_in_bits_vec_1_pred_bpc(ibuf_io_in_bits_vec_1_pred_bpc),
    .io_in_bits_vec_1_valid(ibuf_io_in_bits_vec_1_valid),
    .io_out_ready(ibuf_io_out_ready),
    .io_out_valid(ibuf_io_out_valid),
    .io_out_bits_vec_0_pc(ibuf_io_out_bits_vec_0_pc),
    .io_out_bits_vec_0_inst(ibuf_io_out_bits_vec_0_inst),
    .io_out_bits_vec_0_pred_br(ibuf_io_out_bits_vec_0_pred_br),
    .io_out_bits_vec_0_pred_bpc(ibuf_io_out_bits_vec_0_pred_bpc),
    .io_out_bits_vec_0_valid(ibuf_io_out_bits_vec_0_valid),
    .io_out_bits_vec_1_pc(ibuf_io_out_bits_vec_1_pc),
    .io_out_bits_vec_1_inst(ibuf_io_out_bits_vec_1_inst),
    .io_out_bits_vec_1_pred_br(ibuf_io_out_bits_vec_1_pred_br),
    .io_out_bits_vec_1_pred_bpc(ibuf_io_out_bits_vec_1_pred_bpc),
    .io_out_bits_vec_1_valid(ibuf_io_out_bits_vec_1_valid),
    .io_flush(ibuf_io_flush)
  );
  ysyx_210128_Decode decode ( // @[Core.scala 32:22]
    .clock(decode_clock),
    .reset(decode_reset),
    .io_in_ready(decode_io_in_ready),
    .io_in_valid(decode_io_in_valid),
    .io_in_bits_vec_0_pc(decode_io_in_bits_vec_0_pc),
    .io_in_bits_vec_0_inst(decode_io_in_bits_vec_0_inst),
    .io_in_bits_vec_0_pred_br(decode_io_in_bits_vec_0_pred_br),
    .io_in_bits_vec_0_pred_bpc(decode_io_in_bits_vec_0_pred_bpc),
    .io_in_bits_vec_0_valid(decode_io_in_bits_vec_0_valid),
    .io_in_bits_vec_1_pc(decode_io_in_bits_vec_1_pc),
    .io_in_bits_vec_1_inst(decode_io_in_bits_vec_1_inst),
    .io_in_bits_vec_1_pred_br(decode_io_in_bits_vec_1_pred_br),
    .io_in_bits_vec_1_pred_bpc(decode_io_in_bits_vec_1_pred_bpc),
    .io_in_bits_vec_1_valid(decode_io_in_bits_vec_1_valid),
    .io_out_ready(decode_io_out_ready),
    .io_out_valid(decode_io_out_valid),
    .io_out_bits_vec_0_valid(decode_io_out_bits_vec_0_valid),
    .io_out_bits_vec_0_pc(decode_io_out_bits_vec_0_pc),
    .io_out_bits_vec_0_npc(decode_io_out_bits_vec_0_npc),
    .io_out_bits_vec_0_inst(decode_io_out_bits_vec_0_inst),
    .io_out_bits_vec_0_fu_code(decode_io_out_bits_vec_0_fu_code),
    .io_out_bits_vec_0_alu_code(decode_io_out_bits_vec_0_alu_code),
    .io_out_bits_vec_0_jmp_code(decode_io_out_bits_vec_0_jmp_code),
    .io_out_bits_vec_0_mem_code(decode_io_out_bits_vec_0_mem_code),
    .io_out_bits_vec_0_mem_size(decode_io_out_bits_vec_0_mem_size),
    .io_out_bits_vec_0_sys_code(decode_io_out_bits_vec_0_sys_code),
    .io_out_bits_vec_0_w_type(decode_io_out_bits_vec_0_w_type),
    .io_out_bits_vec_0_rs1_src(decode_io_out_bits_vec_0_rs1_src),
    .io_out_bits_vec_0_rs2_src(decode_io_out_bits_vec_0_rs2_src),
    .io_out_bits_vec_0_rs1_addr(decode_io_out_bits_vec_0_rs1_addr),
    .io_out_bits_vec_0_rs2_addr(decode_io_out_bits_vec_0_rs2_addr),
    .io_out_bits_vec_0_rd_addr(decode_io_out_bits_vec_0_rd_addr),
    .io_out_bits_vec_0_rd_en(decode_io_out_bits_vec_0_rd_en),
    .io_out_bits_vec_0_imm(decode_io_out_bits_vec_0_imm),
    .io_out_bits_vec_0_pred_br(decode_io_out_bits_vec_0_pred_br),
    .io_out_bits_vec_0_pred_bpc(decode_io_out_bits_vec_0_pred_bpc),
    .io_out_bits_vec_1_valid(decode_io_out_bits_vec_1_valid),
    .io_out_bits_vec_1_pc(decode_io_out_bits_vec_1_pc),
    .io_out_bits_vec_1_npc(decode_io_out_bits_vec_1_npc),
    .io_out_bits_vec_1_inst(decode_io_out_bits_vec_1_inst),
    .io_out_bits_vec_1_fu_code(decode_io_out_bits_vec_1_fu_code),
    .io_out_bits_vec_1_alu_code(decode_io_out_bits_vec_1_alu_code),
    .io_out_bits_vec_1_jmp_code(decode_io_out_bits_vec_1_jmp_code),
    .io_out_bits_vec_1_mem_code(decode_io_out_bits_vec_1_mem_code),
    .io_out_bits_vec_1_mem_size(decode_io_out_bits_vec_1_mem_size),
    .io_out_bits_vec_1_sys_code(decode_io_out_bits_vec_1_sys_code),
    .io_out_bits_vec_1_w_type(decode_io_out_bits_vec_1_w_type),
    .io_out_bits_vec_1_rs1_src(decode_io_out_bits_vec_1_rs1_src),
    .io_out_bits_vec_1_rs2_src(decode_io_out_bits_vec_1_rs2_src),
    .io_out_bits_vec_1_rs1_addr(decode_io_out_bits_vec_1_rs1_addr),
    .io_out_bits_vec_1_rs2_addr(decode_io_out_bits_vec_1_rs2_addr),
    .io_out_bits_vec_1_rd_addr(decode_io_out_bits_vec_1_rd_addr),
    .io_out_bits_vec_1_rd_en(decode_io_out_bits_vec_1_rd_en),
    .io_out_bits_vec_1_imm(decode_io_out_bits_vec_1_imm),
    .io_out_bits_vec_1_pred_br(decode_io_out_bits_vec_1_pred_br),
    .io_out_bits_vec_1_pred_bpc(decode_io_out_bits_vec_1_pred_bpc),
    .io_flush(decode_io_flush)
  );
  ysyx_210128_Rename rename ( // @[Core.scala 36:22]
    .clock(rename_clock),
    .reset(rename_reset),
    .io_in_ready(rename_io_in_ready),
    .io_in_valid(rename_io_in_valid),
    .io_in_bits_vec_0_valid(rename_io_in_bits_vec_0_valid),
    .io_in_bits_vec_0_pc(rename_io_in_bits_vec_0_pc),
    .io_in_bits_vec_0_npc(rename_io_in_bits_vec_0_npc),
    .io_in_bits_vec_0_inst(rename_io_in_bits_vec_0_inst),
    .io_in_bits_vec_0_fu_code(rename_io_in_bits_vec_0_fu_code),
    .io_in_bits_vec_0_alu_code(rename_io_in_bits_vec_0_alu_code),
    .io_in_bits_vec_0_jmp_code(rename_io_in_bits_vec_0_jmp_code),
    .io_in_bits_vec_0_mem_code(rename_io_in_bits_vec_0_mem_code),
    .io_in_bits_vec_0_mem_size(rename_io_in_bits_vec_0_mem_size),
    .io_in_bits_vec_0_sys_code(rename_io_in_bits_vec_0_sys_code),
    .io_in_bits_vec_0_w_type(rename_io_in_bits_vec_0_w_type),
    .io_in_bits_vec_0_rs1_src(rename_io_in_bits_vec_0_rs1_src),
    .io_in_bits_vec_0_rs2_src(rename_io_in_bits_vec_0_rs2_src),
    .io_in_bits_vec_0_rs1_addr(rename_io_in_bits_vec_0_rs1_addr),
    .io_in_bits_vec_0_rs2_addr(rename_io_in_bits_vec_0_rs2_addr),
    .io_in_bits_vec_0_rd_addr(rename_io_in_bits_vec_0_rd_addr),
    .io_in_bits_vec_0_rd_en(rename_io_in_bits_vec_0_rd_en),
    .io_in_bits_vec_0_imm(rename_io_in_bits_vec_0_imm),
    .io_in_bits_vec_0_pred_br(rename_io_in_bits_vec_0_pred_br),
    .io_in_bits_vec_0_pred_bpc(rename_io_in_bits_vec_0_pred_bpc),
    .io_in_bits_vec_1_valid(rename_io_in_bits_vec_1_valid),
    .io_in_bits_vec_1_pc(rename_io_in_bits_vec_1_pc),
    .io_in_bits_vec_1_npc(rename_io_in_bits_vec_1_npc),
    .io_in_bits_vec_1_inst(rename_io_in_bits_vec_1_inst),
    .io_in_bits_vec_1_fu_code(rename_io_in_bits_vec_1_fu_code),
    .io_in_bits_vec_1_alu_code(rename_io_in_bits_vec_1_alu_code),
    .io_in_bits_vec_1_jmp_code(rename_io_in_bits_vec_1_jmp_code),
    .io_in_bits_vec_1_mem_code(rename_io_in_bits_vec_1_mem_code),
    .io_in_bits_vec_1_mem_size(rename_io_in_bits_vec_1_mem_size),
    .io_in_bits_vec_1_sys_code(rename_io_in_bits_vec_1_sys_code),
    .io_in_bits_vec_1_w_type(rename_io_in_bits_vec_1_w_type),
    .io_in_bits_vec_1_rs1_src(rename_io_in_bits_vec_1_rs1_src),
    .io_in_bits_vec_1_rs2_src(rename_io_in_bits_vec_1_rs2_src),
    .io_in_bits_vec_1_rs1_addr(rename_io_in_bits_vec_1_rs1_addr),
    .io_in_bits_vec_1_rs2_addr(rename_io_in_bits_vec_1_rs2_addr),
    .io_in_bits_vec_1_rd_addr(rename_io_in_bits_vec_1_rd_addr),
    .io_in_bits_vec_1_rd_en(rename_io_in_bits_vec_1_rd_en),
    .io_in_bits_vec_1_imm(rename_io_in_bits_vec_1_imm),
    .io_in_bits_vec_1_pred_br(rename_io_in_bits_vec_1_pred_br),
    .io_in_bits_vec_1_pred_bpc(rename_io_in_bits_vec_1_pred_bpc),
    .io_out_ready(rename_io_out_ready),
    .io_out_valid(rename_io_out_valid),
    .io_out_bits_vec_0_valid(rename_io_out_bits_vec_0_valid),
    .io_out_bits_vec_0_pc(rename_io_out_bits_vec_0_pc),
    .io_out_bits_vec_0_npc(rename_io_out_bits_vec_0_npc),
    .io_out_bits_vec_0_inst(rename_io_out_bits_vec_0_inst),
    .io_out_bits_vec_0_fu_code(rename_io_out_bits_vec_0_fu_code),
    .io_out_bits_vec_0_alu_code(rename_io_out_bits_vec_0_alu_code),
    .io_out_bits_vec_0_jmp_code(rename_io_out_bits_vec_0_jmp_code),
    .io_out_bits_vec_0_mem_code(rename_io_out_bits_vec_0_mem_code),
    .io_out_bits_vec_0_mem_size(rename_io_out_bits_vec_0_mem_size),
    .io_out_bits_vec_0_sys_code(rename_io_out_bits_vec_0_sys_code),
    .io_out_bits_vec_0_w_type(rename_io_out_bits_vec_0_w_type),
    .io_out_bits_vec_0_rs1_src(rename_io_out_bits_vec_0_rs1_src),
    .io_out_bits_vec_0_rs2_src(rename_io_out_bits_vec_0_rs2_src),
    .io_out_bits_vec_0_rd_addr(rename_io_out_bits_vec_0_rd_addr),
    .io_out_bits_vec_0_rd_en(rename_io_out_bits_vec_0_rd_en),
    .io_out_bits_vec_0_imm(rename_io_out_bits_vec_0_imm),
    .io_out_bits_vec_0_pred_br(rename_io_out_bits_vec_0_pred_br),
    .io_out_bits_vec_0_pred_bpc(rename_io_out_bits_vec_0_pred_bpc),
    .io_out_bits_vec_0_rs1_paddr(rename_io_out_bits_vec_0_rs1_paddr),
    .io_out_bits_vec_0_rs2_paddr(rename_io_out_bits_vec_0_rs2_paddr),
    .io_out_bits_vec_0_rd_paddr(rename_io_out_bits_vec_0_rd_paddr),
    .io_out_bits_vec_0_rd_ppaddr(rename_io_out_bits_vec_0_rd_ppaddr),
    .io_out_bits_vec_1_valid(rename_io_out_bits_vec_1_valid),
    .io_out_bits_vec_1_pc(rename_io_out_bits_vec_1_pc),
    .io_out_bits_vec_1_npc(rename_io_out_bits_vec_1_npc),
    .io_out_bits_vec_1_inst(rename_io_out_bits_vec_1_inst),
    .io_out_bits_vec_1_fu_code(rename_io_out_bits_vec_1_fu_code),
    .io_out_bits_vec_1_alu_code(rename_io_out_bits_vec_1_alu_code),
    .io_out_bits_vec_1_jmp_code(rename_io_out_bits_vec_1_jmp_code),
    .io_out_bits_vec_1_mem_code(rename_io_out_bits_vec_1_mem_code),
    .io_out_bits_vec_1_mem_size(rename_io_out_bits_vec_1_mem_size),
    .io_out_bits_vec_1_sys_code(rename_io_out_bits_vec_1_sys_code),
    .io_out_bits_vec_1_w_type(rename_io_out_bits_vec_1_w_type),
    .io_out_bits_vec_1_rs1_src(rename_io_out_bits_vec_1_rs1_src),
    .io_out_bits_vec_1_rs2_src(rename_io_out_bits_vec_1_rs2_src),
    .io_out_bits_vec_1_rd_addr(rename_io_out_bits_vec_1_rd_addr),
    .io_out_bits_vec_1_rd_en(rename_io_out_bits_vec_1_rd_en),
    .io_out_bits_vec_1_imm(rename_io_out_bits_vec_1_imm),
    .io_out_bits_vec_1_pred_br(rename_io_out_bits_vec_1_pred_br),
    .io_out_bits_vec_1_pred_bpc(rename_io_out_bits_vec_1_pred_bpc),
    .io_out_bits_vec_1_rs1_paddr(rename_io_out_bits_vec_1_rs1_paddr),
    .io_out_bits_vec_1_rs2_paddr(rename_io_out_bits_vec_1_rs2_paddr),
    .io_out_bits_vec_1_rd_paddr(rename_io_out_bits_vec_1_rd_paddr),
    .io_out_bits_vec_1_rd_ppaddr(rename_io_out_bits_vec_1_rd_ppaddr),
    .io_avail_list(rename_io_avail_list),
    .io_flush(rename_io_flush),
    .io_exe_0_valid(rename_io_exe_0_valid),
    .io_exe_0_rd_en(rename_io_exe_0_rd_en),
    .io_exe_0_rd_paddr(rename_io_exe_0_rd_paddr),
    .io_exe_1_valid(rename_io_exe_1_valid),
    .io_exe_1_rd_en(rename_io_exe_1_rd_en),
    .io_exe_1_rd_paddr(rename_io_exe_1_rd_paddr),
    .io_exe_2_valid(rename_io_exe_2_valid),
    .io_exe_2_rd_en(rename_io_exe_2_rd_en),
    .io_exe_2_rd_paddr(rename_io_exe_2_rd_paddr),
    .io_cm_recover(rename_io_cm_recover),
    .io_cm_0_valid(rename_io_cm_0_valid),
    .io_cm_0_rd_addr(rename_io_cm_0_rd_addr),
    .io_cm_0_rd_en(rename_io_cm_0_rd_en),
    .io_cm_0_rd_paddr(rename_io_cm_0_rd_paddr),
    .io_cm_0_rd_ppaddr(rename_io_cm_0_rd_ppaddr),
    .io_cm_1_valid(rename_io_cm_1_valid),
    .io_cm_1_rd_addr(rename_io_cm_1_rd_addr),
    .io_cm_1_rd_en(rename_io_cm_1_rd_en),
    .io_cm_1_rd_paddr(rename_io_cm_1_rd_paddr),
    .io_cm_1_rd_ppaddr(rename_io_cm_1_rd_ppaddr)
  );
  ysyx_210128_StallRegister stall_reg ( // @[Core.scala 42:25]
    .clock(stall_reg_clock),
    .reset(stall_reg_reset),
    .io_flush(stall_reg_io_flush),
    .io_in_ready(stall_reg_io_in_ready),
    .io_in_valid(stall_reg_io_in_valid),
    .io_in_bits_vec_0_valid(stall_reg_io_in_bits_vec_0_valid),
    .io_in_bits_vec_0_pc(stall_reg_io_in_bits_vec_0_pc),
    .io_in_bits_vec_0_npc(stall_reg_io_in_bits_vec_0_npc),
    .io_in_bits_vec_0_inst(stall_reg_io_in_bits_vec_0_inst),
    .io_in_bits_vec_0_fu_code(stall_reg_io_in_bits_vec_0_fu_code),
    .io_in_bits_vec_0_alu_code(stall_reg_io_in_bits_vec_0_alu_code),
    .io_in_bits_vec_0_jmp_code(stall_reg_io_in_bits_vec_0_jmp_code),
    .io_in_bits_vec_0_mem_code(stall_reg_io_in_bits_vec_0_mem_code),
    .io_in_bits_vec_0_mem_size(stall_reg_io_in_bits_vec_0_mem_size),
    .io_in_bits_vec_0_sys_code(stall_reg_io_in_bits_vec_0_sys_code),
    .io_in_bits_vec_0_w_type(stall_reg_io_in_bits_vec_0_w_type),
    .io_in_bits_vec_0_rs1_src(stall_reg_io_in_bits_vec_0_rs1_src),
    .io_in_bits_vec_0_rs2_src(stall_reg_io_in_bits_vec_0_rs2_src),
    .io_in_bits_vec_0_rd_addr(stall_reg_io_in_bits_vec_0_rd_addr),
    .io_in_bits_vec_0_rd_en(stall_reg_io_in_bits_vec_0_rd_en),
    .io_in_bits_vec_0_imm(stall_reg_io_in_bits_vec_0_imm),
    .io_in_bits_vec_0_pred_br(stall_reg_io_in_bits_vec_0_pred_br),
    .io_in_bits_vec_0_pred_bpc(stall_reg_io_in_bits_vec_0_pred_bpc),
    .io_in_bits_vec_0_rs1_paddr(stall_reg_io_in_bits_vec_0_rs1_paddr),
    .io_in_bits_vec_0_rs2_paddr(stall_reg_io_in_bits_vec_0_rs2_paddr),
    .io_in_bits_vec_0_rd_paddr(stall_reg_io_in_bits_vec_0_rd_paddr),
    .io_in_bits_vec_0_rd_ppaddr(stall_reg_io_in_bits_vec_0_rd_ppaddr),
    .io_in_bits_vec_1_valid(stall_reg_io_in_bits_vec_1_valid),
    .io_in_bits_vec_1_pc(stall_reg_io_in_bits_vec_1_pc),
    .io_in_bits_vec_1_npc(stall_reg_io_in_bits_vec_1_npc),
    .io_in_bits_vec_1_inst(stall_reg_io_in_bits_vec_1_inst),
    .io_in_bits_vec_1_fu_code(stall_reg_io_in_bits_vec_1_fu_code),
    .io_in_bits_vec_1_alu_code(stall_reg_io_in_bits_vec_1_alu_code),
    .io_in_bits_vec_1_jmp_code(stall_reg_io_in_bits_vec_1_jmp_code),
    .io_in_bits_vec_1_mem_code(stall_reg_io_in_bits_vec_1_mem_code),
    .io_in_bits_vec_1_mem_size(stall_reg_io_in_bits_vec_1_mem_size),
    .io_in_bits_vec_1_sys_code(stall_reg_io_in_bits_vec_1_sys_code),
    .io_in_bits_vec_1_w_type(stall_reg_io_in_bits_vec_1_w_type),
    .io_in_bits_vec_1_rs1_src(stall_reg_io_in_bits_vec_1_rs1_src),
    .io_in_bits_vec_1_rs2_src(stall_reg_io_in_bits_vec_1_rs2_src),
    .io_in_bits_vec_1_rd_addr(stall_reg_io_in_bits_vec_1_rd_addr),
    .io_in_bits_vec_1_rd_en(stall_reg_io_in_bits_vec_1_rd_en),
    .io_in_bits_vec_1_imm(stall_reg_io_in_bits_vec_1_imm),
    .io_in_bits_vec_1_pred_br(stall_reg_io_in_bits_vec_1_pred_br),
    .io_in_bits_vec_1_pred_bpc(stall_reg_io_in_bits_vec_1_pred_bpc),
    .io_in_bits_vec_1_rs1_paddr(stall_reg_io_in_bits_vec_1_rs1_paddr),
    .io_in_bits_vec_1_rs2_paddr(stall_reg_io_in_bits_vec_1_rs2_paddr),
    .io_in_bits_vec_1_rd_paddr(stall_reg_io_in_bits_vec_1_rd_paddr),
    .io_in_bits_vec_1_rd_ppaddr(stall_reg_io_in_bits_vec_1_rd_ppaddr),
    .io_out_ready(stall_reg_io_out_ready),
    .io_out_valid(stall_reg_io_out_valid),
    .io_out_bits_vec_0_valid(stall_reg_io_out_bits_vec_0_valid),
    .io_out_bits_vec_0_pc(stall_reg_io_out_bits_vec_0_pc),
    .io_out_bits_vec_0_npc(stall_reg_io_out_bits_vec_0_npc),
    .io_out_bits_vec_0_inst(stall_reg_io_out_bits_vec_0_inst),
    .io_out_bits_vec_0_fu_code(stall_reg_io_out_bits_vec_0_fu_code),
    .io_out_bits_vec_0_alu_code(stall_reg_io_out_bits_vec_0_alu_code),
    .io_out_bits_vec_0_jmp_code(stall_reg_io_out_bits_vec_0_jmp_code),
    .io_out_bits_vec_0_mem_code(stall_reg_io_out_bits_vec_0_mem_code),
    .io_out_bits_vec_0_mem_size(stall_reg_io_out_bits_vec_0_mem_size),
    .io_out_bits_vec_0_sys_code(stall_reg_io_out_bits_vec_0_sys_code),
    .io_out_bits_vec_0_w_type(stall_reg_io_out_bits_vec_0_w_type),
    .io_out_bits_vec_0_rs1_src(stall_reg_io_out_bits_vec_0_rs1_src),
    .io_out_bits_vec_0_rs2_src(stall_reg_io_out_bits_vec_0_rs2_src),
    .io_out_bits_vec_0_rd_addr(stall_reg_io_out_bits_vec_0_rd_addr),
    .io_out_bits_vec_0_rd_en(stall_reg_io_out_bits_vec_0_rd_en),
    .io_out_bits_vec_0_imm(stall_reg_io_out_bits_vec_0_imm),
    .io_out_bits_vec_0_pred_br(stall_reg_io_out_bits_vec_0_pred_br),
    .io_out_bits_vec_0_pred_bpc(stall_reg_io_out_bits_vec_0_pred_bpc),
    .io_out_bits_vec_0_rs1_paddr(stall_reg_io_out_bits_vec_0_rs1_paddr),
    .io_out_bits_vec_0_rs2_paddr(stall_reg_io_out_bits_vec_0_rs2_paddr),
    .io_out_bits_vec_0_rd_paddr(stall_reg_io_out_bits_vec_0_rd_paddr),
    .io_out_bits_vec_0_rd_ppaddr(stall_reg_io_out_bits_vec_0_rd_ppaddr),
    .io_out_bits_vec_1_valid(stall_reg_io_out_bits_vec_1_valid),
    .io_out_bits_vec_1_pc(stall_reg_io_out_bits_vec_1_pc),
    .io_out_bits_vec_1_npc(stall_reg_io_out_bits_vec_1_npc),
    .io_out_bits_vec_1_inst(stall_reg_io_out_bits_vec_1_inst),
    .io_out_bits_vec_1_fu_code(stall_reg_io_out_bits_vec_1_fu_code),
    .io_out_bits_vec_1_alu_code(stall_reg_io_out_bits_vec_1_alu_code),
    .io_out_bits_vec_1_jmp_code(stall_reg_io_out_bits_vec_1_jmp_code),
    .io_out_bits_vec_1_mem_code(stall_reg_io_out_bits_vec_1_mem_code),
    .io_out_bits_vec_1_mem_size(stall_reg_io_out_bits_vec_1_mem_size),
    .io_out_bits_vec_1_sys_code(stall_reg_io_out_bits_vec_1_sys_code),
    .io_out_bits_vec_1_w_type(stall_reg_io_out_bits_vec_1_w_type),
    .io_out_bits_vec_1_rs1_src(stall_reg_io_out_bits_vec_1_rs1_src),
    .io_out_bits_vec_1_rs2_src(stall_reg_io_out_bits_vec_1_rs2_src),
    .io_out_bits_vec_1_rd_addr(stall_reg_io_out_bits_vec_1_rd_addr),
    .io_out_bits_vec_1_rd_en(stall_reg_io_out_bits_vec_1_rd_en),
    .io_out_bits_vec_1_imm(stall_reg_io_out_bits_vec_1_imm),
    .io_out_bits_vec_1_pred_br(stall_reg_io_out_bits_vec_1_pred_br),
    .io_out_bits_vec_1_pred_bpc(stall_reg_io_out_bits_vec_1_pred_bpc),
    .io_out_bits_vec_1_rs1_paddr(stall_reg_io_out_bits_vec_1_rs1_paddr),
    .io_out_bits_vec_1_rs2_paddr(stall_reg_io_out_bits_vec_1_rs2_paddr),
    .io_out_bits_vec_1_rd_paddr(stall_reg_io_out_bits_vec_1_rd_paddr),
    .io_out_bits_vec_1_rd_ppaddr(stall_reg_io_out_bits_vec_1_rd_ppaddr)
  );
  ysyx_210128_Rob rob ( // @[Core.scala 46:19]
    .clock(rob_clock),
    .reset(rob_reset),
    .io_in_ready(rob_io_in_ready),
    .io_in_valid(rob_io_in_valid),
    .io_in_bits_vec_0_valid(rob_io_in_bits_vec_0_valid),
    .io_in_bits_vec_0_pc(rob_io_in_bits_vec_0_pc),
    .io_in_bits_vec_0_fu_code(rob_io_in_bits_vec_0_fu_code),
    .io_in_bits_vec_0_sys_code(rob_io_in_bits_vec_0_sys_code),
    .io_in_bits_vec_0_rd_addr(rob_io_in_bits_vec_0_rd_addr),
    .io_in_bits_vec_0_rd_en(rob_io_in_bits_vec_0_rd_en),
    .io_in_bits_vec_0_rd_paddr(rob_io_in_bits_vec_0_rd_paddr),
    .io_in_bits_vec_0_rd_ppaddr(rob_io_in_bits_vec_0_rd_ppaddr),
    .io_in_bits_vec_1_valid(rob_io_in_bits_vec_1_valid),
    .io_in_bits_vec_1_pc(rob_io_in_bits_vec_1_pc),
    .io_in_bits_vec_1_fu_code(rob_io_in_bits_vec_1_fu_code),
    .io_in_bits_vec_1_sys_code(rob_io_in_bits_vec_1_sys_code),
    .io_in_bits_vec_1_rd_addr(rob_io_in_bits_vec_1_rd_addr),
    .io_in_bits_vec_1_rd_en(rob_io_in_bits_vec_1_rd_en),
    .io_in_bits_vec_1_rd_paddr(rob_io_in_bits_vec_1_rd_paddr),
    .io_in_bits_vec_1_rd_ppaddr(rob_io_in_bits_vec_1_rd_ppaddr),
    .io_rob_addr_0(rob_io_rob_addr_0),
    .io_rob_addr_1(rob_io_rob_addr_1),
    .io_exe_0_valid(rob_io_exe_0_valid),
    .io_exe_0_rob_addr(rob_io_exe_0_rob_addr),
    .io_exe_1_valid(rob_io_exe_1_valid),
    .io_exe_1_rob_addr(rob_io_exe_1_rob_addr),
    .io_exe_2_valid(rob_io_exe_2_valid),
    .io_exe_2_rob_addr(rob_io_exe_2_rob_addr),
    .io_exe_ecp_0_jmp_valid(rob_io_exe_ecp_0_jmp_valid),
    .io_exe_ecp_0_jmp(rob_io_exe_ecp_0_jmp),
    .io_exe_ecp_0_jmp_pc(rob_io_exe_ecp_0_jmp_pc),
    .io_exe_ecp_0_mis(rob_io_exe_ecp_0_mis),
    .io_exe_ecp_1_jmp_valid(rob_io_exe_ecp_1_jmp_valid),
    .io_exe_ecp_1_jmp(rob_io_exe_ecp_1_jmp),
    .io_exe_ecp_1_jmp_pc(rob_io_exe_ecp_1_jmp_pc),
    .io_exe_ecp_1_mis(rob_io_exe_ecp_1_mis),
    .io_exe_ecp_2_store_valid(rob_io_exe_ecp_2_store_valid),
    .io_cm_0_valid(rob_io_cm_0_valid),
    .io_cm_0_rd_addr(rob_io_cm_0_rd_addr),
    .io_cm_0_rd_en(rob_io_cm_0_rd_en),
    .io_cm_0_rd_paddr(rob_io_cm_0_rd_paddr),
    .io_cm_0_rd_ppaddr(rob_io_cm_0_rd_ppaddr),
    .io_cm_1_valid(rob_io_cm_1_valid),
    .io_cm_1_rd_addr(rob_io_cm_1_rd_addr),
    .io_cm_1_rd_en(rob_io_cm_1_rd_en),
    .io_cm_1_rd_paddr(rob_io_cm_1_rd_paddr),
    .io_cm_1_rd_ppaddr(rob_io_cm_1_rd_ppaddr),
    .io_jmp_packet_valid(rob_io_jmp_packet_valid),
    .io_jmp_packet_inst_pc(rob_io_jmp_packet_inst_pc),
    .io_jmp_packet_jmp(rob_io_jmp_packet_jmp),
    .io_jmp_packet_jmp_pc(rob_io_jmp_packet_jmp_pc),
    .io_jmp_packet_mis(rob_io_jmp_packet_mis),
    .io_jmp_packet_sys(rob_io_jmp_packet_sys),
    .io_sq_deq_req(rob_io_sq_deq_req),
    .io_flush(rob_io_flush),
    .io_sys_ready(rob_io_sys_ready),
    .csr_mip_mtip_intr_0(rob_csr_mip_mtip_intr_0),
    .intr_mcause_0(rob_intr_mcause_0),
    .intr_mstatus_0(rob_intr_mstatus_0),
    .csr_mtvec_idx_0(rob_csr_mtvec_idx_0),
    .csr_mie_mtie_0(rob_csr_mie_mtie_0),
    .intr_0(rob_intr_0),
    .csr_mstatus_0(rob_csr_mstatus_0),
    .intr_mepc_0(rob_intr_mepc_0)
  );
  ysyx_210128_IssueUnit isu ( // @[Core.scala 47:19]
    .clock(isu_clock),
    .reset(isu_reset),
    .io_flush(isu_io_flush),
    .io_in_ready(isu_io_in_ready),
    .io_in_valid(isu_io_in_valid),
    .io_in_bits_vec_0_valid(isu_io_in_bits_vec_0_valid),
    .io_in_bits_vec_0_pc(isu_io_in_bits_vec_0_pc),
    .io_in_bits_vec_0_npc(isu_io_in_bits_vec_0_npc),
    .io_in_bits_vec_0_inst(isu_io_in_bits_vec_0_inst),
    .io_in_bits_vec_0_fu_code(isu_io_in_bits_vec_0_fu_code),
    .io_in_bits_vec_0_alu_code(isu_io_in_bits_vec_0_alu_code),
    .io_in_bits_vec_0_jmp_code(isu_io_in_bits_vec_0_jmp_code),
    .io_in_bits_vec_0_mem_code(isu_io_in_bits_vec_0_mem_code),
    .io_in_bits_vec_0_mem_size(isu_io_in_bits_vec_0_mem_size),
    .io_in_bits_vec_0_sys_code(isu_io_in_bits_vec_0_sys_code),
    .io_in_bits_vec_0_w_type(isu_io_in_bits_vec_0_w_type),
    .io_in_bits_vec_0_rs1_src(isu_io_in_bits_vec_0_rs1_src),
    .io_in_bits_vec_0_rs2_src(isu_io_in_bits_vec_0_rs2_src),
    .io_in_bits_vec_0_rd_en(isu_io_in_bits_vec_0_rd_en),
    .io_in_bits_vec_0_imm(isu_io_in_bits_vec_0_imm),
    .io_in_bits_vec_0_pred_br(isu_io_in_bits_vec_0_pred_br),
    .io_in_bits_vec_0_pred_bpc(isu_io_in_bits_vec_0_pred_bpc),
    .io_in_bits_vec_0_rs1_paddr(isu_io_in_bits_vec_0_rs1_paddr),
    .io_in_bits_vec_0_rs2_paddr(isu_io_in_bits_vec_0_rs2_paddr),
    .io_in_bits_vec_0_rd_paddr(isu_io_in_bits_vec_0_rd_paddr),
    .io_in_bits_vec_1_valid(isu_io_in_bits_vec_1_valid),
    .io_in_bits_vec_1_pc(isu_io_in_bits_vec_1_pc),
    .io_in_bits_vec_1_npc(isu_io_in_bits_vec_1_npc),
    .io_in_bits_vec_1_inst(isu_io_in_bits_vec_1_inst),
    .io_in_bits_vec_1_fu_code(isu_io_in_bits_vec_1_fu_code),
    .io_in_bits_vec_1_alu_code(isu_io_in_bits_vec_1_alu_code),
    .io_in_bits_vec_1_jmp_code(isu_io_in_bits_vec_1_jmp_code),
    .io_in_bits_vec_1_mem_code(isu_io_in_bits_vec_1_mem_code),
    .io_in_bits_vec_1_mem_size(isu_io_in_bits_vec_1_mem_size),
    .io_in_bits_vec_1_sys_code(isu_io_in_bits_vec_1_sys_code),
    .io_in_bits_vec_1_w_type(isu_io_in_bits_vec_1_w_type),
    .io_in_bits_vec_1_rs1_src(isu_io_in_bits_vec_1_rs1_src),
    .io_in_bits_vec_1_rs2_src(isu_io_in_bits_vec_1_rs2_src),
    .io_in_bits_vec_1_rd_en(isu_io_in_bits_vec_1_rd_en),
    .io_in_bits_vec_1_imm(isu_io_in_bits_vec_1_imm),
    .io_in_bits_vec_1_pred_br(isu_io_in_bits_vec_1_pred_br),
    .io_in_bits_vec_1_pred_bpc(isu_io_in_bits_vec_1_pred_bpc),
    .io_in_bits_vec_1_rs1_paddr(isu_io_in_bits_vec_1_rs1_paddr),
    .io_in_bits_vec_1_rs2_paddr(isu_io_in_bits_vec_1_rs2_paddr),
    .io_in_bits_vec_1_rd_paddr(isu_io_in_bits_vec_1_rd_paddr),
    .io_rob_addr_0(isu_io_rob_addr_0),
    .io_rob_addr_1(isu_io_rob_addr_1),
    .io_out_0_valid(isu_io_out_0_valid),
    .io_out_0_pc(isu_io_out_0_pc),
    .io_out_0_npc(isu_io_out_0_npc),
    .io_out_0_inst(isu_io_out_0_inst),
    .io_out_0_fu_code(isu_io_out_0_fu_code),
    .io_out_0_alu_code(isu_io_out_0_alu_code),
    .io_out_0_jmp_code(isu_io_out_0_jmp_code),
    .io_out_0_sys_code(isu_io_out_0_sys_code),
    .io_out_0_w_type(isu_io_out_0_w_type),
    .io_out_0_rs1_src(isu_io_out_0_rs1_src),
    .io_out_0_rs2_src(isu_io_out_0_rs2_src),
    .io_out_0_rd_en(isu_io_out_0_rd_en),
    .io_out_0_imm(isu_io_out_0_imm),
    .io_out_0_pred_br(isu_io_out_0_pred_br),
    .io_out_0_pred_bpc(isu_io_out_0_pred_bpc),
    .io_out_0_rs1_paddr(isu_io_out_0_rs1_paddr),
    .io_out_0_rs2_paddr(isu_io_out_0_rs2_paddr),
    .io_out_0_rd_paddr(isu_io_out_0_rd_paddr),
    .io_out_0_rob_addr(isu_io_out_0_rob_addr),
    .io_out_1_valid(isu_io_out_1_valid),
    .io_out_1_pc(isu_io_out_1_pc),
    .io_out_1_npc(isu_io_out_1_npc),
    .io_out_1_fu_code(isu_io_out_1_fu_code),
    .io_out_1_alu_code(isu_io_out_1_alu_code),
    .io_out_1_jmp_code(isu_io_out_1_jmp_code),
    .io_out_1_w_type(isu_io_out_1_w_type),
    .io_out_1_rs1_src(isu_io_out_1_rs1_src),
    .io_out_1_rs2_src(isu_io_out_1_rs2_src),
    .io_out_1_rd_en(isu_io_out_1_rd_en),
    .io_out_1_imm(isu_io_out_1_imm),
    .io_out_1_pred_br(isu_io_out_1_pred_br),
    .io_out_1_pred_bpc(isu_io_out_1_pred_bpc),
    .io_out_1_rs1_paddr(isu_io_out_1_rs1_paddr),
    .io_out_1_rs2_paddr(isu_io_out_1_rs2_paddr),
    .io_out_1_rd_paddr(isu_io_out_1_rd_paddr),
    .io_out_1_rob_addr(isu_io_out_1_rob_addr),
    .io_out_2_valid(isu_io_out_2_valid),
    .io_out_2_pc(isu_io_out_2_pc),
    .io_out_2_fu_code(isu_io_out_2_fu_code),
    .io_out_2_alu_code(isu_io_out_2_alu_code),
    .io_out_2_mem_code(isu_io_out_2_mem_code),
    .io_out_2_mem_size(isu_io_out_2_mem_size),
    .io_out_2_w_type(isu_io_out_2_w_type),
    .io_out_2_rs1_src(isu_io_out_2_rs1_src),
    .io_out_2_rs2_src(isu_io_out_2_rs2_src),
    .io_out_2_rd_en(isu_io_out_2_rd_en),
    .io_out_2_imm(isu_io_out_2_imm),
    .io_out_2_rs1_paddr(isu_io_out_2_rs1_paddr),
    .io_out_2_rs2_paddr(isu_io_out_2_rs2_paddr),
    .io_out_2_rd_paddr(isu_io_out_2_rd_paddr),
    .io_out_2_rob_addr(isu_io_out_2_rob_addr),
    .io_avail_list(isu_io_avail_list),
    .io_lsu_ready(isu_io_lsu_ready),
    .io_sys_ready(isu_io_sys_ready)
  );
  ysyx_210128_Prf rf ( // @[Core.scala 70:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_in_0_valid(rf_io_in_0_valid),
    .io_in_0_pc(rf_io_in_0_pc),
    .io_in_0_npc(rf_io_in_0_npc),
    .io_in_0_inst(rf_io_in_0_inst),
    .io_in_0_fu_code(rf_io_in_0_fu_code),
    .io_in_0_alu_code(rf_io_in_0_alu_code),
    .io_in_0_jmp_code(rf_io_in_0_jmp_code),
    .io_in_0_sys_code(rf_io_in_0_sys_code),
    .io_in_0_w_type(rf_io_in_0_w_type),
    .io_in_0_rs1_src(rf_io_in_0_rs1_src),
    .io_in_0_rs2_src(rf_io_in_0_rs2_src),
    .io_in_0_rd_en(rf_io_in_0_rd_en),
    .io_in_0_imm(rf_io_in_0_imm),
    .io_in_0_pred_br(rf_io_in_0_pred_br),
    .io_in_0_pred_bpc(rf_io_in_0_pred_bpc),
    .io_in_0_rs1_paddr(rf_io_in_0_rs1_paddr),
    .io_in_0_rs2_paddr(rf_io_in_0_rs2_paddr),
    .io_in_0_rd_paddr(rf_io_in_0_rd_paddr),
    .io_in_0_rob_addr(rf_io_in_0_rob_addr),
    .io_in_1_valid(rf_io_in_1_valid),
    .io_in_1_pc(rf_io_in_1_pc),
    .io_in_1_npc(rf_io_in_1_npc),
    .io_in_1_fu_code(rf_io_in_1_fu_code),
    .io_in_1_alu_code(rf_io_in_1_alu_code),
    .io_in_1_jmp_code(rf_io_in_1_jmp_code),
    .io_in_1_w_type(rf_io_in_1_w_type),
    .io_in_1_rs1_src(rf_io_in_1_rs1_src),
    .io_in_1_rs2_src(rf_io_in_1_rs2_src),
    .io_in_1_rd_en(rf_io_in_1_rd_en),
    .io_in_1_imm(rf_io_in_1_imm),
    .io_in_1_pred_br(rf_io_in_1_pred_br),
    .io_in_1_pred_bpc(rf_io_in_1_pred_bpc),
    .io_in_1_rs1_paddr(rf_io_in_1_rs1_paddr),
    .io_in_1_rs2_paddr(rf_io_in_1_rs2_paddr),
    .io_in_1_rd_paddr(rf_io_in_1_rd_paddr),
    .io_in_1_rob_addr(rf_io_in_1_rob_addr),
    .io_in_2_valid(rf_io_in_2_valid),
    .io_in_2_pc(rf_io_in_2_pc),
    .io_in_2_fu_code(rf_io_in_2_fu_code),
    .io_in_2_alu_code(rf_io_in_2_alu_code),
    .io_in_2_mem_code(rf_io_in_2_mem_code),
    .io_in_2_mem_size(rf_io_in_2_mem_size),
    .io_in_2_w_type(rf_io_in_2_w_type),
    .io_in_2_rs1_src(rf_io_in_2_rs1_src),
    .io_in_2_rs2_src(rf_io_in_2_rs2_src),
    .io_in_2_rd_en(rf_io_in_2_rd_en),
    .io_in_2_imm(rf_io_in_2_imm),
    .io_in_2_rs1_paddr(rf_io_in_2_rs1_paddr),
    .io_in_2_rs2_paddr(rf_io_in_2_rs2_paddr),
    .io_in_2_rd_paddr(rf_io_in_2_rd_paddr),
    .io_in_2_rob_addr(rf_io_in_2_rob_addr),
    .io_out_0_valid(rf_io_out_0_valid),
    .io_out_0_pc(rf_io_out_0_pc),
    .io_out_0_npc(rf_io_out_0_npc),
    .io_out_0_inst(rf_io_out_0_inst),
    .io_out_0_fu_code(rf_io_out_0_fu_code),
    .io_out_0_alu_code(rf_io_out_0_alu_code),
    .io_out_0_jmp_code(rf_io_out_0_jmp_code),
    .io_out_0_sys_code(rf_io_out_0_sys_code),
    .io_out_0_w_type(rf_io_out_0_w_type),
    .io_out_0_rs1_src(rf_io_out_0_rs1_src),
    .io_out_0_rs2_src(rf_io_out_0_rs2_src),
    .io_out_0_rd_en(rf_io_out_0_rd_en),
    .io_out_0_imm(rf_io_out_0_imm),
    .io_out_0_pred_br(rf_io_out_0_pred_br),
    .io_out_0_pred_bpc(rf_io_out_0_pred_bpc),
    .io_out_0_rd_paddr(rf_io_out_0_rd_paddr),
    .io_out_0_rob_addr(rf_io_out_0_rob_addr),
    .io_out_1_valid(rf_io_out_1_valid),
    .io_out_1_pc(rf_io_out_1_pc),
    .io_out_1_npc(rf_io_out_1_npc),
    .io_out_1_fu_code(rf_io_out_1_fu_code),
    .io_out_1_alu_code(rf_io_out_1_alu_code),
    .io_out_1_jmp_code(rf_io_out_1_jmp_code),
    .io_out_1_w_type(rf_io_out_1_w_type),
    .io_out_1_rs1_src(rf_io_out_1_rs1_src),
    .io_out_1_rs2_src(rf_io_out_1_rs2_src),
    .io_out_1_rd_en(rf_io_out_1_rd_en),
    .io_out_1_imm(rf_io_out_1_imm),
    .io_out_1_pred_br(rf_io_out_1_pred_br),
    .io_out_1_pred_bpc(rf_io_out_1_pred_bpc),
    .io_out_1_rd_paddr(rf_io_out_1_rd_paddr),
    .io_out_1_rob_addr(rf_io_out_1_rob_addr),
    .io_out_2_valid(rf_io_out_2_valid),
    .io_out_2_pc(rf_io_out_2_pc),
    .io_out_2_fu_code(rf_io_out_2_fu_code),
    .io_out_2_alu_code(rf_io_out_2_alu_code),
    .io_out_2_mem_code(rf_io_out_2_mem_code),
    .io_out_2_mem_size(rf_io_out_2_mem_size),
    .io_out_2_w_type(rf_io_out_2_w_type),
    .io_out_2_rs1_src(rf_io_out_2_rs1_src),
    .io_out_2_rs2_src(rf_io_out_2_rs2_src),
    .io_out_2_rd_en(rf_io_out_2_rd_en),
    .io_out_2_imm(rf_io_out_2_imm),
    .io_out_2_rd_paddr(rf_io_out_2_rd_paddr),
    .io_out_2_rob_addr(rf_io_out_2_rob_addr),
    .io_rs1_data_0(rf_io_rs1_data_0),
    .io_rs1_data_1(rf_io_rs1_data_1),
    .io_rs1_data_2(rf_io_rs1_data_2),
    .io_rs2_data_0(rf_io_rs2_data_0),
    .io_rs2_data_1(rf_io_rs2_data_1),
    .io_rs2_data_2(rf_io_rs2_data_2),
    .io_rd_en_0(rf_io_rd_en_0),
    .io_rd_en_1(rf_io_rd_en_1),
    .io_rd_en_2(rf_io_rd_en_2),
    .io_rd_paddr_0(rf_io_rd_paddr_0),
    .io_rd_paddr_1(rf_io_rd_paddr_1),
    .io_rd_paddr_2(rf_io_rd_paddr_2),
    .io_rd_data_0(rf_io_rd_data_0),
    .io_rd_data_1(rf_io_rd_data_1),
    .io_rd_data_2(rf_io_rd_data_2),
    .io_flush(rf_io_flush)
  );
  ysyx_210128_Execution execution ( // @[Core.scala 76:25]
    .clock(execution_clock),
    .reset(execution_reset),
    .io_in_0_valid(execution_io_in_0_valid),
    .io_in_0_pc(execution_io_in_0_pc),
    .io_in_0_npc(execution_io_in_0_npc),
    .io_in_0_inst(execution_io_in_0_inst),
    .io_in_0_fu_code(execution_io_in_0_fu_code),
    .io_in_0_alu_code(execution_io_in_0_alu_code),
    .io_in_0_jmp_code(execution_io_in_0_jmp_code),
    .io_in_0_sys_code(execution_io_in_0_sys_code),
    .io_in_0_w_type(execution_io_in_0_w_type),
    .io_in_0_rs1_src(execution_io_in_0_rs1_src),
    .io_in_0_rs2_src(execution_io_in_0_rs2_src),
    .io_in_0_rd_en(execution_io_in_0_rd_en),
    .io_in_0_imm(execution_io_in_0_imm),
    .io_in_0_pred_br(execution_io_in_0_pred_br),
    .io_in_0_pred_bpc(execution_io_in_0_pred_bpc),
    .io_in_0_rd_paddr(execution_io_in_0_rd_paddr),
    .io_in_0_rob_addr(execution_io_in_0_rob_addr),
    .io_in_1_valid(execution_io_in_1_valid),
    .io_in_1_pc(execution_io_in_1_pc),
    .io_in_1_npc(execution_io_in_1_npc),
    .io_in_1_fu_code(execution_io_in_1_fu_code),
    .io_in_1_alu_code(execution_io_in_1_alu_code),
    .io_in_1_jmp_code(execution_io_in_1_jmp_code),
    .io_in_1_w_type(execution_io_in_1_w_type),
    .io_in_1_rs1_src(execution_io_in_1_rs1_src),
    .io_in_1_rs2_src(execution_io_in_1_rs2_src),
    .io_in_1_rd_en(execution_io_in_1_rd_en),
    .io_in_1_imm(execution_io_in_1_imm),
    .io_in_1_pred_br(execution_io_in_1_pred_br),
    .io_in_1_pred_bpc(execution_io_in_1_pred_bpc),
    .io_in_1_rd_paddr(execution_io_in_1_rd_paddr),
    .io_in_1_rob_addr(execution_io_in_1_rob_addr),
    .io_in_2_valid(execution_io_in_2_valid),
    .io_in_2_pc(execution_io_in_2_pc),
    .io_in_2_fu_code(execution_io_in_2_fu_code),
    .io_in_2_alu_code(execution_io_in_2_alu_code),
    .io_in_2_mem_code(execution_io_in_2_mem_code),
    .io_in_2_mem_size(execution_io_in_2_mem_size),
    .io_in_2_w_type(execution_io_in_2_w_type),
    .io_in_2_rs1_src(execution_io_in_2_rs1_src),
    .io_in_2_rs2_src(execution_io_in_2_rs2_src),
    .io_in_2_rd_en(execution_io_in_2_rd_en),
    .io_in_2_imm(execution_io_in_2_imm),
    .io_in_2_rd_paddr(execution_io_in_2_rd_paddr),
    .io_in_2_rob_addr(execution_io_in_2_rob_addr),
    .io_rs1_data_0(execution_io_rs1_data_0),
    .io_rs1_data_1(execution_io_rs1_data_1),
    .io_rs1_data_2(execution_io_rs1_data_2),
    .io_rs2_data_0(execution_io_rs2_data_0),
    .io_rs2_data_1(execution_io_rs2_data_1),
    .io_rs2_data_2(execution_io_rs2_data_2),
    .io_out_0_valid(execution_io_out_0_valid),
    .io_out_0_rob_addr(execution_io_out_0_rob_addr),
    .io_out_1_valid(execution_io_out_1_valid),
    .io_out_1_rob_addr(execution_io_out_1_rob_addr),
    .io_out_2_valid(execution_io_out_2_valid),
    .io_out_2_rob_addr(execution_io_out_2_rob_addr),
    .io_out_ecp_0_jmp_valid(execution_io_out_ecp_0_jmp_valid),
    .io_out_ecp_0_jmp(execution_io_out_ecp_0_jmp),
    .io_out_ecp_0_jmp_pc(execution_io_out_ecp_0_jmp_pc),
    .io_out_ecp_0_mis(execution_io_out_ecp_0_mis),
    .io_out_ecp_1_jmp_valid(execution_io_out_ecp_1_jmp_valid),
    .io_out_ecp_1_jmp(execution_io_out_ecp_1_jmp),
    .io_out_ecp_1_jmp_pc(execution_io_out_ecp_1_jmp_pc),
    .io_out_ecp_1_mis(execution_io_out_ecp_1_mis),
    .io_out_ecp_2_store_valid(execution_io_out_ecp_2_store_valid),
    .io_rd_en_0(execution_io_rd_en_0),
    .io_rd_en_1(execution_io_rd_en_1),
    .io_rd_en_2(execution_io_rd_en_2),
    .io_rd_paddr_0(execution_io_rd_paddr_0),
    .io_rd_paddr_1(execution_io_rd_paddr_1),
    .io_rd_paddr_2(execution_io_rd_paddr_2),
    .io_rd_data_0(execution_io_rd_data_0),
    .io_rd_data_1(execution_io_rd_data_1),
    .io_rd_data_2(execution_io_rd_data_2),
    .io_flush(execution_io_flush),
    .io_lsu_ready(execution_io_lsu_ready),
    .io_dmem_st_req_ready(execution_io_dmem_st_req_ready),
    .io_dmem_st_req_valid(execution_io_dmem_st_req_valid),
    .io_dmem_st_req_bits_addr(execution_io_dmem_st_req_bits_addr),
    .io_dmem_st_req_bits_wdata(execution_io_dmem_st_req_bits_wdata),
    .io_dmem_st_req_bits_wmask(execution_io_dmem_st_req_bits_wmask),
    .io_dmem_st_req_bits_size(execution_io_dmem_st_req_bits_size),
    .io_dmem_st_resp_ready(execution_io_dmem_st_resp_ready),
    .io_dmem_st_resp_valid(execution_io_dmem_st_resp_valid),
    .io_dmem_ld_req_ready(execution_io_dmem_ld_req_ready),
    .io_dmem_ld_req_valid(execution_io_dmem_ld_req_valid),
    .io_dmem_ld_req_bits_addr(execution_io_dmem_ld_req_bits_addr),
    .io_dmem_ld_req_bits_size(execution_io_dmem_ld_req_bits_size),
    .io_dmem_ld_resp_ready(execution_io_dmem_ld_resp_ready),
    .io_dmem_ld_resp_valid(execution_io_dmem_ld_resp_valid),
    .io_dmem_ld_resp_bits_rdata(execution_io_dmem_ld_resp_bits_rdata),
    .io_lsu_wakeup_uop_valid(execution_io_lsu_wakeup_uop_valid),
    .io_lsu_wakeup_uop_rd_en(execution_io_lsu_wakeup_uop_rd_en),
    .io_lsu_wakeup_uop_rd_paddr(execution_io_lsu_wakeup_uop_rd_paddr),
    .mtip(execution_mtip),
    .intr_mcause(execution_intr_mcause),
    .instr_cnt(execution_instr_cnt),
    .intr_mstatus(execution_intr_mstatus),
    ._T_6_0(execution__T_6_0),
    ._T_5_0(execution__T_5_0),
    .intr(execution_intr),
    .fence_i(execution_fence_i),
    .cycle_cnt(execution_cycle_cnt),
    .mstatus(execution_mstatus),
    .intr_mepc(execution_intr_mepc),
    .mtip_0(execution_mtip_0)
  );
  ysyx_210128_StoreQueue sq ( // @[Core.scala 95:18]
    .clock(sq_clock),
    .reset(sq_reset),
    .io_flush(sq_io_flush),
    .io_in_st_req_ready(sq_io_in_st_req_ready),
    .io_in_st_req_valid(sq_io_in_st_req_valid),
    .io_in_st_req_bits_addr(sq_io_in_st_req_bits_addr),
    .io_in_st_req_bits_wdata(sq_io_in_st_req_bits_wdata),
    .io_in_st_req_bits_wmask(sq_io_in_st_req_bits_wmask),
    .io_in_st_req_bits_size(sq_io_in_st_req_bits_size),
    .io_in_st_resp_ready(sq_io_in_st_resp_ready),
    .io_in_st_resp_valid(sq_io_in_st_resp_valid),
    .io_in_ld_req_ready(sq_io_in_ld_req_ready),
    .io_in_ld_req_valid(sq_io_in_ld_req_valid),
    .io_in_ld_req_bits_addr(sq_io_in_ld_req_bits_addr),
    .io_in_ld_req_bits_size(sq_io_in_ld_req_bits_size),
    .io_in_ld_resp_ready(sq_io_in_ld_resp_ready),
    .io_in_ld_resp_valid(sq_io_in_ld_resp_valid),
    .io_in_ld_resp_bits_rdata(sq_io_in_ld_resp_bits_rdata),
    .io_out_st_req_ready(sq_io_out_st_req_ready),
    .io_out_st_req_valid(sq_io_out_st_req_valid),
    .io_out_st_req_bits_addr(sq_io_out_st_req_bits_addr),
    .io_out_st_req_bits_wdata(sq_io_out_st_req_bits_wdata),
    .io_out_st_req_bits_wmask(sq_io_out_st_req_bits_wmask),
    .io_out_st_req_bits_size(sq_io_out_st_req_bits_size),
    .io_out_st_resp_ready(sq_io_out_st_resp_ready),
    .io_out_st_resp_valid(sq_io_out_st_resp_valid),
    .io_out_ld_req_ready(sq_io_out_ld_req_ready),
    .io_out_ld_req_valid(sq_io_out_ld_req_valid),
    .io_out_ld_req_bits_addr(sq_io_out_ld_req_bits_addr),
    .io_out_ld_req_bits_size(sq_io_out_ld_req_bits_size),
    .io_out_ld_resp_ready(sq_io_out_ld_resp_ready),
    .io_out_ld_resp_valid(sq_io_out_ld_resp_valid),
    .io_out_ld_resp_bits_rdata(sq_io_out_ld_resp_bits_rdata),
    .io_deq_req(sq_io_deq_req),
    .empty_0(sq_empty_0)
  );
  ysyx_210128_CacheBusCrossbarNto1 crossbar2to1 ( // @[Core.scala 101:28]
    .clock(crossbar2to1_clock),
    .io_in_0_req_ready(crossbar2to1_io_in_0_req_ready),
    .io_in_0_req_valid(crossbar2to1_io_in_0_req_valid),
    .io_in_0_req_bits_addr(crossbar2to1_io_in_0_req_bits_addr),
    .io_in_0_req_bits_wdata(crossbar2to1_io_in_0_req_bits_wdata),
    .io_in_0_req_bits_wmask(crossbar2to1_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_size(crossbar2to1_io_in_0_req_bits_size),
    .io_in_0_resp_ready(crossbar2to1_io_in_0_resp_ready),
    .io_in_0_resp_valid(crossbar2to1_io_in_0_resp_valid),
    .io_in_1_req_ready(crossbar2to1_io_in_1_req_ready),
    .io_in_1_req_valid(crossbar2to1_io_in_1_req_valid),
    .io_in_1_req_bits_addr(crossbar2to1_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(crossbar2to1_io_in_1_req_bits_size),
    .io_in_1_resp_ready(crossbar2to1_io_in_1_resp_ready),
    .io_in_1_resp_valid(crossbar2to1_io_in_1_resp_valid),
    .io_in_1_resp_bits_rdata(crossbar2to1_io_in_1_resp_bits_rdata),
    .io_out_req_ready(crossbar2to1_io_out_req_ready),
    .io_out_req_valid(crossbar2to1_io_out_req_valid),
    .io_out_req_bits_id(crossbar2to1_io_out_req_bits_id),
    .io_out_req_bits_addr(crossbar2to1_io_out_req_bits_addr),
    .io_out_req_bits_wdata(crossbar2to1_io_out_req_bits_wdata),
    .io_out_req_bits_wmask(crossbar2to1_io_out_req_bits_wmask),
    .io_out_req_bits_wen(crossbar2to1_io_out_req_bits_wen),
    .io_out_req_bits_size(crossbar2to1_io_out_req_bits_size),
    .io_out_resp_ready(crossbar2to1_io_out_resp_ready),
    .io_out_resp_valid(crossbar2to1_io_out_resp_valid),
    .io_out_resp_bits_id(crossbar2to1_io_out_resp_bits_id),
    .io_out_resp_bits_rdata(crossbar2to1_io_out_resp_bits_rdata)
  );
  ysyx_210128_CacheBusCrossbar1to2_1 crossbar1to2 ( // @[Core.scala 105:28]
    .clock(crossbar1to2_clock),
    .reset(crossbar1to2_reset),
    .io_in_req_ready(crossbar1to2_io_in_req_ready),
    .io_in_req_valid(crossbar1to2_io_in_req_valid),
    .io_in_req_bits_id(crossbar1to2_io_in_req_bits_id),
    .io_in_req_bits_addr(crossbar1to2_io_in_req_bits_addr),
    .io_in_req_bits_wdata(crossbar1to2_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(crossbar1to2_io_in_req_bits_wmask),
    .io_in_req_bits_wen(crossbar1to2_io_in_req_bits_wen),
    .io_in_req_bits_size(crossbar1to2_io_in_req_bits_size),
    .io_in_resp_ready(crossbar1to2_io_in_resp_ready),
    .io_in_resp_valid(crossbar1to2_io_in_resp_valid),
    .io_in_resp_bits_id(crossbar1to2_io_in_resp_bits_id),
    .io_in_resp_bits_rdata(crossbar1to2_io_in_resp_bits_rdata),
    .io_out_0_req_ready(crossbar1to2_io_out_0_req_ready),
    .io_out_0_req_valid(crossbar1to2_io_out_0_req_valid),
    .io_out_0_req_bits_id(crossbar1to2_io_out_0_req_bits_id),
    .io_out_0_req_bits_addr(crossbar1to2_io_out_0_req_bits_addr),
    .io_out_0_req_bits_wdata(crossbar1to2_io_out_0_req_bits_wdata),
    .io_out_0_req_bits_wmask(crossbar1to2_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wen(crossbar1to2_io_out_0_req_bits_wen),
    .io_out_0_req_bits_size(crossbar1to2_io_out_0_req_bits_size),
    .io_out_0_resp_ready(crossbar1to2_io_out_0_resp_ready),
    .io_out_0_resp_valid(crossbar1to2_io_out_0_resp_valid),
    .io_out_0_resp_bits_id(crossbar1to2_io_out_0_resp_bits_id),
    .io_out_0_resp_bits_rdata(crossbar1to2_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(crossbar1to2_io_out_1_req_ready),
    .io_out_1_req_valid(crossbar1to2_io_out_1_req_valid),
    .io_out_1_req_bits_id(crossbar1to2_io_out_1_req_bits_id),
    .io_out_1_req_bits_addr(crossbar1to2_io_out_1_req_bits_addr),
    .io_out_1_req_bits_wdata(crossbar1to2_io_out_1_req_bits_wdata),
    .io_out_1_req_bits_wmask(crossbar1to2_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wen(crossbar1to2_io_out_1_req_bits_wen),
    .io_out_1_req_bits_size(crossbar1to2_io_out_1_req_bits_size),
    .io_out_1_resp_ready(crossbar1to2_io_out_1_resp_ready),
    .io_out_1_resp_valid(crossbar1to2_io_out_1_resp_valid),
    .io_out_1_resp_bits_id(crossbar1to2_io_out_1_resp_bits_id),
    .io_out_1_resp_bits_rdata(crossbar1to2_io_out_1_resp_bits_rdata),
    .io_to_1(crossbar1to2_io_to_1)
  );
  ysyx_210128_CacheController_1 dcache ( // @[Core.scala 112:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_in_req_ready(dcache_io_in_req_ready),
    .io_in_req_valid(dcache_io_in_req_valid),
    .io_in_req_bits_id(dcache_io_in_req_bits_id),
    .io_in_req_bits_addr(dcache_io_in_req_bits_addr),
    .io_in_req_bits_wdata(dcache_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(dcache_io_in_req_bits_wmask),
    .io_in_req_bits_wen(dcache_io_in_req_bits_wen),
    .io_in_req_bits_size(dcache_io_in_req_bits_size),
    .io_in_resp_ready(dcache_io_in_resp_ready),
    .io_in_resp_valid(dcache_io_in_resp_valid),
    .io_in_resp_bits_id(dcache_io_in_resp_bits_id),
    .io_in_resp_bits_rdata(dcache_io_in_resp_bits_rdata),
    .io_out_cache_req_ready(dcache_io_out_cache_req_ready),
    .io_out_cache_req_valid(dcache_io_out_cache_req_valid),
    .io_out_cache_req_bits_addr(dcache_io_out_cache_req_bits_addr),
    .io_out_cache_req_bits_aen(dcache_io_out_cache_req_bits_aen),
    .io_out_cache_req_bits_wdata(dcache_io_out_cache_req_bits_wdata),
    .io_out_cache_req_bits_wlast(dcache_io_out_cache_req_bits_wlast),
    .io_out_cache_req_bits_wen(dcache_io_out_cache_req_bits_wen),
    .io_out_cache_resp_ready(dcache_io_out_cache_resp_ready),
    .io_out_cache_resp_valid(dcache_io_out_cache_resp_valid),
    .io_out_cache_resp_bits_rdata(dcache_io_out_cache_resp_bits_rdata),
    .io_out_cache_resp_bits_rlast(dcache_io_out_cache_resp_bits_rlast),
    .io_out_uncache_req_ready(dcache_io_out_uncache_req_ready),
    .io_out_uncache_req_valid(dcache_io_out_uncache_req_valid),
    .io_out_uncache_req_bits_addr(dcache_io_out_uncache_req_bits_addr),
    .io_out_uncache_req_bits_wdata(dcache_io_out_uncache_req_bits_wdata),
    .io_out_uncache_req_bits_wmask(dcache_io_out_uncache_req_bits_wmask),
    .io_out_uncache_req_bits_wen(dcache_io_out_uncache_req_bits_wen),
    .io_out_uncache_req_bits_size(dcache_io_out_uncache_req_bits_size),
    .io_out_uncache_resp_ready(dcache_io_out_uncache_resp_ready),
    .io_out_uncache_resp_valid(dcache_io_out_uncache_resp_valid),
    .io_out_uncache_resp_bits_rdata(dcache_io_out_uncache_resp_bits_rdata),
    .fence_i(dcache_fence_i),
    ._WIRE_10(dcache__WIRE_10),
    .empty(dcache_empty)
  );
  ysyx_210128_Clint clint ( // @[Core.scala 117:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io_in_req_ready(clint_io_in_req_ready),
    .io_in_req_valid(clint_io_in_req_valid),
    .io_in_req_bits_id(clint_io_in_req_bits_id),
    .io_in_req_bits_addr(clint_io_in_req_bits_addr),
    .io_in_req_bits_wdata(clint_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(clint_io_in_req_bits_wmask),
    .io_in_req_bits_wen(clint_io_in_req_bits_wen),
    .io_in_resp_ready(clint_io_in_resp_ready),
    .io_in_resp_valid(clint_io_in_resp_valid),
    .io_in_resp_bits_id(clint_io_in_resp_bits_id),
    .io_in_resp_bits_rdata(clint_io_in_resp_bits_rdata),
    .mtip_1(clint_mtip_1)
  );
  assign io_core_bus_0_req_valid = icache_io_out_cache_req_valid; // @[Core.scala 21:23]
  assign io_core_bus_0_req_bits_addr = icache_io_out_cache_req_bits_addr; // @[Core.scala 21:23]
  assign io_core_bus_0_req_bits_aen = icache_io_out_cache_req_bits_aen; // @[Core.scala 21:23]
  assign io_core_bus_0_req_bits_wdata = icache_io_out_cache_req_bits_wdata; // @[Core.scala 21:23]
  assign io_core_bus_0_req_bits_wlast = icache_io_out_cache_req_bits_wlast; // @[Core.scala 21:23]
  assign io_core_bus_0_req_bits_wen = icache_io_out_cache_req_bits_wen; // @[Core.scala 21:23]
  assign io_core_bus_0_resp_ready = icache_io_out_cache_resp_ready; // @[Core.scala 21:23]
  assign io_core_bus_1_req_valid = dcache_io_out_cache_req_valid; // @[Core.scala 114:23]
  assign io_core_bus_1_req_bits_addr = dcache_io_out_cache_req_bits_addr; // @[Core.scala 114:23]
  assign io_core_bus_1_req_bits_aen = dcache_io_out_cache_req_bits_aen; // @[Core.scala 114:23]
  assign io_core_bus_1_req_bits_wdata = dcache_io_out_cache_req_bits_wdata; // @[Core.scala 114:23]
  assign io_core_bus_1_req_bits_wlast = dcache_io_out_cache_req_bits_wlast; // @[Core.scala 114:23]
  assign io_core_bus_1_req_bits_wen = dcache_io_out_cache_req_bits_wen; // @[Core.scala 114:23]
  assign io_core_bus_1_resp_ready = dcache_io_out_cache_resp_ready; // @[Core.scala 114:23]
  assign io_core_bus_2_req_valid = icache_io_out_uncache_req_valid; // @[Core.scala 22:25]
  assign io_core_bus_2_req_bits_addr = icache_io_out_uncache_req_bits_addr; // @[Core.scala 22:25]
  assign io_core_bus_2_req_bits_size = icache_io_out_uncache_req_bits_size; // @[Core.scala 22:25]
  assign io_core_bus_2_resp_ready = icache_io_out_uncache_resp_ready; // @[Core.scala 22:25]
  assign io_core_bus_3_req_valid = dcache_io_out_uncache_req_valid; // @[Core.scala 115:25]
  assign io_core_bus_3_req_bits_addr = dcache_io_out_uncache_req_bits_addr; // @[Core.scala 115:25]
  assign io_core_bus_3_req_bits_wdata = dcache_io_out_uncache_req_bits_wdata; // @[Core.scala 115:25]
  assign io_core_bus_3_req_bits_wmask = dcache_io_out_uncache_req_bits_wmask; // @[Core.scala 115:25]
  assign io_core_bus_3_req_bits_wen = dcache_io_out_uncache_req_bits_wen; // @[Core.scala 115:25]
  assign io_core_bus_3_req_bits_size = dcache_io_out_uncache_req_bits_size; // @[Core.scala 115:25]
  assign io_core_bus_3_resp_ready = dcache_io_out_uncache_resp_ready; // @[Core.scala 115:25]
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_io_imem_req_ready = icache_io_in_req_ready; // @[Core.scala 20:16]
  assign fetch_io_imem_resp_valid = icache_io_in_resp_valid; // @[Core.scala 20:16]
  assign fetch_io_imem_resp_bits_rdata = icache_io_in_resp_bits_rdata; // @[Core.scala 20:16]
  assign fetch_io_imem_resp_bits_user = icache_io_in_resp_bits_user; // @[Core.scala 20:16]
  assign fetch_io_jmp_packet_valid = rob_io_jmp_packet_valid; // @[Core.scala 56:23]
  assign fetch_io_jmp_packet_inst_pc = rob_io_jmp_packet_inst_pc; // @[Core.scala 56:23]
  assign fetch_io_jmp_packet_jmp = rob_io_jmp_packet_jmp; // @[Core.scala 56:23]
  assign fetch_io_jmp_packet_jmp_pc = rob_io_jmp_packet_jmp_pc; // @[Core.scala 56:23]
  assign fetch_io_jmp_packet_mis = rob_io_jmp_packet_mis; // @[Core.scala 56:23]
  assign fetch_io_jmp_packet_sys = rob_io_jmp_packet_sys; // @[Core.scala 56:23]
  assign fetch_io_out_ready = ibuf_io_in_ready; // @[Core.scala 27:14]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_in_req_valid = fetch_io_imem_req_valid; // @[Core.scala 20:16]
  assign icache_io_in_req_bits_addr = fetch_io_imem_req_bits_addr; // @[Core.scala 20:16]
  assign icache_io_in_req_bits_user = fetch_io_imem_req_bits_user; // @[Core.scala 20:16]
  assign icache_io_in_resp_ready = fetch_io_imem_resp_ready; // @[Core.scala 20:16]
  assign icache_io_out_cache_req_ready = io_core_bus_0_req_ready; // @[Core.scala 21:23]
  assign icache_io_out_cache_resp_valid = io_core_bus_0_resp_valid; // @[Core.scala 21:23]
  assign icache_io_out_cache_resp_bits_rdata = io_core_bus_0_resp_bits_rdata; // @[Core.scala 21:23]
  assign icache_io_out_cache_resp_bits_rlast = io_core_bus_0_resp_bits_rlast; // @[Core.scala 21:23]
  assign icache_io_out_uncache_req_ready = io_core_bus_2_req_ready; // @[Core.scala 22:25]
  assign icache_io_out_uncache_resp_valid = io_core_bus_2_resp_valid; // @[Core.scala 22:25]
  assign icache_io_out_uncache_resp_bits_rdata = io_core_bus_2_resp_bits_rdata; // @[Core.scala 22:25]
  assign icache_fence_i = execution_fence_i;
  assign icache__WIRE_10 = dcache__WIRE_10;
  assign icache_empty = sq_empty_0;
  assign ibuf_clock = clock;
  assign ibuf_reset = reset;
  assign ibuf_io_in_valid = fetch_io_out_valid; // @[Core.scala 27:14]
  assign ibuf_io_in_bits_vec_0_pc = fetch_io_out_bits_vec_0_pc; // @[Core.scala 27:14]
  assign ibuf_io_in_bits_vec_0_inst = fetch_io_out_bits_vec_0_inst; // @[Core.scala 27:14]
  assign ibuf_io_in_bits_vec_0_pred_br = fetch_io_out_bits_vec_0_pred_br; // @[Core.scala 27:14]
  assign ibuf_io_in_bits_vec_0_pred_bpc = fetch_io_out_bits_vec_0_pred_bpc; // @[Core.scala 27:14]
  assign ibuf_io_in_bits_vec_0_valid = fetch_io_out_bits_vec_0_valid; // @[Core.scala 27:14]
  assign ibuf_io_in_bits_vec_1_pc = fetch_io_out_bits_vec_1_pc; // @[Core.scala 27:14]
  assign ibuf_io_in_bits_vec_1_inst = fetch_io_out_bits_vec_1_inst; // @[Core.scala 27:14]
  assign ibuf_io_in_bits_vec_1_pred_br = fetch_io_out_bits_vec_1_pred_br; // @[Core.scala 27:14]
  assign ibuf_io_in_bits_vec_1_pred_bpc = fetch_io_out_bits_vec_1_pred_bpc; // @[Core.scala 27:14]
  assign ibuf_io_in_bits_vec_1_valid = fetch_io_out_bits_vec_1_valid; // @[Core.scala 27:14]
  assign ibuf_io_out_ready = decode_io_in_ready; // @[Core.scala 33:16]
  assign ibuf_io_flush = rob_io_jmp_packet_mis; // @[Core.scala 28:17]
  assign decode_clock = clock;
  assign decode_reset = reset;
  assign decode_io_in_valid = ibuf_io_out_valid; // @[Core.scala 33:16]
  assign decode_io_in_bits_vec_0_pc = ibuf_io_out_bits_vec_0_pc; // @[Core.scala 33:16]
  assign decode_io_in_bits_vec_0_inst = ibuf_io_out_bits_vec_0_inst; // @[Core.scala 33:16]
  assign decode_io_in_bits_vec_0_pred_br = ibuf_io_out_bits_vec_0_pred_br; // @[Core.scala 33:16]
  assign decode_io_in_bits_vec_0_pred_bpc = ibuf_io_out_bits_vec_0_pred_bpc; // @[Core.scala 33:16]
  assign decode_io_in_bits_vec_0_valid = ibuf_io_out_bits_vec_0_valid; // @[Core.scala 33:16]
  assign decode_io_in_bits_vec_1_pc = ibuf_io_out_bits_vec_1_pc; // @[Core.scala 33:16]
  assign decode_io_in_bits_vec_1_inst = ibuf_io_out_bits_vec_1_inst; // @[Core.scala 33:16]
  assign decode_io_in_bits_vec_1_pred_br = ibuf_io_out_bits_vec_1_pred_br; // @[Core.scala 33:16]
  assign decode_io_in_bits_vec_1_pred_bpc = ibuf_io_out_bits_vec_1_pred_bpc; // @[Core.scala 33:16]
  assign decode_io_in_bits_vec_1_valid = ibuf_io_out_bits_vec_1_valid; // @[Core.scala 33:16]
  assign decode_io_out_ready = rename_io_in_ready; // @[Core.scala 37:16]
  assign decode_io_flush = rob_io_jmp_packet_mis; // @[Core.scala 34:19]
  assign rename_clock = clock;
  assign rename_reset = reset;
  assign rename_io_in_valid = decode_io_out_valid; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_valid = decode_io_out_bits_vec_0_valid; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_pc = decode_io_out_bits_vec_0_pc; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_npc = decode_io_out_bits_vec_0_npc; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_inst = decode_io_out_bits_vec_0_inst; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_fu_code = decode_io_out_bits_vec_0_fu_code; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_alu_code = decode_io_out_bits_vec_0_alu_code; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_jmp_code = decode_io_out_bits_vec_0_jmp_code; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_mem_code = decode_io_out_bits_vec_0_mem_code; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_mem_size = decode_io_out_bits_vec_0_mem_size; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_sys_code = decode_io_out_bits_vec_0_sys_code; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_w_type = decode_io_out_bits_vec_0_w_type; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_rs1_src = decode_io_out_bits_vec_0_rs1_src; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_rs2_src = decode_io_out_bits_vec_0_rs2_src; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_rs1_addr = decode_io_out_bits_vec_0_rs1_addr; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_rs2_addr = decode_io_out_bits_vec_0_rs2_addr; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_rd_addr = decode_io_out_bits_vec_0_rd_addr; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_rd_en = decode_io_out_bits_vec_0_rd_en; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_imm = decode_io_out_bits_vec_0_imm; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_pred_br = decode_io_out_bits_vec_0_pred_br; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_0_pred_bpc = decode_io_out_bits_vec_0_pred_bpc; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_valid = decode_io_out_bits_vec_1_valid; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_pc = decode_io_out_bits_vec_1_pc; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_npc = decode_io_out_bits_vec_1_npc; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_inst = decode_io_out_bits_vec_1_inst; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_fu_code = decode_io_out_bits_vec_1_fu_code; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_alu_code = decode_io_out_bits_vec_1_alu_code; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_jmp_code = decode_io_out_bits_vec_1_jmp_code; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_mem_code = decode_io_out_bits_vec_1_mem_code; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_mem_size = decode_io_out_bits_vec_1_mem_size; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_sys_code = decode_io_out_bits_vec_1_sys_code; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_w_type = decode_io_out_bits_vec_1_w_type; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_rs1_src = decode_io_out_bits_vec_1_rs1_src; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_rs2_src = decode_io_out_bits_vec_1_rs2_src; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_rs1_addr = decode_io_out_bits_vec_1_rs1_addr; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_rs2_addr = decode_io_out_bits_vec_1_rs2_addr; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_rd_addr = decode_io_out_bits_vec_1_rd_addr; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_rd_en = decode_io_out_bits_vec_1_rd_en; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_imm = decode_io_out_bits_vec_1_imm; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_pred_br = decode_io_out_bits_vec_1_pred_br; // @[Core.scala 37:16]
  assign rename_io_in_bits_vec_1_pred_bpc = decode_io_out_bits_vec_1_pred_bpc; // @[Core.scala 37:16]
  assign rename_io_out_ready = stall_reg_io_in_ready; // @[Core.scala 43:19]
  assign rename_io_flush = rob_io_jmp_packet_mis; // @[Core.scala 38:19]
  assign rename_io_exe_0_valid = isu_io_out_0_valid; // @[Core.scala 84:24]
  assign rename_io_exe_0_rd_en = isu_io_out_0_rd_en; // @[Core.scala 84:24]
  assign rename_io_exe_0_rd_paddr = isu_io_out_0_rd_paddr; // @[Core.scala 84:24]
  assign rename_io_exe_1_valid = isu_io_out_1_valid; // @[Core.scala 84:24]
  assign rename_io_exe_1_rd_en = isu_io_out_1_rd_en; // @[Core.scala 84:24]
  assign rename_io_exe_1_rd_paddr = isu_io_out_1_rd_paddr; // @[Core.scala 84:24]
  assign rename_io_exe_2_valid = execution_io_lsu_wakeup_uop_valid; // @[Core.scala 86:24]
  assign rename_io_exe_2_rd_en = execution_io_lsu_wakeup_uop_rd_en; // @[Core.scala 86:24]
  assign rename_io_exe_2_rd_paddr = execution_io_lsu_wakeup_uop_rd_paddr; // @[Core.scala 86:24]
  assign rename_io_cm_recover = REG; // @[Core.scala 53:24]
  assign rename_io_cm_0_valid = rob_io_cm_0_valid; // @[Core.scala 54:16]
  assign rename_io_cm_0_rd_addr = rob_io_cm_0_rd_addr; // @[Core.scala 54:16]
  assign rename_io_cm_0_rd_en = rob_io_cm_0_rd_en; // @[Core.scala 54:16]
  assign rename_io_cm_0_rd_paddr = rob_io_cm_0_rd_paddr; // @[Core.scala 54:16]
  assign rename_io_cm_0_rd_ppaddr = rob_io_cm_0_rd_ppaddr; // @[Core.scala 54:16]
  assign rename_io_cm_1_valid = rob_io_cm_1_valid; // @[Core.scala 54:16]
  assign rename_io_cm_1_rd_addr = rob_io_cm_1_rd_addr; // @[Core.scala 54:16]
  assign rename_io_cm_1_rd_en = rob_io_cm_1_rd_en; // @[Core.scala 54:16]
  assign rename_io_cm_1_rd_paddr = rob_io_cm_1_rd_paddr; // @[Core.scala 54:16]
  assign rename_io_cm_1_rd_ppaddr = rob_io_cm_1_rd_ppaddr; // @[Core.scala 54:16]
  assign stall_reg_clock = clock;
  assign stall_reg_reset = reset;
  assign stall_reg_io_flush = rob_io_jmp_packet_mis; // @[Core.scala 44:22]
  assign stall_reg_io_in_valid = rename_io_out_valid; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_valid = rename_io_out_bits_vec_0_valid; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_pc = rename_io_out_bits_vec_0_pc; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_npc = rename_io_out_bits_vec_0_npc; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_inst = rename_io_out_bits_vec_0_inst; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_fu_code = rename_io_out_bits_vec_0_fu_code; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_alu_code = rename_io_out_bits_vec_0_alu_code; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_jmp_code = rename_io_out_bits_vec_0_jmp_code; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_mem_code = rename_io_out_bits_vec_0_mem_code; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_mem_size = rename_io_out_bits_vec_0_mem_size; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_sys_code = rename_io_out_bits_vec_0_sys_code; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_w_type = rename_io_out_bits_vec_0_w_type; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_rs1_src = rename_io_out_bits_vec_0_rs1_src; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_rs2_src = rename_io_out_bits_vec_0_rs2_src; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_rd_addr = rename_io_out_bits_vec_0_rd_addr; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_rd_en = rename_io_out_bits_vec_0_rd_en; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_imm = rename_io_out_bits_vec_0_imm; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_pred_br = rename_io_out_bits_vec_0_pred_br; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_pred_bpc = rename_io_out_bits_vec_0_pred_bpc; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_rs1_paddr = rename_io_out_bits_vec_0_rs1_paddr; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_rs2_paddr = rename_io_out_bits_vec_0_rs2_paddr; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_rd_paddr = rename_io_out_bits_vec_0_rd_paddr; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_0_rd_ppaddr = rename_io_out_bits_vec_0_rd_ppaddr; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_valid = rename_io_out_bits_vec_1_valid; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_pc = rename_io_out_bits_vec_1_pc; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_npc = rename_io_out_bits_vec_1_npc; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_inst = rename_io_out_bits_vec_1_inst; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_fu_code = rename_io_out_bits_vec_1_fu_code; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_alu_code = rename_io_out_bits_vec_1_alu_code; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_jmp_code = rename_io_out_bits_vec_1_jmp_code; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_mem_code = rename_io_out_bits_vec_1_mem_code; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_mem_size = rename_io_out_bits_vec_1_mem_size; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_sys_code = rename_io_out_bits_vec_1_sys_code; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_w_type = rename_io_out_bits_vec_1_w_type; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_rs1_src = rename_io_out_bits_vec_1_rs1_src; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_rs2_src = rename_io_out_bits_vec_1_rs2_src; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_rd_addr = rename_io_out_bits_vec_1_rd_addr; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_rd_en = rename_io_out_bits_vec_1_rd_en; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_imm = rename_io_out_bits_vec_1_imm; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_pred_br = rename_io_out_bits_vec_1_pred_br; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_pred_bpc = rename_io_out_bits_vec_1_pred_bpc; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_rs1_paddr = rename_io_out_bits_vec_1_rs1_paddr; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_rs2_paddr = rename_io_out_bits_vec_1_rs2_paddr; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_rd_paddr = rename_io_out_bits_vec_1_rd_paddr; // @[Core.scala 43:19]
  assign stall_reg_io_in_bits_vec_1_rd_ppaddr = rename_io_out_bits_vec_1_rd_ppaddr; // @[Core.scala 43:19]
  assign stall_reg_io_out_ready = rob_io_in_ready & isu_io_in_ready; // @[Core.scala 66:45]
  assign rob_clock = clock;
  assign rob_reset = reset;
  assign rob_io_in_valid = stall_reg_io_out_valid & isu_io_in_ready; // @[Core.scala 50:45]
  assign rob_io_in_bits_vec_0_valid = stall_reg_io_out_bits_vec_0_valid; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_0_pc = stall_reg_io_out_bits_vec_0_pc; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_0_fu_code = stall_reg_io_out_bits_vec_0_fu_code; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_0_sys_code = stall_reg_io_out_bits_vec_0_sys_code; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_0_rd_addr = stall_reg_io_out_bits_vec_0_rd_addr; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_0_rd_en = stall_reg_io_out_bits_vec_0_rd_en; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_0_rd_paddr = stall_reg_io_out_bits_vec_0_rd_paddr; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_0_rd_ppaddr = stall_reg_io_out_bits_vec_0_rd_ppaddr; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_1_valid = stall_reg_io_out_bits_vec_1_valid; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_1_pc = stall_reg_io_out_bits_vec_1_pc; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_1_fu_code = stall_reg_io_out_bits_vec_1_fu_code; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_1_sys_code = stall_reg_io_out_bits_vec_1_sys_code; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_1_rd_addr = stall_reg_io_out_bits_vec_1_rd_addr; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_1_rd_en = stall_reg_io_out_bits_vec_1_rd_en; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_1_rd_paddr = stall_reg_io_out_bits_vec_1_rd_paddr; // @[Core.scala 49:18]
  assign rob_io_in_bits_vec_1_rd_ppaddr = stall_reg_io_out_bits_vec_1_rd_ppaddr; // @[Core.scala 49:18]
  assign rob_io_exe_0_valid = execution_io_out_0_valid; // @[Core.scala 90:14]
  assign rob_io_exe_0_rob_addr = execution_io_out_0_rob_addr; // @[Core.scala 90:14]
  assign rob_io_exe_1_valid = execution_io_out_1_valid; // @[Core.scala 90:14]
  assign rob_io_exe_1_rob_addr = execution_io_out_1_rob_addr; // @[Core.scala 90:14]
  assign rob_io_exe_2_valid = execution_io_out_2_valid; // @[Core.scala 90:14]
  assign rob_io_exe_2_rob_addr = execution_io_out_2_rob_addr; // @[Core.scala 90:14]
  assign rob_io_exe_ecp_0_jmp_valid = execution_io_out_ecp_0_jmp_valid; // @[Core.scala 91:18]
  assign rob_io_exe_ecp_0_jmp = execution_io_out_ecp_0_jmp; // @[Core.scala 91:18]
  assign rob_io_exe_ecp_0_jmp_pc = execution_io_out_ecp_0_jmp_pc; // @[Core.scala 91:18]
  assign rob_io_exe_ecp_0_mis = execution_io_out_ecp_0_mis; // @[Core.scala 91:18]
  assign rob_io_exe_ecp_1_jmp_valid = execution_io_out_ecp_1_jmp_valid; // @[Core.scala 91:18]
  assign rob_io_exe_ecp_1_jmp = execution_io_out_ecp_1_jmp; // @[Core.scala 91:18]
  assign rob_io_exe_ecp_1_jmp_pc = execution_io_out_ecp_1_jmp_pc; // @[Core.scala 91:18]
  assign rob_io_exe_ecp_1_mis = execution_io_out_ecp_1_mis; // @[Core.scala 91:18]
  assign rob_io_exe_ecp_2_store_valid = execution_io_out_ecp_2_store_valid; // @[Core.scala 91:18]
  assign rob_io_flush = rob_io_jmp_packet_mis; // @[Core.scala 51:16]
  assign rob_csr_mip_mtip_intr_0 = execution_mtip;
  assign rob_csr_mtvec_idx_0 = execution__T_6_0;
  assign rob_csr_mie_mtie_0 = execution__T_5_0;
  assign rob_csr_mstatus_0 = execution_mstatus;
  assign isu_clock = clock;
  assign isu_reset = reset;
  assign isu_io_flush = rob_io_jmp_packet_mis; // @[Core.scala 62:16]
  assign isu_io_in_valid = stall_reg_io_out_valid & rob_io_in_ready; // @[Core.scala 60:45]
  assign isu_io_in_bits_vec_0_valid = stall_reg_io_out_bits_vec_0_valid; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_pc = stall_reg_io_out_bits_vec_0_pc; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_npc = stall_reg_io_out_bits_vec_0_npc; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_inst = stall_reg_io_out_bits_vec_0_inst; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_fu_code = stall_reg_io_out_bits_vec_0_fu_code; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_alu_code = stall_reg_io_out_bits_vec_0_alu_code; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_jmp_code = stall_reg_io_out_bits_vec_0_jmp_code; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_mem_code = stall_reg_io_out_bits_vec_0_mem_code; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_mem_size = stall_reg_io_out_bits_vec_0_mem_size; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_sys_code = stall_reg_io_out_bits_vec_0_sys_code; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_w_type = stall_reg_io_out_bits_vec_0_w_type; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_rs1_src = stall_reg_io_out_bits_vec_0_rs1_src; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_rs2_src = stall_reg_io_out_bits_vec_0_rs2_src; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_rd_en = stall_reg_io_out_bits_vec_0_rd_en; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_imm = stall_reg_io_out_bits_vec_0_imm; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_pred_br = stall_reg_io_out_bits_vec_0_pred_br; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_pred_bpc = stall_reg_io_out_bits_vec_0_pred_bpc; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_rs1_paddr = stall_reg_io_out_bits_vec_0_rs1_paddr; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_rs2_paddr = stall_reg_io_out_bits_vec_0_rs2_paddr; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_0_rd_paddr = stall_reg_io_out_bits_vec_0_rd_paddr; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_valid = stall_reg_io_out_bits_vec_1_valid; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_pc = stall_reg_io_out_bits_vec_1_pc; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_npc = stall_reg_io_out_bits_vec_1_npc; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_inst = stall_reg_io_out_bits_vec_1_inst; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_fu_code = stall_reg_io_out_bits_vec_1_fu_code; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_alu_code = stall_reg_io_out_bits_vec_1_alu_code; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_jmp_code = stall_reg_io_out_bits_vec_1_jmp_code; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_mem_code = stall_reg_io_out_bits_vec_1_mem_code; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_mem_size = stall_reg_io_out_bits_vec_1_mem_size; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_sys_code = stall_reg_io_out_bits_vec_1_sys_code; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_w_type = stall_reg_io_out_bits_vec_1_w_type; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_rs1_src = stall_reg_io_out_bits_vec_1_rs1_src; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_rs2_src = stall_reg_io_out_bits_vec_1_rs2_src; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_rd_en = stall_reg_io_out_bits_vec_1_rd_en; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_imm = stall_reg_io_out_bits_vec_1_imm; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_pred_br = stall_reg_io_out_bits_vec_1_pred_br; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_pred_bpc = stall_reg_io_out_bits_vec_1_pred_bpc; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_rs1_paddr = stall_reg_io_out_bits_vec_1_rs1_paddr; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_rs2_paddr = stall_reg_io_out_bits_vec_1_rs2_paddr; // @[Core.scala 59:18]
  assign isu_io_in_bits_vec_1_rd_paddr = stall_reg_io_out_bits_vec_1_rd_paddr; // @[Core.scala 59:18]
  assign isu_io_rob_addr_0 = rob_io_rob_addr_0; // @[Core.scala 61:19]
  assign isu_io_rob_addr_1 = rob_io_rob_addr_1; // @[Core.scala 61:19]
  assign isu_io_avail_list = rename_io_avail_list; // @[Core.scala 63:21]
  assign isu_io_lsu_ready = execution_io_lsu_ready; // @[Core.scala 93:20]
  assign isu_io_sys_ready = rob_io_sys_ready; // @[Core.scala 64:20]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_in_0_valid = isu_io_out_0_valid; // @[Core.scala 71:12]
  assign rf_io_in_0_pc = isu_io_out_0_pc; // @[Core.scala 71:12]
  assign rf_io_in_0_npc = isu_io_out_0_npc; // @[Core.scala 71:12]
  assign rf_io_in_0_inst = isu_io_out_0_inst; // @[Core.scala 71:12]
  assign rf_io_in_0_fu_code = isu_io_out_0_fu_code; // @[Core.scala 71:12]
  assign rf_io_in_0_alu_code = isu_io_out_0_alu_code; // @[Core.scala 71:12]
  assign rf_io_in_0_jmp_code = isu_io_out_0_jmp_code; // @[Core.scala 71:12]
  assign rf_io_in_0_sys_code = isu_io_out_0_sys_code; // @[Core.scala 71:12]
  assign rf_io_in_0_w_type = isu_io_out_0_w_type; // @[Core.scala 71:12]
  assign rf_io_in_0_rs1_src = isu_io_out_0_rs1_src; // @[Core.scala 71:12]
  assign rf_io_in_0_rs2_src = isu_io_out_0_rs2_src; // @[Core.scala 71:12]
  assign rf_io_in_0_rd_en = isu_io_out_0_rd_en; // @[Core.scala 71:12]
  assign rf_io_in_0_imm = isu_io_out_0_imm; // @[Core.scala 71:12]
  assign rf_io_in_0_pred_br = isu_io_out_0_pred_br; // @[Core.scala 71:12]
  assign rf_io_in_0_pred_bpc = isu_io_out_0_pred_bpc; // @[Core.scala 71:12]
  assign rf_io_in_0_rs1_paddr = isu_io_out_0_rs1_paddr; // @[Core.scala 71:12]
  assign rf_io_in_0_rs2_paddr = isu_io_out_0_rs2_paddr; // @[Core.scala 71:12]
  assign rf_io_in_0_rd_paddr = isu_io_out_0_rd_paddr; // @[Core.scala 71:12]
  assign rf_io_in_0_rob_addr = isu_io_out_0_rob_addr; // @[Core.scala 71:12]
  assign rf_io_in_1_valid = isu_io_out_1_valid; // @[Core.scala 71:12]
  assign rf_io_in_1_pc = isu_io_out_1_pc; // @[Core.scala 71:12]
  assign rf_io_in_1_npc = isu_io_out_1_npc; // @[Core.scala 71:12]
  assign rf_io_in_1_fu_code = isu_io_out_1_fu_code; // @[Core.scala 71:12]
  assign rf_io_in_1_alu_code = isu_io_out_1_alu_code; // @[Core.scala 71:12]
  assign rf_io_in_1_jmp_code = isu_io_out_1_jmp_code; // @[Core.scala 71:12]
  assign rf_io_in_1_w_type = isu_io_out_1_w_type; // @[Core.scala 71:12]
  assign rf_io_in_1_rs1_src = isu_io_out_1_rs1_src; // @[Core.scala 71:12]
  assign rf_io_in_1_rs2_src = isu_io_out_1_rs2_src; // @[Core.scala 71:12]
  assign rf_io_in_1_rd_en = isu_io_out_1_rd_en; // @[Core.scala 71:12]
  assign rf_io_in_1_imm = isu_io_out_1_imm; // @[Core.scala 71:12]
  assign rf_io_in_1_pred_br = isu_io_out_1_pred_br; // @[Core.scala 71:12]
  assign rf_io_in_1_pred_bpc = isu_io_out_1_pred_bpc; // @[Core.scala 71:12]
  assign rf_io_in_1_rs1_paddr = isu_io_out_1_rs1_paddr; // @[Core.scala 71:12]
  assign rf_io_in_1_rs2_paddr = isu_io_out_1_rs2_paddr; // @[Core.scala 71:12]
  assign rf_io_in_1_rd_paddr = isu_io_out_1_rd_paddr; // @[Core.scala 71:12]
  assign rf_io_in_1_rob_addr = isu_io_out_1_rob_addr; // @[Core.scala 71:12]
  assign rf_io_in_2_valid = isu_io_out_2_valid; // @[Core.scala 71:12]
  assign rf_io_in_2_pc = isu_io_out_2_pc; // @[Core.scala 71:12]
  assign rf_io_in_2_fu_code = isu_io_out_2_fu_code; // @[Core.scala 71:12]
  assign rf_io_in_2_alu_code = isu_io_out_2_alu_code; // @[Core.scala 71:12]
  assign rf_io_in_2_mem_code = isu_io_out_2_mem_code; // @[Core.scala 71:12]
  assign rf_io_in_2_mem_size = isu_io_out_2_mem_size; // @[Core.scala 71:12]
  assign rf_io_in_2_w_type = isu_io_out_2_w_type; // @[Core.scala 71:12]
  assign rf_io_in_2_rs1_src = isu_io_out_2_rs1_src; // @[Core.scala 71:12]
  assign rf_io_in_2_rs2_src = isu_io_out_2_rs2_src; // @[Core.scala 71:12]
  assign rf_io_in_2_rd_en = isu_io_out_2_rd_en; // @[Core.scala 71:12]
  assign rf_io_in_2_imm = isu_io_out_2_imm; // @[Core.scala 71:12]
  assign rf_io_in_2_rs1_paddr = isu_io_out_2_rs1_paddr; // @[Core.scala 71:12]
  assign rf_io_in_2_rs2_paddr = isu_io_out_2_rs2_paddr; // @[Core.scala 71:12]
  assign rf_io_in_2_rd_paddr = isu_io_out_2_rd_paddr; // @[Core.scala 71:12]
  assign rf_io_in_2_rob_addr = isu_io_out_2_rob_addr; // @[Core.scala 71:12]
  assign rf_io_rd_en_0 = execution_io_rd_en_0; // @[Core.scala 122:15]
  assign rf_io_rd_en_1 = execution_io_rd_en_1; // @[Core.scala 122:15]
  assign rf_io_rd_en_2 = execution_io_rd_en_2; // @[Core.scala 122:15]
  assign rf_io_rd_paddr_0 = execution_io_rd_paddr_0; // @[Core.scala 123:18]
  assign rf_io_rd_paddr_1 = execution_io_rd_paddr_1; // @[Core.scala 123:18]
  assign rf_io_rd_paddr_2 = execution_io_rd_paddr_2; // @[Core.scala 123:18]
  assign rf_io_rd_data_0 = execution_io_rd_data_0; // @[Core.scala 124:17]
  assign rf_io_rd_data_1 = execution_io_rd_data_1; // @[Core.scala 124:17]
  assign rf_io_rd_data_2 = execution_io_rd_data_2; // @[Core.scala 124:17]
  assign rf_io_flush = rob_io_jmp_packet_mis; // @[Core.scala 72:15]
  assign execution_clock = clock;
  assign execution_reset = reset;
  assign execution_io_in_0_valid = rf_io_out_0_valid; // @[Core.scala 77:19]
  assign execution_io_in_0_pc = rf_io_out_0_pc; // @[Core.scala 77:19]
  assign execution_io_in_0_npc = rf_io_out_0_npc; // @[Core.scala 77:19]
  assign execution_io_in_0_inst = rf_io_out_0_inst; // @[Core.scala 77:19]
  assign execution_io_in_0_fu_code = rf_io_out_0_fu_code; // @[Core.scala 77:19]
  assign execution_io_in_0_alu_code = rf_io_out_0_alu_code; // @[Core.scala 77:19]
  assign execution_io_in_0_jmp_code = rf_io_out_0_jmp_code; // @[Core.scala 77:19]
  assign execution_io_in_0_sys_code = rf_io_out_0_sys_code; // @[Core.scala 77:19]
  assign execution_io_in_0_w_type = rf_io_out_0_w_type; // @[Core.scala 77:19]
  assign execution_io_in_0_rs1_src = rf_io_out_0_rs1_src; // @[Core.scala 77:19]
  assign execution_io_in_0_rs2_src = rf_io_out_0_rs2_src; // @[Core.scala 77:19]
  assign execution_io_in_0_rd_en = rf_io_out_0_rd_en; // @[Core.scala 77:19]
  assign execution_io_in_0_imm = rf_io_out_0_imm; // @[Core.scala 77:19]
  assign execution_io_in_0_pred_br = rf_io_out_0_pred_br; // @[Core.scala 77:19]
  assign execution_io_in_0_pred_bpc = rf_io_out_0_pred_bpc; // @[Core.scala 77:19]
  assign execution_io_in_0_rd_paddr = rf_io_out_0_rd_paddr; // @[Core.scala 77:19]
  assign execution_io_in_0_rob_addr = rf_io_out_0_rob_addr; // @[Core.scala 77:19]
  assign execution_io_in_1_valid = rf_io_out_1_valid; // @[Core.scala 77:19]
  assign execution_io_in_1_pc = rf_io_out_1_pc; // @[Core.scala 77:19]
  assign execution_io_in_1_npc = rf_io_out_1_npc; // @[Core.scala 77:19]
  assign execution_io_in_1_fu_code = rf_io_out_1_fu_code; // @[Core.scala 77:19]
  assign execution_io_in_1_alu_code = rf_io_out_1_alu_code; // @[Core.scala 77:19]
  assign execution_io_in_1_jmp_code = rf_io_out_1_jmp_code; // @[Core.scala 77:19]
  assign execution_io_in_1_w_type = rf_io_out_1_w_type; // @[Core.scala 77:19]
  assign execution_io_in_1_rs1_src = rf_io_out_1_rs1_src; // @[Core.scala 77:19]
  assign execution_io_in_1_rs2_src = rf_io_out_1_rs2_src; // @[Core.scala 77:19]
  assign execution_io_in_1_rd_en = rf_io_out_1_rd_en; // @[Core.scala 77:19]
  assign execution_io_in_1_imm = rf_io_out_1_imm; // @[Core.scala 77:19]
  assign execution_io_in_1_pred_br = rf_io_out_1_pred_br; // @[Core.scala 77:19]
  assign execution_io_in_1_pred_bpc = rf_io_out_1_pred_bpc; // @[Core.scala 77:19]
  assign execution_io_in_1_rd_paddr = rf_io_out_1_rd_paddr; // @[Core.scala 77:19]
  assign execution_io_in_1_rob_addr = rf_io_out_1_rob_addr; // @[Core.scala 77:19]
  assign execution_io_in_2_valid = rf_io_out_2_valid; // @[Core.scala 77:19]
  assign execution_io_in_2_pc = rf_io_out_2_pc; // @[Core.scala 77:19]
  assign execution_io_in_2_fu_code = rf_io_out_2_fu_code; // @[Core.scala 77:19]
  assign execution_io_in_2_alu_code = rf_io_out_2_alu_code; // @[Core.scala 77:19]
  assign execution_io_in_2_mem_code = rf_io_out_2_mem_code; // @[Core.scala 77:19]
  assign execution_io_in_2_mem_size = rf_io_out_2_mem_size; // @[Core.scala 77:19]
  assign execution_io_in_2_w_type = rf_io_out_2_w_type; // @[Core.scala 77:19]
  assign execution_io_in_2_rs1_src = rf_io_out_2_rs1_src; // @[Core.scala 77:19]
  assign execution_io_in_2_rs2_src = rf_io_out_2_rs2_src; // @[Core.scala 77:19]
  assign execution_io_in_2_rd_en = rf_io_out_2_rd_en; // @[Core.scala 77:19]
  assign execution_io_in_2_imm = rf_io_out_2_imm; // @[Core.scala 77:19]
  assign execution_io_in_2_rd_paddr = rf_io_out_2_rd_paddr; // @[Core.scala 77:19]
  assign execution_io_in_2_rob_addr = rf_io_out_2_rob_addr; // @[Core.scala 77:19]
  assign execution_io_rs1_data_0 = rf_io_rs1_data_0; // @[Core.scala 79:25]
  assign execution_io_rs1_data_1 = rf_io_rs1_data_1; // @[Core.scala 79:25]
  assign execution_io_rs1_data_2 = rf_io_rs1_data_2; // @[Core.scala 79:25]
  assign execution_io_rs2_data_0 = rf_io_rs2_data_0; // @[Core.scala 80:25]
  assign execution_io_rs2_data_1 = rf_io_rs2_data_1; // @[Core.scala 80:25]
  assign execution_io_rs2_data_2 = rf_io_rs2_data_2; // @[Core.scala 80:25]
  assign execution_io_flush = rob_io_jmp_packet_mis; // @[Core.scala 78:22]
  assign execution_io_dmem_st_req_ready = sq_io_in_st_req_ready; // @[Core.scala 97:15]
  assign execution_io_dmem_st_resp_valid = sq_io_in_st_resp_valid; // @[Core.scala 97:15]
  assign execution_io_dmem_ld_req_ready = sq_io_in_ld_req_ready; // @[Core.scala 98:15]
  assign execution_io_dmem_ld_resp_valid = sq_io_in_ld_resp_valid; // @[Core.scala 98:15]
  assign execution_io_dmem_ld_resp_bits_rdata = sq_io_in_ld_resp_bits_rdata; // @[Core.scala 98:15]
  assign execution_intr_mcause = rob_intr_mcause_0;
  assign execution_instr_cnt = instr_cnt;
  assign execution_intr_mstatus = rob_intr_mstatus_0;
  assign execution_intr = rob_intr_0;
  assign execution_cycle_cnt = cycle_cnt;
  assign execution_intr_mepc = rob_intr_mepc_0;
  assign execution_mtip_0 = clint_mtip_1;
  assign sq_clock = clock;
  assign sq_reset = reset;
  assign sq_io_flush = rob_io_jmp_packet_mis; // @[Core.scala 96:15]
  assign sq_io_in_st_req_valid = execution_io_dmem_st_req_valid; // @[Core.scala 97:15]
  assign sq_io_in_st_req_bits_addr = execution_io_dmem_st_req_bits_addr; // @[Core.scala 97:15]
  assign sq_io_in_st_req_bits_wdata = execution_io_dmem_st_req_bits_wdata; // @[Core.scala 97:15]
  assign sq_io_in_st_req_bits_wmask = execution_io_dmem_st_req_bits_wmask; // @[Core.scala 97:15]
  assign sq_io_in_st_req_bits_size = execution_io_dmem_st_req_bits_size; // @[Core.scala 97:15]
  assign sq_io_in_st_resp_ready = execution_io_dmem_st_resp_ready; // @[Core.scala 97:15]
  assign sq_io_in_ld_req_valid = execution_io_dmem_ld_req_valid; // @[Core.scala 98:15]
  assign sq_io_in_ld_req_bits_addr = execution_io_dmem_ld_req_bits_addr; // @[Core.scala 98:15]
  assign sq_io_in_ld_req_bits_size = execution_io_dmem_ld_req_bits_size; // @[Core.scala 98:15]
  assign sq_io_in_ld_resp_ready = execution_io_dmem_ld_resp_ready; // @[Core.scala 98:15]
  assign sq_io_out_st_req_ready = crossbar2to1_io_in_0_req_ready; // @[Core.scala 102:25]
  assign sq_io_out_st_resp_valid = crossbar2to1_io_in_0_resp_valid; // @[Core.scala 102:25]
  assign sq_io_out_ld_req_ready = crossbar2to1_io_in_1_req_ready; // @[Core.scala 103:25]
  assign sq_io_out_ld_resp_valid = crossbar2to1_io_in_1_resp_valid; // @[Core.scala 103:25]
  assign sq_io_out_ld_resp_bits_rdata = crossbar2to1_io_in_1_resp_bits_rdata; // @[Core.scala 103:25]
  assign sq_io_deq_req = rob_io_sq_deq_req; // @[Core.scala 99:17]
  assign crossbar2to1_clock = clock;
  assign crossbar2to1_io_in_0_req_valid = sq_io_out_st_req_valid; // @[Core.scala 102:25]
  assign crossbar2to1_io_in_0_req_bits_addr = sq_io_out_st_req_bits_addr; // @[Core.scala 102:25]
  assign crossbar2to1_io_in_0_req_bits_wdata = sq_io_out_st_req_bits_wdata; // @[Core.scala 102:25]
  assign crossbar2to1_io_in_0_req_bits_wmask = sq_io_out_st_req_bits_wmask; // @[Core.scala 102:25]
  assign crossbar2to1_io_in_0_req_bits_size = sq_io_out_st_req_bits_size; // @[Core.scala 102:25]
  assign crossbar2to1_io_in_0_resp_ready = sq_io_out_st_resp_ready; // @[Core.scala 102:25]
  assign crossbar2to1_io_in_1_req_valid = sq_io_out_ld_req_valid; // @[Core.scala 103:25]
  assign crossbar2to1_io_in_1_req_bits_addr = sq_io_out_ld_req_bits_addr; // @[Core.scala 103:25]
  assign crossbar2to1_io_in_1_req_bits_size = sq_io_out_ld_req_bits_size; // @[Core.scala 103:25]
  assign crossbar2to1_io_in_1_resp_ready = sq_io_out_ld_resp_ready; // @[Core.scala 103:25]
  assign crossbar2to1_io_out_req_ready = crossbar1to2_io_in_req_ready; // @[Core.scala 106:22]
  assign crossbar2to1_io_out_resp_valid = crossbar1to2_io_in_resp_valid; // @[Core.scala 106:22]
  assign crossbar2to1_io_out_resp_bits_id = crossbar1to2_io_in_resp_bits_id; // @[Core.scala 106:22]
  assign crossbar2to1_io_out_resp_bits_rdata = crossbar1to2_io_in_resp_bits_rdata; // @[Core.scala 106:22]
  assign crossbar1to2_clock = clock;
  assign crossbar1to2_reset = reset;
  assign crossbar1to2_io_in_req_valid = crossbar2to1_io_out_req_valid; // @[Core.scala 106:22]
  assign crossbar1to2_io_in_req_bits_id = crossbar2to1_io_out_req_bits_id; // @[Core.scala 106:22]
  assign crossbar1to2_io_in_req_bits_addr = crossbar2to1_io_out_req_bits_addr; // @[Core.scala 106:22]
  assign crossbar1to2_io_in_req_bits_wdata = crossbar2to1_io_out_req_bits_wdata; // @[Core.scala 106:22]
  assign crossbar1to2_io_in_req_bits_wmask = crossbar2to1_io_out_req_bits_wmask; // @[Core.scala 106:22]
  assign crossbar1to2_io_in_req_bits_wen = crossbar2to1_io_out_req_bits_wen; // @[Core.scala 106:22]
  assign crossbar1to2_io_in_req_bits_size = crossbar2to1_io_out_req_bits_size; // @[Core.scala 106:22]
  assign crossbar1to2_io_in_resp_ready = crossbar2to1_io_out_resp_ready; // @[Core.scala 106:22]
  assign crossbar1to2_io_out_0_req_ready = dcache_io_in_req_ready; // @[Core.scala 113:16]
  assign crossbar1to2_io_out_0_resp_valid = dcache_io_in_resp_valid; // @[Core.scala 113:16]
  assign crossbar1to2_io_out_0_resp_bits_id = dcache_io_in_resp_bits_id; // @[Core.scala 113:16]
  assign crossbar1to2_io_out_0_resp_bits_rdata = dcache_io_in_resp_bits_rdata; // @[Core.scala 113:16]
  assign crossbar1to2_io_out_1_req_ready = clint_io_in_req_ready; // @[Core.scala 118:15]
  assign crossbar1to2_io_out_1_resp_valid = clint_io_in_resp_valid; // @[Core.scala 118:15]
  assign crossbar1to2_io_out_1_resp_bits_id = clint_io_in_resp_bits_id; // @[Core.scala 118:15]
  assign crossbar1to2_io_out_1_resp_bits_rdata = clint_io_in_resp_bits_rdata; // @[Core.scala 118:15]
  assign crossbar1to2_io_to_1 = crossbar1to2_io_in_req_bits_addr >= 32'h2000000 & crossbar1to2_io_in_req_bits_addr < 32'h2010000
    ; // @[Core.scala 109:57]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_in_req_valid = crossbar1to2_io_out_0_req_valid; // @[Core.scala 113:16]
  assign dcache_io_in_req_bits_id = crossbar1to2_io_out_0_req_bits_id; // @[Core.scala 113:16]
  assign dcache_io_in_req_bits_addr = crossbar1to2_io_out_0_req_bits_addr; // @[Core.scala 113:16]
  assign dcache_io_in_req_bits_wdata = crossbar1to2_io_out_0_req_bits_wdata; // @[Core.scala 113:16]
  assign dcache_io_in_req_bits_wmask = crossbar1to2_io_out_0_req_bits_wmask; // @[Core.scala 113:16]
  assign dcache_io_in_req_bits_wen = crossbar1to2_io_out_0_req_bits_wen; // @[Core.scala 113:16]
  assign dcache_io_in_req_bits_size = crossbar1to2_io_out_0_req_bits_size; // @[Core.scala 113:16]
  assign dcache_io_in_resp_ready = crossbar1to2_io_out_0_resp_ready; // @[Core.scala 113:16]
  assign dcache_io_out_cache_req_ready = io_core_bus_1_req_ready; // @[Core.scala 114:23]
  assign dcache_io_out_cache_resp_valid = io_core_bus_1_resp_valid; // @[Core.scala 114:23]
  assign dcache_io_out_cache_resp_bits_rdata = io_core_bus_1_resp_bits_rdata; // @[Core.scala 114:23]
  assign dcache_io_out_cache_resp_bits_rlast = io_core_bus_1_resp_bits_rlast; // @[Core.scala 114:23]
  assign dcache_io_out_uncache_req_ready = io_core_bus_3_req_ready; // @[Core.scala 115:25]
  assign dcache_io_out_uncache_resp_valid = io_core_bus_3_resp_valid; // @[Core.scala 115:25]
  assign dcache_io_out_uncache_resp_bits_rdata = io_core_bus_3_resp_bits_rdata; // @[Core.scala 115:25]
  assign dcache_fence_i = execution_fence_i;
  assign dcache_empty = sq_empty_0;
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io_in_req_valid = crossbar1to2_io_out_1_req_valid; // @[Core.scala 118:15]
  assign clint_io_in_req_bits_id = crossbar1to2_io_out_1_req_bits_id; // @[Core.scala 118:15]
  assign clint_io_in_req_bits_addr = crossbar1to2_io_out_1_req_bits_addr; // @[Core.scala 118:15]
  assign clint_io_in_req_bits_wdata = crossbar1to2_io_out_1_req_bits_wdata; // @[Core.scala 118:15]
  assign clint_io_in_req_bits_wmask = crossbar1to2_io_out_1_req_bits_wmask; // @[Core.scala 118:15]
  assign clint_io_in_req_bits_wen = crossbar1to2_io_out_1_req_bits_wen; // @[Core.scala 118:15]
  assign clint_io_in_resp_ready = crossbar1to2_io_out_1_resp_ready; // @[Core.scala 118:15]
  always @(posedge clock) begin
    REG <= rob_io_jmp_packet_mis; // @[Core.scala 53:34]
    if (reset) begin // @[Core.scala 132:26]
      cycle_cnt <= 64'h0; // @[Core.scala 132:26]
    end else begin
      cycle_cnt <= _T_8; // @[Core.scala 138:13]
    end
    if (reset) begin // @[Core.scala 133:26]
      instr_cnt <= 64'h0; // @[Core.scala 133:26]
    end else begin
      instr_cnt <= _T_12; // @[Core.scala 139:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  cycle_cnt = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  instr_cnt = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_RRArbiter_1(
  input         clock,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input         io_in_0_bits_aen,
  input  [63:0] io_in_0_bits_wdata,
  input         io_in_0_bits_wlast,
  input         io_in_0_bits_wen,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input         io_in_1_bits_aen,
  input  [63:0] io_in_1_bits_wdata,
  input         io_in_1_bits_wlast,
  input         io_in_1_bits_wen,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_addr,
  input  [1:0]  io_in_2_bits_size,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_addr,
  input  [63:0] io_in_3_bits_wdata,
  input  [7:0]  io_in_3_bits_wmask,
  input         io_in_3_bits_wen,
  input  [1:0]  io_in_3_bits_size,
  input         io_out_ready,
  output        io_out_valid,
  output [3:0]  io_out_bits_id,
  output [31:0] io_out_bits_addr,
  output        io_out_bits_aen,
  output [63:0] io_out_bits_wdata,
  output [7:0]  io_out_bits_wmask,
  output        io_out_bits_wlast,
  output        io_out_bits_wen,
  output [7:0]  io_out_bits_len,
  output [1:0]  io_out_bits_size,
  output [1:0]  io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_1 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:{16,16}]
  wire  _GEN_2 = 2'h2 == io_chosen ? io_in_2_valid : _GEN_1; // @[Arbiter.scala 41:{16,16}]
  wire [1:0] _GEN_6 = 2'h2 == io_chosen ? io_in_2_bits_size : 2'h3; // @[Arbiter.scala 42:{15,15}]
  wire [7:0] _GEN_10 = 2'h2 == io_chosen ? 8'h0 : 8'h1; // @[Arbiter.scala 42:{15,15}]
  wire  _GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_wen : io_in_0_bits_wen; // @[Arbiter.scala 42:{15,15}]
  wire  _GEN_14 = 2'h2 == io_chosen ? 1'h0 : _GEN_13; // @[Arbiter.scala 42:{15,15}]
  wire  _GEN_17 = 2'h1 == io_chosen ? io_in_1_bits_wlast : io_in_0_bits_wlast; // @[Arbiter.scala 42:{15,15}]
  wire [7:0] _GEN_22 = 2'h2 == io_chosen ? 8'h0 : 8'hff; // @[Arbiter.scala 42:{15,15}]
  wire [63:0] _GEN_25 = 2'h1 == io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[Arbiter.scala 42:{15,15}]
  wire [63:0] _GEN_26 = 2'h2 == io_chosen ? 64'h0 : _GEN_25; // @[Arbiter.scala 42:{15,15}]
  wire  _GEN_29 = 2'h1 == io_chosen ? io_in_1_bits_aen : io_in_0_bits_aen; // @[Arbiter.scala 42:{15,15}]
  wire [31:0] _GEN_33 = 2'h1 == io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:{15,15}]
  wire [31:0] _GEN_34 = 2'h2 == io_chosen ? io_in_2_bits_addr : _GEN_33; // @[Arbiter.scala 42:{15,15}]
  wire [3:0] _GEN_37 = 2'h1 == io_chosen ? 4'h2 : 4'h1; // @[Arbiter.scala 42:{15,15}]
  wire [3:0] _GEN_38 = 2'h2 == io_chosen ? 4'h3 : _GEN_37; // @[Arbiter.scala 42:{15,15}]
  wire  _ctrl_validMask_grantMask_lastGrant_T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg [1:0] lastGrant; // @[Reg.scala 15:16]
  wire  grantMask_1 = 2'h1 > lastGrant; // @[Arbiter.scala 67:49]
  wire  grantMask_2 = 2'h2 > lastGrant; // @[Arbiter.scala 67:49]
  wire  grantMask_3 = 2'h3 > lastGrant; // @[Arbiter.scala 67:49]
  wire  validMask_1 = io_in_1_valid & grantMask_1; // @[Arbiter.scala 68:75]
  wire  validMask_2 = io_in_2_valid & grantMask_2; // @[Arbiter.scala 68:75]
  wire  validMask_3 = io_in_3_valid & grantMask_3; // @[Arbiter.scala 68:75]
  wire [1:0] _GEN_41 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 77:{27,36}]
  wire [1:0] _GEN_42 = io_in_1_valid ? 2'h1 : _GEN_41; // @[Arbiter.scala 77:{27,36}]
  wire [1:0] _GEN_43 = io_in_0_valid ? 2'h0 : _GEN_42; // @[Arbiter.scala 77:{27,36}]
  wire [1:0] _GEN_44 = validMask_3 ? 2'h3 : _GEN_43; // @[Arbiter.scala 79:{25,34}]
  wire [1:0] _GEN_45 = validMask_2 ? 2'h2 : _GEN_44; // @[Arbiter.scala 79:{25,34}]
  assign io_out_valid = 2'h3 == io_chosen ? io_in_3_valid : _GEN_2; // @[Arbiter.scala 41:{16,16}]
  assign io_out_bits_id = 2'h3 == io_chosen ? 4'h4 : _GEN_38; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_addr = 2'h3 == io_chosen ? io_in_3_bits_addr : _GEN_34; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_aen = 2'h3 == io_chosen | (2'h2 == io_chosen | _GEN_29); // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wdata = 2'h3 == io_chosen ? io_in_3_bits_wdata : _GEN_26; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wmask = 2'h3 == io_chosen ? io_in_3_bits_wmask : _GEN_22; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wlast = 2'h3 == io_chosen | (2'h2 == io_chosen | _GEN_17); // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_wen = 2'h3 == io_chosen ? io_in_3_bits_wen : _GEN_14; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_len = 2'h3 == io_chosen ? 8'h0 : _GEN_10; // @[Arbiter.scala 42:{15,15}]
  assign io_out_bits_size = 2'h3 == io_chosen ? io_in_3_bits_size : _GEN_6; // @[Arbiter.scala 42:{15,15}]
  assign io_chosen = validMask_1 ? 2'h1 : _GEN_45; // @[Arbiter.scala 79:{25,34}]
  always @(posedge clock) begin
    if (_ctrl_validMask_grantMask_lastGrant_T) begin // @[Reg.scala 16:19]
      lastGrant <= io_chosen; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lastGrant = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_210128_CoreBusCrossbarNto1(
  input         clock,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [31:0] io_in_0_req_bits_addr,
  input         io_in_0_req_bits_aen,
  input  [63:0] io_in_0_req_bits_wdata,
  input         io_in_0_req_bits_wlast,
  input         io_in_0_req_bits_wen,
  input         io_in_0_resp_ready,
  output        io_in_0_resp_valid,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_0_resp_bits_rlast,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [31:0] io_in_1_req_bits_addr,
  input         io_in_1_req_bits_aen,
  input  [63:0] io_in_1_req_bits_wdata,
  input         io_in_1_req_bits_wlast,
  input         io_in_1_req_bits_wen,
  input         io_in_1_resp_ready,
  output        io_in_1_resp_valid,
  output [63:0] io_in_1_resp_bits_rdata,
  output        io_in_1_resp_bits_rlast,
  output        io_in_2_req_ready,
  input         io_in_2_req_valid,
  input  [31:0] io_in_2_req_bits_addr,
  input  [1:0]  io_in_2_req_bits_size,
  input         io_in_2_resp_ready,
  output        io_in_2_resp_valid,
  output [63:0] io_in_2_resp_bits_rdata,
  output        io_in_3_req_ready,
  input         io_in_3_req_valid,
  input  [31:0] io_in_3_req_bits_addr,
  input  [63:0] io_in_3_req_bits_wdata,
  input  [7:0]  io_in_3_req_bits_wmask,
  input         io_in_3_req_bits_wen,
  input  [1:0]  io_in_3_req_bits_size,
  input         io_in_3_resp_ready,
  output        io_in_3_resp_valid,
  output [63:0] io_in_3_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [3:0]  io_out_req_bits_id,
  output [31:0] io_out_req_bits_addr,
  output        io_out_req_bits_aen,
  output [63:0] io_out_req_bits_wdata,
  output [7:0]  io_out_req_bits_wmask,
  output        io_out_req_bits_wlast,
  output        io_out_req_bits_wen,
  output [7:0]  io_out_req_bits_len,
  output [1:0]  io_out_req_bits_size,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_id,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_out_resp_bits_rlast
);
  wire  arbiter_clock; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_0_valid; // @[Crossbar.scala 12:23]
  wire [31:0] arbiter_io_in_0_bits_addr; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_0_bits_aen; // @[Crossbar.scala 12:23]
  wire [63:0] arbiter_io_in_0_bits_wdata; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_0_bits_wlast; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_0_bits_wen; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_1_valid; // @[Crossbar.scala 12:23]
  wire [31:0] arbiter_io_in_1_bits_addr; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_1_bits_aen; // @[Crossbar.scala 12:23]
  wire [63:0] arbiter_io_in_1_bits_wdata; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_1_bits_wlast; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_1_bits_wen; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_2_valid; // @[Crossbar.scala 12:23]
  wire [31:0] arbiter_io_in_2_bits_addr; // @[Crossbar.scala 12:23]
  wire [1:0] arbiter_io_in_2_bits_size; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_3_valid; // @[Crossbar.scala 12:23]
  wire [31:0] arbiter_io_in_3_bits_addr; // @[Crossbar.scala 12:23]
  wire [63:0] arbiter_io_in_3_bits_wdata; // @[Crossbar.scala 12:23]
  wire [7:0] arbiter_io_in_3_bits_wmask; // @[Crossbar.scala 12:23]
  wire  arbiter_io_in_3_bits_wen; // @[Crossbar.scala 12:23]
  wire [1:0] arbiter_io_in_3_bits_size; // @[Crossbar.scala 12:23]
  wire  arbiter_io_out_ready; // @[Crossbar.scala 12:23]
  wire  arbiter_io_out_valid; // @[Crossbar.scala 12:23]
  wire [3:0] arbiter_io_out_bits_id; // @[Crossbar.scala 12:23]
  wire [31:0] arbiter_io_out_bits_addr; // @[Crossbar.scala 12:23]
  wire  arbiter_io_out_bits_aen; // @[Crossbar.scala 12:23]
  wire [63:0] arbiter_io_out_bits_wdata; // @[Crossbar.scala 12:23]
  wire [7:0] arbiter_io_out_bits_wmask; // @[Crossbar.scala 12:23]
  wire  arbiter_io_out_bits_wlast; // @[Crossbar.scala 12:23]
  wire  arbiter_io_out_bits_wen; // @[Crossbar.scala 12:23]
  wire [7:0] arbiter_io_out_bits_len; // @[Crossbar.scala 12:23]
  wire [1:0] arbiter_io_out_bits_size; // @[Crossbar.scala 12:23]
  wire [1:0] arbiter_io_chosen; // @[Crossbar.scala 12:23]
  wire  _GEN_0 = io_out_resp_bits_id == 4'h1 & io_in_0_resp_ready; // @[Crossbar.scala 32:23 35:46 36:25]
  wire  _GEN_2 = io_out_resp_bits_id == 4'h2 ? io_in_1_resp_ready : _GEN_0; // @[Crossbar.scala 35:46 36:25]
  wire  _GEN_4 = io_out_resp_bits_id == 4'h3 ? io_in_2_resp_ready : _GEN_2; // @[Crossbar.scala 35:46 36:25]
  ysyx_210128_RRArbiter_1 arbiter ( // @[Crossbar.scala 12:23]
    .clock(arbiter_clock),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_0_bits_addr(arbiter_io_in_0_bits_addr),
    .io_in_0_bits_aen(arbiter_io_in_0_bits_aen),
    .io_in_0_bits_wdata(arbiter_io_in_0_bits_wdata),
    .io_in_0_bits_wlast(arbiter_io_in_0_bits_wlast),
    .io_in_0_bits_wen(arbiter_io_in_0_bits_wen),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_1_bits_addr(arbiter_io_in_1_bits_addr),
    .io_in_1_bits_aen(arbiter_io_in_1_bits_aen),
    .io_in_1_bits_wdata(arbiter_io_in_1_bits_wdata),
    .io_in_1_bits_wlast(arbiter_io_in_1_bits_wlast),
    .io_in_1_bits_wen(arbiter_io_in_1_bits_wen),
    .io_in_2_valid(arbiter_io_in_2_valid),
    .io_in_2_bits_addr(arbiter_io_in_2_bits_addr),
    .io_in_2_bits_size(arbiter_io_in_2_bits_size),
    .io_in_3_valid(arbiter_io_in_3_valid),
    .io_in_3_bits_addr(arbiter_io_in_3_bits_addr),
    .io_in_3_bits_wdata(arbiter_io_in_3_bits_wdata),
    .io_in_3_bits_wmask(arbiter_io_in_3_bits_wmask),
    .io_in_3_bits_wen(arbiter_io_in_3_bits_wen),
    .io_in_3_bits_size(arbiter_io_in_3_bits_size),
    .io_out_ready(arbiter_io_out_ready),
    .io_out_valid(arbiter_io_out_valid),
    .io_out_bits_id(arbiter_io_out_bits_id),
    .io_out_bits_addr(arbiter_io_out_bits_addr),
    .io_out_bits_aen(arbiter_io_out_bits_aen),
    .io_out_bits_wdata(arbiter_io_out_bits_wdata),
    .io_out_bits_wmask(arbiter_io_out_bits_wmask),
    .io_out_bits_wlast(arbiter_io_out_bits_wlast),
    .io_out_bits_wen(arbiter_io_out_bits_wen),
    .io_out_bits_len(arbiter_io_out_bits_len),
    .io_out_bits_size(arbiter_io_out_bits_size),
    .io_chosen(arbiter_io_chosen)
  );
  assign io_in_0_req_ready = arbiter_io_chosen == 2'h0 & io_out_req_ready; // @[Crossbar.scala 20:55]
  assign io_in_0_resp_valid = io_out_resp_bits_id == 4'h1 & io_out_resp_valid; // @[Crossbar.scala 31:25 35:46 37:27]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 30:24]
  assign io_in_0_resp_bits_rlast = io_out_resp_bits_rlast; // @[Crossbar.scala 30:24]
  assign io_in_1_req_ready = arbiter_io_chosen == 2'h1 & io_out_req_ready; // @[Crossbar.scala 20:55]
  assign io_in_1_resp_valid = io_out_resp_bits_id == 4'h2 & io_out_resp_valid; // @[Crossbar.scala 31:25 35:46 37:27]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 30:24]
  assign io_in_1_resp_bits_rlast = io_out_resp_bits_rlast; // @[Crossbar.scala 30:24]
  assign io_in_2_req_ready = arbiter_io_chosen == 2'h2 & io_out_req_ready; // @[Crossbar.scala 20:55]
  assign io_in_2_resp_valid = io_out_resp_bits_id == 4'h3 & io_out_resp_valid; // @[Crossbar.scala 31:25 35:46 37:27]
  assign io_in_2_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 30:24]
  assign io_in_3_req_ready = arbiter_io_chosen == 2'h3 & io_out_req_ready; // @[Crossbar.scala 20:55]
  assign io_in_3_resp_valid = io_out_resp_bits_id == 4'h4 & io_out_resp_valid; // @[Crossbar.scala 31:25 35:46 37:27]
  assign io_in_3_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 30:24]
  assign io_out_req_valid = arbiter_io_out_valid; // @[Crossbar.scala 24:13]
  assign io_out_req_bits_id = arbiter_io_out_bits_id; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_addr = arbiter_io_out_bits_addr; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_aen = arbiter_io_out_bits_aen; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_wdata = arbiter_io_out_bits_wdata; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_wmask = arbiter_io_out_bits_wmask; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_wlast = arbiter_io_out_bits_wlast; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_wen = arbiter_io_out_bits_wen; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_len = arbiter_io_out_bits_len; // @[Crossbar.scala 23:12]
  assign io_out_req_bits_size = arbiter_io_out_bits_size; // @[Crossbar.scala 23:12]
  assign io_out_resp_ready = io_out_resp_bits_id == 4'h4 ? io_in_3_resp_ready : _GEN_4; // @[Crossbar.scala 35:46 36:25]
  assign arbiter_clock = clock;
  assign arbiter_io_in_0_valid = io_in_0_req_valid; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_0_bits_aen = io_in_0_req_bits_aen; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_0_bits_wlast = io_in_0_req_bits_wlast; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_0_bits_wen = io_in_0_req_bits_wen; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_1_valid = io_in_1_req_valid; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_1_bits_aen = io_in_1_req_bits_aen; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_1_bits_wlast = io_in_1_req_bits_wlast; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_1_bits_wen = io_in_1_req_bits_wen; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_2_valid = io_in_2_req_valid; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_2_bits_addr = io_in_2_req_bits_addr; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_2_bits_size = io_in_2_req_bits_size; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_3_valid = io_in_3_req_valid; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_3_bits_addr = io_in_3_req_bits_addr; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_3_bits_wdata = io_in_3_req_bits_wdata; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_3_bits_wmask = io_in_3_req_bits_wmask; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_3_bits_wen = io_in_3_req_bits_wen; // @[Crossbar.scala 15:22]
  assign arbiter_io_in_3_bits_size = io_in_3_req_bits_size; // @[Crossbar.scala 15:22]
  assign arbiter_io_out_ready = io_out_req_ready; // @[Crossbar.scala 25:13]
endmodule
module ysyx_210128_CoreBus2Axi(
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [3:0]  io_in_req_bits_id,
  input  [31:0] io_in_req_bits_addr,
  input         io_in_req_bits_aen,
  input  [63:0] io_in_req_bits_wdata,
  input  [7:0]  io_in_req_bits_wmask,
  input         io_in_req_bits_wlast,
  input         io_in_req_bits_wen,
  input  [7:0]  io_in_req_bits_len,
  input  [1:0]  io_in_req_bits_size,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_id,
  output [63:0] io_in_resp_bits_rdata,
  output        io_in_resp_bits_rlast,
  input         io_out_aw_ready,
  output        io_out_aw_valid,
  output [3:0]  io_out_aw_bits_id,
  output [31:0] io_out_aw_bits_addr,
  output [7:0]  io_out_aw_bits_len,
  output [2:0]  io_out_aw_bits_size,
  input         io_out_w_ready,
  output        io_out_w_valid,
  output [63:0] io_out_w_bits_data,
  output [7:0]  io_out_w_bits_strb,
  output        io_out_w_bits_last,
  output        io_out_b_ready,
  input         io_out_b_valid,
  input  [3:0]  io_out_b_bits_id,
  input         io_out_ar_ready,
  output        io_out_ar_valid,
  output [3:0]  io_out_ar_bits_id,
  output [31:0] io_out_ar_bits_addr,
  output [7:0]  io_out_ar_bits_len,
  output [2:0]  io_out_ar_bits_size,
  output        io_out_r_ready,
  input         io_out_r_valid,
  input  [3:0]  io_out_r_bits_id,
  input  [63:0] io_out_r_bits_data,
  input         io_out_r_bits_last
);
  wire  _T = io_in_req_valid & io_in_req_bits_aen; // @[CoreBus.scala 47:37]
  wire  _T_9 = io_in_req_bits_wen ? io_out_aw_ready & io_out_w_ready : io_out_ar_ready; // @[CoreBus.scala 87:26]
  wire  _T_10 = io_in_req_bits_wen & io_out_w_ready; // @[CoreBus.scala 88:26]
  wire  _GEN_1 = io_out_r_valid & io_in_resp_ready; // @[CoreBus.scala 103:25 105:17 113:17]
  wire [3:0] _GEN_3 = io_out_r_valid ? io_out_r_bits_id : 4'h0; // @[CoreBus.scala 103:25 107:21 115:21]
  wire [63:0] _GEN_4 = io_out_r_valid ? io_out_r_bits_data : 64'h0; // @[CoreBus.scala 103:25 108:24 116:24]
  wire  _GEN_5 = io_out_r_valid & io_out_r_bits_last; // @[CoreBus.scala 103:25 110:24 118:24]
  assign io_in_req_ready = io_in_req_bits_aen ? _T_9 : _T_10; // @[CoreBus.scala 86:22]
  assign io_in_resp_valid = io_out_b_valid ? io_out_b_valid : io_out_r_valid; // @[CoreBus.scala 95:18 98:19]
  assign io_in_resp_bits_id = io_out_b_valid ? io_out_b_bits_id : _GEN_3; // @[CoreBus.scala 95:18 99:21]
  assign io_in_resp_bits_rdata = io_out_b_valid ? 64'h0 : _GEN_4; // @[CoreBus.scala 95:18 100:24]
  assign io_in_resp_bits_rlast = io_out_b_valid ? 1'h0 : _GEN_5; // @[CoreBus.scala 95:18 102:24]
  assign io_out_aw_valid = io_in_req_valid & io_in_req_bits_aen & io_in_req_bits_wen; // @[CoreBus.scala 47:56]
  assign io_out_aw_bits_id = io_in_req_bits_id; // @[CoreBus.scala 49:21]
  assign io_out_aw_bits_addr = io_in_req_bits_addr; // @[CoreBus.scala 48:21]
  assign io_out_aw_bits_len = io_in_req_bits_len; // @[CoreBus.scala 50:21]
  assign io_out_aw_bits_size = {1'h0,io_in_req_bits_size}; // @[Cat.scala 30:58]
  assign io_out_w_valid = io_in_req_valid & io_in_req_bits_wen; // @[CoreBus.scala 62:37]
  assign io_out_w_bits_data = io_in_req_bits_wdata; // @[CoreBus.scala 63:21]
  assign io_out_w_bits_strb = io_in_req_bits_wmask; // @[CoreBus.scala 64:21]
  assign io_out_w_bits_last = io_in_req_bits_wlast; // @[CoreBus.scala 65:21]
  assign io_out_b_ready = io_out_b_valid & io_in_resp_ready; // @[CoreBus.scala 95:18 96:17]
  assign io_out_ar_valid = _T & ~io_in_req_bits_wen; // @[CoreBus.scala 67:56]
  assign io_out_ar_bits_id = io_in_req_bits_id; // @[CoreBus.scala 69:21]
  assign io_out_ar_bits_addr = io_in_req_bits_addr; // @[CoreBus.scala 68:21]
  assign io_out_ar_bits_len = io_in_req_bits_len; // @[CoreBus.scala 70:21]
  assign io_out_ar_bits_size = {1'h0,io_in_req_bits_size}; // @[Cat.scala 30:58]
  assign io_out_r_ready = io_out_b_valid ? 1'h0 : _GEN_1; // @[CoreBus.scala 95:18 97:17]
endmodule
module ysyx_210128(
  input         clock,
  input         reset,
  input         io_interrupt,
  input         io_master_awready,
  output        io_master_awvalid,
  output [3:0]  io_master_awid,
  output [31:0] io_master_awaddr,
  output [7:0]  io_master_awlen,
  output [2:0]  io_master_awsize,
  output [1:0]  io_master_awburst,
  input         io_master_wready,
  output        io_master_wvalid,
  output [63:0] io_master_wdata,
  output [7:0]  io_master_wstrb,
  output        io_master_wlast,
  output        io_master_bready,
  input         io_master_bvalid,
  input  [3:0]  io_master_bid,
  input  [1:0]  io_master_bresp,
  input         io_master_arready,
  output        io_master_arvalid,
  output [3:0]  io_master_arid,
  output [31:0] io_master_araddr,
  output [7:0]  io_master_arlen,
  output [2:0]  io_master_arsize,
  output [1:0]  io_master_arburst,
  output        io_master_rready,
  input         io_master_rvalid,
  input  [3:0]  io_master_rid,
  input  [1:0]  io_master_rresp,
  input  [63:0] io_master_rdata,
  input         io_master_rlast,
  output        io_slave_awready,
  input         io_slave_awvalid,
  input  [3:0]  io_slave_awid,
  input  [31:0] io_slave_awaddr,
  input  [7:0]  io_slave_awlen,
  input  [2:0]  io_slave_awsize,
  input  [1:0]  io_slave_awburst,
  output        io_slave_wready,
  input         io_slave_wvalid,
  input  [63:0] io_slave_wdata,
  input  [7:0]  io_slave_wstrb,
  input         io_slave_wlast,
  input         io_slave_bready,
  output        io_slave_bvalid,
  output [3:0]  io_slave_bid,
  output [1:0]  io_slave_bresp,
  output        io_slave_arready,
  input         io_slave_arvalid,
  input  [3:0]  io_slave_arid,
  input  [31:0] io_slave_araddr,
  input  [7:0]  io_slave_arlen,
  input  [2:0]  io_slave_arsize,
  input  [1:0]  io_slave_arburst,
  input         io_slave_rready,
  output        io_slave_rvalid,
  output [3:0]  io_slave_rid,
  output [1:0]  io_slave_rresp,
  output [63:0] io_slave_rdata,
  output        io_slave_rlast
);
  wire  core_clock; // @[RealTop.scala 13:20]
  wire  core_reset; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_0_req_ready; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_0_req_valid; // @[RealTop.scala 13:20]
  wire [31:0] core_io_core_bus_0_req_bits_addr; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_0_req_bits_aen; // @[RealTop.scala 13:20]
  wire [63:0] core_io_core_bus_0_req_bits_wdata; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_0_req_bits_wlast; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_0_req_bits_wen; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_0_resp_ready; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_0_resp_valid; // @[RealTop.scala 13:20]
  wire [63:0] core_io_core_bus_0_resp_bits_rdata; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_0_resp_bits_rlast; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_1_req_ready; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_1_req_valid; // @[RealTop.scala 13:20]
  wire [31:0] core_io_core_bus_1_req_bits_addr; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_1_req_bits_aen; // @[RealTop.scala 13:20]
  wire [63:0] core_io_core_bus_1_req_bits_wdata; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_1_req_bits_wlast; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_1_req_bits_wen; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_1_resp_ready; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_1_resp_valid; // @[RealTop.scala 13:20]
  wire [63:0] core_io_core_bus_1_resp_bits_rdata; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_1_resp_bits_rlast; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_2_req_ready; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_2_req_valid; // @[RealTop.scala 13:20]
  wire [31:0] core_io_core_bus_2_req_bits_addr; // @[RealTop.scala 13:20]
  wire [1:0] core_io_core_bus_2_req_bits_size; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_2_resp_ready; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_2_resp_valid; // @[RealTop.scala 13:20]
  wire [63:0] core_io_core_bus_2_resp_bits_rdata; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_3_req_ready; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_3_req_valid; // @[RealTop.scala 13:20]
  wire [31:0] core_io_core_bus_3_req_bits_addr; // @[RealTop.scala 13:20]
  wire [63:0] core_io_core_bus_3_req_bits_wdata; // @[RealTop.scala 13:20]
  wire [7:0] core_io_core_bus_3_req_bits_wmask; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_3_req_bits_wen; // @[RealTop.scala 13:20]
  wire [1:0] core_io_core_bus_3_req_bits_size; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_3_resp_ready; // @[RealTop.scala 13:20]
  wire  core_io_core_bus_3_resp_valid; // @[RealTop.scala 13:20]
  wire [63:0] core_io_core_bus_3_resp_bits_rdata; // @[RealTop.scala 13:20]
  wire  crossbar_clock; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_0_req_ready; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_0_req_valid; // @[RealTop.scala 15:24]
  wire [31:0] crossbar_io_in_0_req_bits_addr; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_0_req_bits_aen; // @[RealTop.scala 15:24]
  wire [63:0] crossbar_io_in_0_req_bits_wdata; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_0_req_bits_wlast; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_0_req_bits_wen; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_0_resp_ready; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_0_resp_valid; // @[RealTop.scala 15:24]
  wire [63:0] crossbar_io_in_0_resp_bits_rdata; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_0_resp_bits_rlast; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_1_req_ready; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_1_req_valid; // @[RealTop.scala 15:24]
  wire [31:0] crossbar_io_in_1_req_bits_addr; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_1_req_bits_aen; // @[RealTop.scala 15:24]
  wire [63:0] crossbar_io_in_1_req_bits_wdata; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_1_req_bits_wlast; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_1_req_bits_wen; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_1_resp_ready; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_1_resp_valid; // @[RealTop.scala 15:24]
  wire [63:0] crossbar_io_in_1_resp_bits_rdata; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_1_resp_bits_rlast; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_2_req_ready; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_2_req_valid; // @[RealTop.scala 15:24]
  wire [31:0] crossbar_io_in_2_req_bits_addr; // @[RealTop.scala 15:24]
  wire [1:0] crossbar_io_in_2_req_bits_size; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_2_resp_ready; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_2_resp_valid; // @[RealTop.scala 15:24]
  wire [63:0] crossbar_io_in_2_resp_bits_rdata; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_3_req_ready; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_3_req_valid; // @[RealTop.scala 15:24]
  wire [31:0] crossbar_io_in_3_req_bits_addr; // @[RealTop.scala 15:24]
  wire [63:0] crossbar_io_in_3_req_bits_wdata; // @[RealTop.scala 15:24]
  wire [7:0] crossbar_io_in_3_req_bits_wmask; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_3_req_bits_wen; // @[RealTop.scala 15:24]
  wire [1:0] crossbar_io_in_3_req_bits_size; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_3_resp_ready; // @[RealTop.scala 15:24]
  wire  crossbar_io_in_3_resp_valid; // @[RealTop.scala 15:24]
  wire [63:0] crossbar_io_in_3_resp_bits_rdata; // @[RealTop.scala 15:24]
  wire  crossbar_io_out_req_ready; // @[RealTop.scala 15:24]
  wire  crossbar_io_out_req_valid; // @[RealTop.scala 15:24]
  wire [3:0] crossbar_io_out_req_bits_id; // @[RealTop.scala 15:24]
  wire [31:0] crossbar_io_out_req_bits_addr; // @[RealTop.scala 15:24]
  wire  crossbar_io_out_req_bits_aen; // @[RealTop.scala 15:24]
  wire [63:0] crossbar_io_out_req_bits_wdata; // @[RealTop.scala 15:24]
  wire [7:0] crossbar_io_out_req_bits_wmask; // @[RealTop.scala 15:24]
  wire  crossbar_io_out_req_bits_wlast; // @[RealTop.scala 15:24]
  wire  crossbar_io_out_req_bits_wen; // @[RealTop.scala 15:24]
  wire [7:0] crossbar_io_out_req_bits_len; // @[RealTop.scala 15:24]
  wire [1:0] crossbar_io_out_req_bits_size; // @[RealTop.scala 15:24]
  wire  crossbar_io_out_resp_ready; // @[RealTop.scala 15:24]
  wire  crossbar_io_out_resp_valid; // @[RealTop.scala 15:24]
  wire [3:0] crossbar_io_out_resp_bits_id; // @[RealTop.scala 15:24]
  wire [63:0] crossbar_io_out_resp_bits_rdata; // @[RealTop.scala 15:24]
  wire  crossbar_io_out_resp_bits_rlast; // @[RealTop.scala 15:24]
  wire  core2axi_io_in_req_ready; // @[RealTop.scala 18:24]
  wire  core2axi_io_in_req_valid; // @[RealTop.scala 18:24]
  wire [3:0] core2axi_io_in_req_bits_id; // @[RealTop.scala 18:24]
  wire [31:0] core2axi_io_in_req_bits_addr; // @[RealTop.scala 18:24]
  wire  core2axi_io_in_req_bits_aen; // @[RealTop.scala 18:24]
  wire [63:0] core2axi_io_in_req_bits_wdata; // @[RealTop.scala 18:24]
  wire [7:0] core2axi_io_in_req_bits_wmask; // @[RealTop.scala 18:24]
  wire  core2axi_io_in_req_bits_wlast; // @[RealTop.scala 18:24]
  wire  core2axi_io_in_req_bits_wen; // @[RealTop.scala 18:24]
  wire [7:0] core2axi_io_in_req_bits_len; // @[RealTop.scala 18:24]
  wire [1:0] core2axi_io_in_req_bits_size; // @[RealTop.scala 18:24]
  wire  core2axi_io_in_resp_ready; // @[RealTop.scala 18:24]
  wire  core2axi_io_in_resp_valid; // @[RealTop.scala 18:24]
  wire [3:0] core2axi_io_in_resp_bits_id; // @[RealTop.scala 18:24]
  wire [63:0] core2axi_io_in_resp_bits_rdata; // @[RealTop.scala 18:24]
  wire  core2axi_io_in_resp_bits_rlast; // @[RealTop.scala 18:24]
  wire  core2axi_io_out_aw_ready; // @[RealTop.scala 18:24]
  wire  core2axi_io_out_aw_valid; // @[RealTop.scala 18:24]
  wire [3:0] core2axi_io_out_aw_bits_id; // @[RealTop.scala 18:24]
  wire [31:0] core2axi_io_out_aw_bits_addr; // @[RealTop.scala 18:24]
  wire [7:0] core2axi_io_out_aw_bits_len; // @[RealTop.scala 18:24]
  wire [2:0] core2axi_io_out_aw_bits_size; // @[RealTop.scala 18:24]
  wire  core2axi_io_out_w_ready; // @[RealTop.scala 18:24]
  wire  core2axi_io_out_w_valid; // @[RealTop.scala 18:24]
  wire [63:0] core2axi_io_out_w_bits_data; // @[RealTop.scala 18:24]
  wire [7:0] core2axi_io_out_w_bits_strb; // @[RealTop.scala 18:24]
  wire  core2axi_io_out_w_bits_last; // @[RealTop.scala 18:24]
  wire  core2axi_io_out_b_ready; // @[RealTop.scala 18:24]
  wire  core2axi_io_out_b_valid; // @[RealTop.scala 18:24]
  wire [3:0] core2axi_io_out_b_bits_id; // @[RealTop.scala 18:24]
  wire  core2axi_io_out_ar_ready; // @[RealTop.scala 18:24]
  wire  core2axi_io_out_ar_valid; // @[RealTop.scala 18:24]
  wire [3:0] core2axi_io_out_ar_bits_id; // @[RealTop.scala 18:24]
  wire [31:0] core2axi_io_out_ar_bits_addr; // @[RealTop.scala 18:24]
  wire [7:0] core2axi_io_out_ar_bits_len; // @[RealTop.scala 18:24]
  wire [2:0] core2axi_io_out_ar_bits_size; // @[RealTop.scala 18:24]
  wire  core2axi_io_out_r_ready; // @[RealTop.scala 18:24]
  wire  core2axi_io_out_r_valid; // @[RealTop.scala 18:24]
  wire [3:0] core2axi_io_out_r_bits_id; // @[RealTop.scala 18:24]
  wire [63:0] core2axi_io_out_r_bits_data; // @[RealTop.scala 18:24]
  wire  core2axi_io_out_r_bits_last; // @[RealTop.scala 18:24]
  ysyx_210128_Core core ( // @[RealTop.scala 13:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_core_bus_0_req_ready(core_io_core_bus_0_req_ready),
    .io_core_bus_0_req_valid(core_io_core_bus_0_req_valid),
    .io_core_bus_0_req_bits_addr(core_io_core_bus_0_req_bits_addr),
    .io_core_bus_0_req_bits_aen(core_io_core_bus_0_req_bits_aen),
    .io_core_bus_0_req_bits_wdata(core_io_core_bus_0_req_bits_wdata),
    .io_core_bus_0_req_bits_wlast(core_io_core_bus_0_req_bits_wlast),
    .io_core_bus_0_req_bits_wen(core_io_core_bus_0_req_bits_wen),
    .io_core_bus_0_resp_ready(core_io_core_bus_0_resp_ready),
    .io_core_bus_0_resp_valid(core_io_core_bus_0_resp_valid),
    .io_core_bus_0_resp_bits_rdata(core_io_core_bus_0_resp_bits_rdata),
    .io_core_bus_0_resp_bits_rlast(core_io_core_bus_0_resp_bits_rlast),
    .io_core_bus_1_req_ready(core_io_core_bus_1_req_ready),
    .io_core_bus_1_req_valid(core_io_core_bus_1_req_valid),
    .io_core_bus_1_req_bits_addr(core_io_core_bus_1_req_bits_addr),
    .io_core_bus_1_req_bits_aen(core_io_core_bus_1_req_bits_aen),
    .io_core_bus_1_req_bits_wdata(core_io_core_bus_1_req_bits_wdata),
    .io_core_bus_1_req_bits_wlast(core_io_core_bus_1_req_bits_wlast),
    .io_core_bus_1_req_bits_wen(core_io_core_bus_1_req_bits_wen),
    .io_core_bus_1_resp_ready(core_io_core_bus_1_resp_ready),
    .io_core_bus_1_resp_valid(core_io_core_bus_1_resp_valid),
    .io_core_bus_1_resp_bits_rdata(core_io_core_bus_1_resp_bits_rdata),
    .io_core_bus_1_resp_bits_rlast(core_io_core_bus_1_resp_bits_rlast),
    .io_core_bus_2_req_ready(core_io_core_bus_2_req_ready),
    .io_core_bus_2_req_valid(core_io_core_bus_2_req_valid),
    .io_core_bus_2_req_bits_addr(core_io_core_bus_2_req_bits_addr),
    .io_core_bus_2_req_bits_size(core_io_core_bus_2_req_bits_size),
    .io_core_bus_2_resp_ready(core_io_core_bus_2_resp_ready),
    .io_core_bus_2_resp_valid(core_io_core_bus_2_resp_valid),
    .io_core_bus_2_resp_bits_rdata(core_io_core_bus_2_resp_bits_rdata),
    .io_core_bus_3_req_ready(core_io_core_bus_3_req_ready),
    .io_core_bus_3_req_valid(core_io_core_bus_3_req_valid),
    .io_core_bus_3_req_bits_addr(core_io_core_bus_3_req_bits_addr),
    .io_core_bus_3_req_bits_wdata(core_io_core_bus_3_req_bits_wdata),
    .io_core_bus_3_req_bits_wmask(core_io_core_bus_3_req_bits_wmask),
    .io_core_bus_3_req_bits_wen(core_io_core_bus_3_req_bits_wen),
    .io_core_bus_3_req_bits_size(core_io_core_bus_3_req_bits_size),
    .io_core_bus_3_resp_ready(core_io_core_bus_3_resp_ready),
    .io_core_bus_3_resp_valid(core_io_core_bus_3_resp_valid),
    .io_core_bus_3_resp_bits_rdata(core_io_core_bus_3_resp_bits_rdata)
  );
  ysyx_210128_CoreBusCrossbarNto1 crossbar ( // @[RealTop.scala 15:24]
    .clock(crossbar_clock),
    .io_in_0_req_ready(crossbar_io_in_0_req_ready),
    .io_in_0_req_valid(crossbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(crossbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_aen(crossbar_io_in_0_req_bits_aen),
    .io_in_0_req_bits_wdata(crossbar_io_in_0_req_bits_wdata),
    .io_in_0_req_bits_wlast(crossbar_io_in_0_req_bits_wlast),
    .io_in_0_req_bits_wen(crossbar_io_in_0_req_bits_wen),
    .io_in_0_resp_ready(crossbar_io_in_0_resp_ready),
    .io_in_0_resp_valid(crossbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(crossbar_io_in_0_resp_bits_rdata),
    .io_in_0_resp_bits_rlast(crossbar_io_in_0_resp_bits_rlast),
    .io_in_1_req_ready(crossbar_io_in_1_req_ready),
    .io_in_1_req_valid(crossbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(crossbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_aen(crossbar_io_in_1_req_bits_aen),
    .io_in_1_req_bits_wdata(crossbar_io_in_1_req_bits_wdata),
    .io_in_1_req_bits_wlast(crossbar_io_in_1_req_bits_wlast),
    .io_in_1_req_bits_wen(crossbar_io_in_1_req_bits_wen),
    .io_in_1_resp_ready(crossbar_io_in_1_resp_ready),
    .io_in_1_resp_valid(crossbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_rdata(crossbar_io_in_1_resp_bits_rdata),
    .io_in_1_resp_bits_rlast(crossbar_io_in_1_resp_bits_rlast),
    .io_in_2_req_ready(crossbar_io_in_2_req_ready),
    .io_in_2_req_valid(crossbar_io_in_2_req_valid),
    .io_in_2_req_bits_addr(crossbar_io_in_2_req_bits_addr),
    .io_in_2_req_bits_size(crossbar_io_in_2_req_bits_size),
    .io_in_2_resp_ready(crossbar_io_in_2_resp_ready),
    .io_in_2_resp_valid(crossbar_io_in_2_resp_valid),
    .io_in_2_resp_bits_rdata(crossbar_io_in_2_resp_bits_rdata),
    .io_in_3_req_ready(crossbar_io_in_3_req_ready),
    .io_in_3_req_valid(crossbar_io_in_3_req_valid),
    .io_in_3_req_bits_addr(crossbar_io_in_3_req_bits_addr),
    .io_in_3_req_bits_wdata(crossbar_io_in_3_req_bits_wdata),
    .io_in_3_req_bits_wmask(crossbar_io_in_3_req_bits_wmask),
    .io_in_3_req_bits_wen(crossbar_io_in_3_req_bits_wen),
    .io_in_3_req_bits_size(crossbar_io_in_3_req_bits_size),
    .io_in_3_resp_ready(crossbar_io_in_3_resp_ready),
    .io_in_3_resp_valid(crossbar_io_in_3_resp_valid),
    .io_in_3_resp_bits_rdata(crossbar_io_in_3_resp_bits_rdata),
    .io_out_req_ready(crossbar_io_out_req_ready),
    .io_out_req_valid(crossbar_io_out_req_valid),
    .io_out_req_bits_id(crossbar_io_out_req_bits_id),
    .io_out_req_bits_addr(crossbar_io_out_req_bits_addr),
    .io_out_req_bits_aen(crossbar_io_out_req_bits_aen),
    .io_out_req_bits_wdata(crossbar_io_out_req_bits_wdata),
    .io_out_req_bits_wmask(crossbar_io_out_req_bits_wmask),
    .io_out_req_bits_wlast(crossbar_io_out_req_bits_wlast),
    .io_out_req_bits_wen(crossbar_io_out_req_bits_wen),
    .io_out_req_bits_len(crossbar_io_out_req_bits_len),
    .io_out_req_bits_size(crossbar_io_out_req_bits_size),
    .io_out_resp_ready(crossbar_io_out_resp_ready),
    .io_out_resp_valid(crossbar_io_out_resp_valid),
    .io_out_resp_bits_id(crossbar_io_out_resp_bits_id),
    .io_out_resp_bits_rdata(crossbar_io_out_resp_bits_rdata),
    .io_out_resp_bits_rlast(crossbar_io_out_resp_bits_rlast)
  );
  ysyx_210128_CoreBus2Axi core2axi ( // @[RealTop.scala 18:24]
    .io_in_req_ready(core2axi_io_in_req_ready),
    .io_in_req_valid(core2axi_io_in_req_valid),
    .io_in_req_bits_id(core2axi_io_in_req_bits_id),
    .io_in_req_bits_addr(core2axi_io_in_req_bits_addr),
    .io_in_req_bits_aen(core2axi_io_in_req_bits_aen),
    .io_in_req_bits_wdata(core2axi_io_in_req_bits_wdata),
    .io_in_req_bits_wmask(core2axi_io_in_req_bits_wmask),
    .io_in_req_bits_wlast(core2axi_io_in_req_bits_wlast),
    .io_in_req_bits_wen(core2axi_io_in_req_bits_wen),
    .io_in_req_bits_len(core2axi_io_in_req_bits_len),
    .io_in_req_bits_size(core2axi_io_in_req_bits_size),
    .io_in_resp_ready(core2axi_io_in_resp_ready),
    .io_in_resp_valid(core2axi_io_in_resp_valid),
    .io_in_resp_bits_id(core2axi_io_in_resp_bits_id),
    .io_in_resp_bits_rdata(core2axi_io_in_resp_bits_rdata),
    .io_in_resp_bits_rlast(core2axi_io_in_resp_bits_rlast),
    .io_out_aw_ready(core2axi_io_out_aw_ready),
    .io_out_aw_valid(core2axi_io_out_aw_valid),
    .io_out_aw_bits_id(core2axi_io_out_aw_bits_id),
    .io_out_aw_bits_addr(core2axi_io_out_aw_bits_addr),
    .io_out_aw_bits_len(core2axi_io_out_aw_bits_len),
    .io_out_aw_bits_size(core2axi_io_out_aw_bits_size),
    .io_out_w_ready(core2axi_io_out_w_ready),
    .io_out_w_valid(core2axi_io_out_w_valid),
    .io_out_w_bits_data(core2axi_io_out_w_bits_data),
    .io_out_w_bits_strb(core2axi_io_out_w_bits_strb),
    .io_out_w_bits_last(core2axi_io_out_w_bits_last),
    .io_out_b_ready(core2axi_io_out_b_ready),
    .io_out_b_valid(core2axi_io_out_b_valid),
    .io_out_b_bits_id(core2axi_io_out_b_bits_id),
    .io_out_ar_ready(core2axi_io_out_ar_ready),
    .io_out_ar_valid(core2axi_io_out_ar_valid),
    .io_out_ar_bits_id(core2axi_io_out_ar_bits_id),
    .io_out_ar_bits_addr(core2axi_io_out_ar_bits_addr),
    .io_out_ar_bits_len(core2axi_io_out_ar_bits_len),
    .io_out_ar_bits_size(core2axi_io_out_ar_bits_size),
    .io_out_r_ready(core2axi_io_out_r_ready),
    .io_out_r_valid(core2axi_io_out_r_valid),
    .io_out_r_bits_id(core2axi_io_out_r_bits_id),
    .io_out_r_bits_data(core2axi_io_out_r_bits_data),
    .io_out_r_bits_last(core2axi_io_out_r_bits_last)
  );
  assign io_master_awvalid = core2axi_io_out_aw_valid; // @[RealTop.scala 20:16]
  assign io_master_awid = core2axi_io_out_aw_bits_id; // @[RealTop.scala 20:16]
  assign io_master_awaddr = core2axi_io_out_aw_bits_addr; // @[RealTop.scala 20:16]
  assign io_master_awlen = core2axi_io_out_aw_bits_len; // @[RealTop.scala 20:16]
  assign io_master_awsize = core2axi_io_out_aw_bits_size; // @[RealTop.scala 20:16]
  assign io_master_awburst = 2'h1; // @[RealTop.scala 20:16]
  assign io_master_wvalid = core2axi_io_out_w_valid; // @[RealTop.scala 20:16]
  assign io_master_wdata = core2axi_io_out_w_bits_data; // @[RealTop.scala 20:16]
  assign io_master_wstrb = core2axi_io_out_w_bits_strb; // @[RealTop.scala 20:16]
  assign io_master_wlast = core2axi_io_out_w_bits_last; // @[RealTop.scala 20:16]
  assign io_master_bready = core2axi_io_out_b_ready; // @[RealTop.scala 20:16]
  assign io_master_arvalid = core2axi_io_out_ar_valid; // @[RealTop.scala 20:16]
  assign io_master_arid = core2axi_io_out_ar_bits_id; // @[RealTop.scala 20:16]
  assign io_master_araddr = core2axi_io_out_ar_bits_addr; // @[RealTop.scala 20:16]
  assign io_master_arlen = core2axi_io_out_ar_bits_len; // @[RealTop.scala 20:16]
  assign io_master_arsize = core2axi_io_out_ar_bits_size; // @[RealTop.scala 20:16]
  assign io_master_arburst = 2'h1; // @[RealTop.scala 20:16]
  assign io_master_rready = core2axi_io_out_r_ready; // @[RealTop.scala 20:16]
  assign io_slave_awready = 1'h0; // @[RealTop.scala 23:21]
  assign io_slave_wready = 1'h0; // @[RealTop.scala 24:21]
  assign io_slave_bvalid = 1'h0; // @[RealTop.scala 25:21]
  assign io_slave_bid = 4'h0; // @[RealTop.scala 27:21]
  assign io_slave_bresp = 2'h0; // @[RealTop.scala 26:21]
  assign io_slave_arready = 1'h0; // @[RealTop.scala 28:21]
  assign io_slave_rvalid = 1'h0; // @[RealTop.scala 29:21]
  assign io_slave_rid = 4'h0; // @[RealTop.scala 33:21]
  assign io_slave_rresp = 2'h0; // @[RealTop.scala 30:21]
  assign io_slave_rdata = 64'h0; // @[RealTop.scala 31:21]
  assign io_slave_rlast = 1'h0; // @[RealTop.scala 32:21]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_core_bus_0_req_ready = crossbar_io_in_0_req_ready; // @[RealTop.scala 16:18]
  assign core_io_core_bus_0_resp_valid = crossbar_io_in_0_resp_valid; // @[RealTop.scala 16:18]
  assign core_io_core_bus_0_resp_bits_rdata = crossbar_io_in_0_resp_bits_rdata; // @[RealTop.scala 16:18]
  assign core_io_core_bus_0_resp_bits_rlast = crossbar_io_in_0_resp_bits_rlast; // @[RealTop.scala 16:18]
  assign core_io_core_bus_1_req_ready = crossbar_io_in_1_req_ready; // @[RealTop.scala 16:18]
  assign core_io_core_bus_1_resp_valid = crossbar_io_in_1_resp_valid; // @[RealTop.scala 16:18]
  assign core_io_core_bus_1_resp_bits_rdata = crossbar_io_in_1_resp_bits_rdata; // @[RealTop.scala 16:18]
  assign core_io_core_bus_1_resp_bits_rlast = crossbar_io_in_1_resp_bits_rlast; // @[RealTop.scala 16:18]
  assign core_io_core_bus_2_req_ready = crossbar_io_in_2_req_ready; // @[RealTop.scala 16:18]
  assign core_io_core_bus_2_resp_valid = crossbar_io_in_2_resp_valid; // @[RealTop.scala 16:18]
  assign core_io_core_bus_2_resp_bits_rdata = crossbar_io_in_2_resp_bits_rdata; // @[RealTop.scala 16:18]
  assign core_io_core_bus_3_req_ready = crossbar_io_in_3_req_ready; // @[RealTop.scala 16:18]
  assign core_io_core_bus_3_resp_valid = crossbar_io_in_3_resp_valid; // @[RealTop.scala 16:18]
  assign core_io_core_bus_3_resp_bits_rdata = crossbar_io_in_3_resp_bits_rdata; // @[RealTop.scala 16:18]
  assign crossbar_clock = clock;
  assign crossbar_io_in_0_req_valid = core_io_core_bus_0_req_valid; // @[RealTop.scala 16:18]
  assign crossbar_io_in_0_req_bits_addr = core_io_core_bus_0_req_bits_addr; // @[RealTop.scala 16:18]
  assign crossbar_io_in_0_req_bits_aen = core_io_core_bus_0_req_bits_aen; // @[RealTop.scala 16:18]
  assign crossbar_io_in_0_req_bits_wdata = core_io_core_bus_0_req_bits_wdata; // @[RealTop.scala 16:18]
  assign crossbar_io_in_0_req_bits_wlast = core_io_core_bus_0_req_bits_wlast; // @[RealTop.scala 16:18]
  assign crossbar_io_in_0_req_bits_wen = core_io_core_bus_0_req_bits_wen; // @[RealTop.scala 16:18]
  assign crossbar_io_in_0_resp_ready = core_io_core_bus_0_resp_ready; // @[RealTop.scala 16:18]
  assign crossbar_io_in_1_req_valid = core_io_core_bus_1_req_valid; // @[RealTop.scala 16:18]
  assign crossbar_io_in_1_req_bits_addr = core_io_core_bus_1_req_bits_addr; // @[RealTop.scala 16:18]
  assign crossbar_io_in_1_req_bits_aen = core_io_core_bus_1_req_bits_aen; // @[RealTop.scala 16:18]
  assign crossbar_io_in_1_req_bits_wdata = core_io_core_bus_1_req_bits_wdata; // @[RealTop.scala 16:18]
  assign crossbar_io_in_1_req_bits_wlast = core_io_core_bus_1_req_bits_wlast; // @[RealTop.scala 16:18]
  assign crossbar_io_in_1_req_bits_wen = core_io_core_bus_1_req_bits_wen; // @[RealTop.scala 16:18]
  assign crossbar_io_in_1_resp_ready = core_io_core_bus_1_resp_ready; // @[RealTop.scala 16:18]
  assign crossbar_io_in_2_req_valid = core_io_core_bus_2_req_valid; // @[RealTop.scala 16:18]
  assign crossbar_io_in_2_req_bits_addr = core_io_core_bus_2_req_bits_addr; // @[RealTop.scala 16:18]
  assign crossbar_io_in_2_req_bits_size = core_io_core_bus_2_req_bits_size; // @[RealTop.scala 16:18]
  assign crossbar_io_in_2_resp_ready = core_io_core_bus_2_resp_ready; // @[RealTop.scala 16:18]
  assign crossbar_io_in_3_req_valid = core_io_core_bus_3_req_valid; // @[RealTop.scala 16:18]
  assign crossbar_io_in_3_req_bits_addr = core_io_core_bus_3_req_bits_addr; // @[RealTop.scala 16:18]
  assign crossbar_io_in_3_req_bits_wdata = core_io_core_bus_3_req_bits_wdata; // @[RealTop.scala 16:18]
  assign crossbar_io_in_3_req_bits_wmask = core_io_core_bus_3_req_bits_wmask; // @[RealTop.scala 16:18]
  assign crossbar_io_in_3_req_bits_wen = core_io_core_bus_3_req_bits_wen; // @[RealTop.scala 16:18]
  assign crossbar_io_in_3_req_bits_size = core_io_core_bus_3_req_bits_size; // @[RealTop.scala 16:18]
  assign crossbar_io_in_3_resp_ready = core_io_core_bus_3_resp_ready; // @[RealTop.scala 16:18]
  assign crossbar_io_out_req_ready = core2axi_io_in_req_ready; // @[RealTop.scala 19:15]
  assign crossbar_io_out_resp_valid = core2axi_io_in_resp_valid; // @[RealTop.scala 19:15]
  assign crossbar_io_out_resp_bits_id = core2axi_io_in_resp_bits_id; // @[RealTop.scala 19:15]
  assign crossbar_io_out_resp_bits_rdata = core2axi_io_in_resp_bits_rdata; // @[RealTop.scala 19:15]
  assign crossbar_io_out_resp_bits_rlast = core2axi_io_in_resp_bits_rlast; // @[RealTop.scala 19:15]
  assign core2axi_io_in_req_valid = crossbar_io_out_req_valid; // @[RealTop.scala 19:15]
  assign core2axi_io_in_req_bits_id = crossbar_io_out_req_bits_id; // @[RealTop.scala 19:15]
  assign core2axi_io_in_req_bits_addr = crossbar_io_out_req_bits_addr; // @[RealTop.scala 19:15]
  assign core2axi_io_in_req_bits_aen = crossbar_io_out_req_bits_aen; // @[RealTop.scala 19:15]
  assign core2axi_io_in_req_bits_wdata = crossbar_io_out_req_bits_wdata; // @[RealTop.scala 19:15]
  assign core2axi_io_in_req_bits_wmask = crossbar_io_out_req_bits_wmask; // @[RealTop.scala 19:15]
  assign core2axi_io_in_req_bits_wlast = crossbar_io_out_req_bits_wlast; // @[RealTop.scala 19:15]
  assign core2axi_io_in_req_bits_wen = crossbar_io_out_req_bits_wen; // @[RealTop.scala 19:15]
  assign core2axi_io_in_req_bits_len = crossbar_io_out_req_bits_len; // @[RealTop.scala 19:15]
  assign core2axi_io_in_req_bits_size = crossbar_io_out_req_bits_size; // @[RealTop.scala 19:15]
  assign core2axi_io_in_resp_ready = crossbar_io_out_resp_ready; // @[RealTop.scala 19:15]
  assign core2axi_io_out_aw_ready = io_master_awready; // @[RealTop.scala 20:16]
  assign core2axi_io_out_w_ready = io_master_wready; // @[RealTop.scala 20:16]
  assign core2axi_io_out_b_valid = io_master_bvalid; // @[RealTop.scala 20:16]
  assign core2axi_io_out_b_bits_id = io_master_bid; // @[RealTop.scala 20:16]
  assign core2axi_io_out_ar_ready = io_master_arready; // @[RealTop.scala 20:16]
  assign core2axi_io_out_r_valid = io_master_rvalid; // @[RealTop.scala 20:16]
  assign core2axi_io_out_r_bits_id = io_master_rid; // @[RealTop.scala 20:16]
  assign core2axi_io_out_r_bits_data = io_master_rdata; // @[RealTop.scala 20:16]
  assign core2axi_io_out_r_bits_last = io_master_rlast; // @[RealTop.scala 20:16]
endmodule
