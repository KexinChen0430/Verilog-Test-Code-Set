module ass(a, b, out);
    input [1:0] a;
    output [1:0] out;
    assign out = a;
endmodule