module  add2 ( count,sum,a,b,cin );
  input a, b; 
  output  count; 
  output sum; 
  assign {count,sum} = a + b; 
endmodule 