module page33;

integer a;              // integer value
time last_chng;        // time value
real float ;// a variable to store a real value
realtime rtime ;// a variable to store time as a real value

endmodule