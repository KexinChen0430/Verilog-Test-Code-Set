module page251;

specify
$nochange( posedge clk, data, 0, 0) ;
endspecify
endmodule